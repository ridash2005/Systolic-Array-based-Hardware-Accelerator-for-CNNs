VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Systolic4x4_serial_io
  CLASS BLOCK ;
  FOREIGN Systolic4x4_serial_io ;
  ORIGIN 0.000 0.000 ;
  SIZE 672.655 BY 683.375 ;
  PIN A_in_frame_sync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END A_in_frame_sync
  PIN A_in_serial_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END A_in_serial_clk
  PIN A_in_serial_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END A_in_serial_data
  PIN B_in_frame_sync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END B_in_frame_sync
  PIN B_in_serial_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END B_in_serial_clk
  PIN B_in_serial_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END B_in_serial_data
  PIN C_out_frame_sync
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END C_out_frame_sync
  PIN C_out_serial_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 25.850 679.375 26.130 683.375 ;
    END
  END C_out_serial_clk
  PIN C_out_serial_data
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 244.810 679.375 245.090 683.375 ;
    END
  END C_out_serial_data
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 672.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 667.240 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 667.240 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 667.240 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 667.240 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 667.240 644.350 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 672.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 667.240 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 667.240 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 667.240 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 667.240 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 667.240 641.050 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 196.510 679.375 196.790 683.375 ;
    END
  END done
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END rst_n
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END start
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 667.190 672.030 ;
      LAYER li1 ;
        RECT 5.520 10.795 667.000 671.925 ;
      LAYER met1 ;
        RECT 0.530 0.380 667.300 672.080 ;
      LAYER met2 ;
        RECT 0.550 679.095 25.570 679.375 ;
        RECT 26.410 679.095 196.230 679.375 ;
        RECT 197.070 679.095 244.530 679.375 ;
        RECT 245.370 679.095 665.520 679.375 ;
        RECT 0.550 4.280 665.520 679.095 ;
        RECT 0.550 0.350 19.130 4.280 ;
        RECT 19.970 0.350 186.570 4.280 ;
        RECT 187.410 0.350 665.520 4.280 ;
      LAYER met3 ;
        RECT 0.525 650.440 652.675 672.005 ;
        RECT 4.400 649.040 652.675 650.440 ;
        RECT 0.525 592.640 652.675 649.040 ;
        RECT 4.400 591.240 652.675 592.640 ;
        RECT 0.525 449.840 652.675 591.240 ;
        RECT 4.400 448.440 652.675 449.840 ;
        RECT 0.525 446.440 652.675 448.440 ;
        RECT 4.400 445.040 652.675 446.440 ;
        RECT 0.525 398.840 652.675 445.040 ;
        RECT 4.400 397.440 652.675 398.840 ;
        RECT 0.525 337.640 652.675 397.440 ;
        RECT 4.400 336.240 652.675 337.640 ;
        RECT 0.525 242.440 652.675 336.240 ;
        RECT 4.400 241.040 652.675 242.440 ;
        RECT 0.525 239.040 652.675 241.040 ;
        RECT 4.400 237.640 652.675 239.040 ;
        RECT 0.525 10.715 652.675 237.640 ;
      LAYER met4 ;
        RECT 3.975 82.455 20.640 618.625 ;
        RECT 23.040 82.455 23.940 618.625 ;
        RECT 26.340 82.455 174.240 618.625 ;
        RECT 176.640 82.455 177.540 618.625 ;
        RECT 179.940 82.455 327.840 618.625 ;
        RECT 330.240 82.455 331.140 618.625 ;
        RECT 333.540 82.455 481.440 618.625 ;
        RECT 483.840 82.455 484.740 618.625 ;
        RECT 487.140 82.455 635.040 618.625 ;
        RECT 637.440 82.455 638.340 618.625 ;
        RECT 640.740 82.455 642.785 618.625 ;
  END
END Systolic4x4_serial_io
END LIBRARY

