VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Systolic4x4_serial_io
  CLASS BLOCK ;
  FOREIGN Systolic4x4_serial_io ;
  ORIGIN 0.000 0.000 ;
  SIZE 191.040 BY 201.760 ;
  PIN A_in_frame_sync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 187.040 81.640 191.040 82.240 ;
    END
  END A_in_frame_sync
  PIN A_in_serial_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END A_in_serial_clk
  PIN A_in_serial_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END A_in_serial_data
  PIN B_in_frame_sync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 197.760 148.490 201.760 ;
    END
  END B_in_frame_sync
  PIN B_in_serial_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 197.760 154.930 201.760 ;
    END
  END B_in_serial_clk
  PIN B_in_serial_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 197.760 125.950 201.760 ;
    END
  END B_in_serial_data
  PIN C_out_frame_sync
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END C_out_frame_sync
  PIN C_out_serial_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END C_out_serial_clk
  PIN C_out_serial_data
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 187.040 30.640 191.040 31.240 ;
    END
  END C_out_serial_data
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 190.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 190.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 185.620 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 185.620 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 190.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 190.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 185.620 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 185.620 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END done
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END rst_n
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END start
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 185.570 190.485 ;
      LAYER li1 ;
        RECT 5.520 10.795 185.380 190.485 ;
      LAYER met1 ;
        RECT 4.210 10.640 185.380 190.640 ;
      LAYER met2 ;
        RECT 4.230 197.480 125.390 198.290 ;
        RECT 126.230 197.480 147.930 198.290 ;
        RECT 148.770 197.480 154.370 198.290 ;
        RECT 155.210 197.480 183.910 198.290 ;
        RECT 4.230 4.280 183.910 197.480 ;
        RECT 4.230 4.000 51.330 4.280 ;
        RECT 52.170 4.000 115.730 4.280 ;
        RECT 116.570 4.000 183.910 4.280 ;
      LAYER met3 ;
        RECT 3.990 184.640 187.040 190.565 ;
        RECT 4.400 183.240 187.040 184.640 ;
        RECT 3.990 147.240 187.040 183.240 ;
        RECT 4.400 145.840 187.040 147.240 ;
        RECT 3.990 126.840 187.040 145.840 ;
        RECT 4.400 125.440 187.040 126.840 ;
        RECT 3.990 120.040 187.040 125.440 ;
        RECT 4.400 118.640 187.040 120.040 ;
        RECT 3.990 89.440 187.040 118.640 ;
        RECT 4.400 88.040 187.040 89.440 ;
        RECT 3.990 82.640 187.040 88.040 ;
        RECT 3.990 81.240 186.640 82.640 ;
        RECT 3.990 72.440 187.040 81.240 ;
        RECT 4.400 71.040 187.040 72.440 ;
        RECT 3.990 31.640 187.040 71.040 ;
        RECT 3.990 30.240 186.640 31.640 ;
        RECT 3.990 10.715 187.040 30.240 ;
  END
END Systolic4x4_serial_io
END LIBRARY

