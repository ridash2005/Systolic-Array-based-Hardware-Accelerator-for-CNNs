* NGSPICE file created from Systolic4x4_serial_io.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

.subckt Systolic4x4_serial_io A_in_frame_sync A_in_serial_clk A_in_serial_data B_in_frame_sync
+ B_in_serial_clk B_in_serial_data C_out_frame_sync C_out_serial_clk C_out_serial_data
+ VGND VPWR clk done rst_n start
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer7 net22 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer481 _0415_ VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer492 _0416_ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkbuf_2
X_1270_ clknet_4_10_0_B_in_serial_clk _0217_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0985_ deser_B.kept_shift_reg\[104\] deser_B.kept_shift_reg\[105\] net845 VGND VGND
+ VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
X_1399_ clknet_2_1__leaf_clk _0343_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ deser_A.kept_shift_reg\[61\] deser_A.kept_shift_reg\[62\] net808 VGND VGND
+ VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_4
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1253_ clknet_4_12_0_B_in_serial_clk _0200_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1322_ clknet_4_4_0_B_in_serial_clk _0269_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1184_ clknet_4_4_0_A_in_serial_clk _0132_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0968_ deser_B.kept_shift_reg\[87\] deser_B.kept_shift_reg\[88\] net10 VGND VGND
+ VPWR VPWR _0283_ sky130_fd_sc_hd__mux2_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0899_ deser_B.kept_shift_reg\[18\] deser_B.kept_shift_reg\[19\] net11 VGND VGND
+ VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0822_ deser_A.kept_shift_reg\[113\] deser_A.kept_shift_reg\[114\] net735 VGND VGND
+ VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0753_ deser_A.kept_shift_reg\[44\] deser_A.kept_shift_reg\[45\] net730 VGND VGND
+ VPWR VPWR _0096_ sky130_fd_sc_hd__mux2_2
X_0684_ _0511_ _0501_ _0417_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__and3_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1236_ clknet_4_12_0_B_in_serial_clk _0184_ net15 VGND VGND VPWR VPWR deser_B.bit_idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1305_ clknet_4_0_0_B_in_serial_clk _0252_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_6_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_6_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1167_ clknet_4_15_0_A_in_serial_clk _0115_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
Xclone793 net24 VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__clkbuf_16
X_1098_ clknet_4_9_0_A_in_serial_clk _0047_ net14 VGND VGND VPWR VPWR deser_A.kept_bit_idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1021_ ser_C.bit_idx\[3\] ser_C.bit_idx\[4\] _0379_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__and3_1
X_0805_ deser_A.kept_shift_reg\[96\] deser_A.kept_shift_reg\[97\] net734 VGND VGND
+ VPWR VPWR _0148_ sky130_fd_sc_hd__mux2_4
X_0598_ _0451_ _0452_ systolic_inst.cycle_cnt\[10\] VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__mux2_1
X_0667_ net22 net1 VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__and2b_1
X_0736_ deser_A.kept_shift_reg\[27\] deser_A.kept_shift_reg\[28\] net17 VGND VGND
+ VPWR VPWR _0079_ sky130_fd_sc_hd__mux2_1
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1219_ clknet_4_1_0_A_in_serial_clk _0167_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer800 _0363_ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_14_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_45_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer17 _0363_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer28 net739 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_8
X_1004_ deser_B.kept_shift_reg\[123\] deser_B.kept_shift_reg\[124\] net27 VGND VGND
+ VPWR VPWR _0319_ sky130_fd_sc_hd__mux2_1
XFILLER_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0719_ deser_A.kept_shift_reg\[10\] deser_A.kept_shift_reg\[11\] net18 VGND VGND
+ VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_4
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput7 net7 VGND VGND VPWR VPWR C_out_frame_sync sky130_fd_sc_hd__buf_1
Xclkbuf_4_7_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_7_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer493 _0417_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_1
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer8 net22 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_8
XFILLER_47_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0984_ deser_B.kept_shift_reg\[103\] deser_B.kept_shift_reg\[104\] net47 VGND VGND
+ VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_15_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_15_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1398_ clknet_2_1__leaf_clk _0342_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1252_ clknet_4_13_0_B_in_serial_clk _0199_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1321_ clknet_4_1_0_B_in_serial_clk _0268_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1183_ clknet_4_6_0_A_in_serial_clk _0131_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0967_ deser_B.kept_shift_reg\[86\] deser_B.kept_shift_reg\[87\] net10 VGND VGND
+ VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
XFILLER_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0898_ deser_B.kept_shift_reg\[17\] deser_B.kept_shift_reg\[18\] net640 VGND VGND
+ VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0821_ deser_A.kept_shift_reg\[112\] deser_A.kept_shift_reg\[113\] net12 VGND VGND
+ VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
X_0752_ deser_A.kept_shift_reg\[43\] deser_A.kept_shift_reg\[44\] net728 VGND VGND
+ VPWR VPWR _0095_ sky130_fd_sc_hd__mux2_2
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ _0420_ net508 deser_A.bit_idx\[5\] deser_A.bit_idx\[6\] VGND VGND VPWR VPWR
+ _0511_ sky130_fd_sc_hd__a31o_1
X_1235_ clknet_4_13_0_B_in_serial_clk _0183_ net15 VGND VGND VPWR VPWR deser_B.bit_idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1304_ clknet_4_2_0_B_in_serial_clk _0251_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_1166_ clknet_4_15_0_A_in_serial_clk _0114_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1097_ clknet_4_10_0_A_in_serial_clk _0046_ net14 VGND VGND VPWR VPWR deser_A.kept_bit_idx\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1020_ ser_C.bit_idx\[3\] _0379_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__xor2_1
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0804_ deser_A.kept_shift_reg\[95\] deser_A.kept_shift_reg\[96\] net12 VGND VGND
+ VPWR VPWR _0147_ sky130_fd_sc_hd__mux2_1
X_0735_ deser_A.kept_shift_reg\[26\] deser_A.kept_shift_reg\[27\] net808 VGND VGND
+ VPWR VPWR _0078_ sky130_fd_sc_hd__mux2_4
X_0597_ systolic_inst.cycle_cnt\[9\] _0453_ _0452_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__o21a_1
X_0666_ net17 _0419_ net491 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux2_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1149_ clknet_4_7_0_A_in_serial_clk _0097_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_1218_ clknet_4_4_0_A_in_serial_clk _0166_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ deser_B.kept_shift_reg\[122\] deser_B.kept_shift_reg\[123\] net847 VGND VGND
+ VPWR VPWR _0318_ sky130_fd_sc_hd__mux2_1
Xrebuffer18 deser_B.receiving VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_8
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0718_ deser_A.kept_shift_reg\[9\] deser_A.kept_shift_reg\[10\] net25 VGND VGND VPWR
+ VPWR _0061_ sky130_fd_sc_hd__mux2_2
X_0649_ systolic_inst.cycle_cnt\[26\] _0483_ _0486_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__and3_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR C_out_serial_clk sky130_fd_sc_hd__buf_1
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer483 _0347_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer9 net24 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ deser_B.kept_shift_reg\[102\] deser_B.kept_shift_reg\[103\] net10 VGND VGND
+ VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1397_ clknet_2_1__leaf_clk _0341_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1320_ clknet_4_1_0_B_in_serial_clk _0267_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_1251_ clknet_4_13_0_B_in_serial_clk _0198_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1182_ clknet_4_6_0_A_in_serial_clk _0130_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0966_ deser_B.kept_shift_reg\[85\] deser_B.kept_shift_reg\[86\] net47 VGND VGND
+ VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
X_0897_ deser_B.kept_shift_reg\[16\] deser_B.kept_shift_reg\[17\] net11 VGND VGND
+ VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0820_ deser_A.kept_shift_reg\[111\] deser_A.kept_shift_reg\[112\] net730 VGND VGND
+ VPWR VPWR _0163_ sky130_fd_sc_hd__mux2_4
X_0751_ deser_A.kept_shift_reg\[42\] deser_A.kept_shift_reg\[43\] net12 VGND VGND
+ VPWR VPWR _0094_ sky130_fd_sc_hd__mux2_1
X_1303_ clknet_4_2_0_B_in_serial_clk _0250_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_0682_ _0501_ _0510_ _0509_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and3_1
XFILLER_64_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1234_ clknet_4_13_0_B_in_serial_clk _0182_ net15 VGND VGND VPWR VPWR deser_B.bit_idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1165_ clknet_4_15_0_A_in_serial_clk _0113_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_1096_ clknet_4_8_0_A_in_serial_clk _0045_ net14 VGND VGND VPWR VPWR deser_A.kept_bit_idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_0949_ deser_B.kept_shift_reg\[68\] deser_B.kept_shift_reg\[69\] net10 VGND VGND
+ VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
XFILLER_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0665_ _0499_ _0401_ _0498_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux2_1
X_0803_ deser_A.kept_shift_reg\[94\] deser_A.kept_shift_reg\[95\] net12 VGND VGND
+ VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_1
X_0734_ deser_A.kept_shift_reg\[25\] deser_A.kept_shift_reg\[26\] net740 VGND VGND
+ VPWR VPWR _0077_ sky130_fd_sc_hd__mux2_2
X_0596_ systolic_inst.cycle_cnt\[8\] _0428_ _0447_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__and3_1
X_1079_ clknet_2_3__leaf_clk _0028_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_1217_ clknet_4_4_0_A_in_serial_clk _0165_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1148_ clknet_4_7_0_A_in_serial_clk _0096_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer802 deser_A.receiving VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__buf_2
XFILLER_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_7 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1002_ deser_B.kept_shift_reg\[121\] deser_B.kept_shift_reg\[122\] net27 VGND VGND
+ VPWR VPWR _0317_ sky130_fd_sc_hd__mux2_1
Xrebuffer19 net34 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlymetal6s2s_1
X_0648_ systolic_inst.cycle_cnt\[26\] _0436_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__nand2_1
X_0717_ deser_A.kept_shift_reg\[8\] deser_A.kept_shift_reg\[9\] net23 VGND VGND VPWR
+ VPWR _0060_ sky130_fd_sc_hd__mux2_2
X_0579_ _0439_ _0440_ systolic_inst.cycle_cnt\[4\] VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_33_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput9 net9 VGND VGND VPWR VPWR done sky130_fd_sc_hd__buf_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer484 _0347_ VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0982_ deser_B.kept_shift_reg\[101\] deser_B.kept_shift_reg\[102\] net10 VGND VGND
+ VPWR VPWR _0297_ sky130_fd_sc_hd__mux2_1
XFILLER_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1396_ clknet_2_1__leaf_clk _0340_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ clknet_4_13_0_B_in_serial_clk _0197_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1181_ clknet_4_6_0_A_in_serial_clk _0129_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0965_ deser_B.kept_shift_reg\[84\] deser_B.kept_shift_reg\[85\] net10 VGND VGND
+ VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
X_0896_ deser_B.kept_shift_reg\[15\] deser_B.kept_shift_reg\[16\] net11 VGND VGND
+ VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
XFILLER_55_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1379_ clknet_2_2__leaf_clk _0004_ net5 VGND VGND VPWR VPWR systolic_inst.ce_local
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_2_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0681_ _0420_ _0415_ deser_A.bit_idx\[4\] deser_A.bit_idx\[5\] VGND VGND VPWR VPWR
+ _0510_ sky130_fd_sc_hd__a31o_1
X_0750_ deser_A.kept_shift_reg\[41\] deser_A.kept_shift_reg\[42\] net730 VGND VGND
+ VPWR VPWR _0093_ sky130_fd_sc_hd__mux2_4
X_1233_ clknet_4_13_0_B_in_serial_clk _0181_ net15 VGND VGND VPWR VPWR deser_B.bit_idx\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1302_ clknet_4_2_0_B_in_serial_clk _0249_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1164_ clknet_4_15_0_A_in_serial_clk _0112_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_1095_ clknet_4_10_0_A_in_serial_clk _0044_ net14 VGND VGND VPWR VPWR deser_A.bit_idx\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0948_ deser_B.kept_shift_reg\[67\] deser_B.kept_shift_reg\[68\] net10 VGND VGND
+ VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
XFILLER_20_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0879_ deser_B.kept_bit_idx\[7\] _0373_ _0371_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux2_4
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0802_ deser_A.kept_shift_reg\[93\] deser_A.kept_shift_reg\[94\] net730 VGND VGND
+ VPWR VPWR _0145_ sky130_fd_sc_hd__mux2_4
X_0664_ _0401_ _0435_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__nor2_1
X_0733_ deser_A.kept_shift_reg\[24\] deser_A.kept_shift_reg\[25\] net40 VGND VGND
+ VPWR VPWR _0076_ sky130_fd_sc_hd__mux2_1
X_0595_ _0435_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__nor2_1
X_1216_ clknet_4_4_0_A_in_serial_clk _0164_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_1078_ clknet_2_3__leaf_clk _0027_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1147_ clknet_4_7_0_A_in_serial_clk _0095_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_42_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_1_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_49_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ deser_B.kept_shift_reg\[120\] deser_B.kept_shift_reg\[121\] net847 VGND VGND
+ VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0578_ _0438_ _0440_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__and2_1
X_0647_ _0436_ _0485_ _0487_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__and3_1
X_0716_ deser_A.kept_shift_reg\[7\] deser_A.kept_shift_reg\[8\] net17 VGND VGND VPWR
+ VPWR _0059_ sky130_fd_sc_hd__mux2_1
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer485 deser_B.bit_idx\[0\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer474 deser_A.bit_idx\[0\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ deser_B.kept_shift_reg\[100\] deser_B.kept_shift_reg\[101\] net47 VGND VGND
+ VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1395_ clknet_2_1__leaf_clk _0339_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_2_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_58_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1180_ clknet_4_7_0_A_in_serial_clk _0128_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0964_ deser_B.kept_shift_reg\[83\] deser_B.kept_shift_reg\[84\] net47 VGND VGND
+ VPWR VPWR _0279_ sky130_fd_sc_hd__mux2_1
X_0895_ deser_B.kept_shift_reg\[14\] deser_B.kept_shift_reg\[15\] net640 VGND VGND
+ VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_4
X_1378_ clknet_4_8_0_A_in_serial_clk _0325_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0680_ deser_A.bit_idx\[5\] _0416_ _0420_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__nand3_1
X_1232_ clknet_4_13_0_B_in_serial_clk _0180_ net15 VGND VGND VPWR VPWR deser_B.bit_idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_10_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_10_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1301_ clknet_4_2_0_B_in_serial_clk _0248_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1163_ clknet_4_15_0_A_in_serial_clk _0111_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
Xclone753 net24 VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__buf_12
X_1094_ clknet_4_10_0_A_in_serial_clk _0043_ net14 VGND VGND VPWR VPWR deser_A.bit_idx\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_0947_ deser_B.kept_shift_reg\[66\] deser_B.kept_shift_reg\[67\] net10 VGND VGND
+ VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_1
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0878_ deser_B.kept_bit_idx\[7\] _0348_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__nand2_1
XFILLER_28_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_4
XFILLER_61_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0801_ deser_A.kept_shift_reg\[92\] deser_A.kept_shift_reg\[93\] net732 VGND VGND
+ VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_4
X_0663_ _0497_ _0400_ _0496_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_1
X_0594_ systolic_inst.cycle_cnt\[8\] systolic_inst.cycle_cnt\[9\] _0448_ VGND VGND
+ VPWR VPWR _0451_ sky130_fd_sc_hd__and3_1
X_0732_ deser_A.kept_shift_reg\[23\] deser_A.kept_shift_reg\[24\] net40 VGND VGND
+ VPWR VPWR _0075_ sky130_fd_sc_hd__mux2_1
X_1215_ clknet_4_4_0_A_in_serial_clk _0163_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_1146_ clknet_4_7_0_A_in_serial_clk _0094_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_1077_ clknet_2_1__leaf_clk _0026_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer804 deser_B.receiving VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_9 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1000_ deser_B.kept_shift_reg\[119\] deser_B.kept_shift_reg\[120\] net845 VGND VGND
+ VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0715_ deser_A.kept_shift_reg\[6\] deser_A.kept_shift_reg\[7\] net23 VGND VGND VPWR
+ VPWR _0058_ sky130_fd_sc_hd__mux2_1
X_0577_ _0435_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__nor2_1
X_0646_ _0483_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__nand2_1
X_1129_ clknet_4_12_0_A_in_serial_clk _0077_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0629_ _0472_ _0475_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__and2_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer475 deser_A.bit_idx\[0\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer486 net501 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0980_ deser_B.kept_shift_reg\[99\] deser_B.kept_shift_reg\[100\] net47 VGND VGND
+ VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_1
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1394_ clknet_2_1__leaf_clk _0338_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0894_ deser_B.kept_shift_reg\[13\] deser_B.kept_shift_reg\[14\] net11 VGND VGND
+ VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
X_0963_ deser_B.kept_shift_reg\[82\] deser_B.kept_shift_reg\[83\] net47 VGND VGND
+ VPWR VPWR _0278_ sky130_fd_sc_hd__mux2_1
X_1377_ clknet_4_13_0_B_in_serial_clk _0324_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1300_ clknet_4_2_0_B_in_serial_clk _0247_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_1162_ clknet_4_15_0_A_in_serial_clk _0110_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_1231_ clknet_4_2_0_A_in_serial_clk _0179_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1093_ clknet_4_10_0_A_in_serial_clk _0042_ net14 VGND VGND VPWR VPWR deser_A.bit_idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_0877_ _0371_ _0372_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__and2_1
X_0946_ deser_B.kept_shift_reg\[65\] deser_B.kept_shift_reg\[66\] net47 VGND VGND
+ VPWR VPWR _0261_ sky130_fd_sc_hd__mux2_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0800_ deser_A.kept_shift_reg\[91\] deser_A.kept_shift_reg\[92\] net735 VGND VGND
+ VPWR VPWR _0143_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_12_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0731_ deser_A.kept_shift_reg\[22\] deser_A.kept_shift_reg\[23\] net44 VGND VGND
+ VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_2
X_0662_ systolic_inst.cycle_cnt\[28\] systolic_inst.cycle_cnt\[29\] systolic_inst.cycle_cnt\[30\]
+ _0492_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__and4_1
X_0593_ systolic_inst.cycle_cnt\[8\] _0448_ _0450_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1145_ clknet_4_6_0_A_in_serial_clk _0093_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_1214_ clknet_4_5_0_A_in_serial_clk _0162_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[110\]
+ sky130_fd_sc_hd__dfrtp_1
Xrebuffer805 deser_B.receiving VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__buf_1
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1076_ clknet_2_1__leaf_clk _0025_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_0929_ deser_B.kept_shift_reg\[48\] deser_B.kept_shift_reg\[49\] net642 VGND VGND
+ VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_4
Xclkbuf_4_9_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_9_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0645_ systolic_inst.cycle_cnt\[24\] systolic_inst.cycle_cnt\[25\] VGND VGND VPWR
+ VPWR _0486_ sky130_fd_sc_hd__and2_1
XFILLER_30_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0714_ deser_A.kept_shift_reg\[5\] deser_A.kept_shift_reg\[6\] net24 VGND VGND VPWR
+ VPWR _0057_ sky130_fd_sc_hd__mux2_1
X_0576_ systolic_inst.cycle_cnt\[2\] systolic_inst.cycle_cnt\[3\] _0434_ VGND VGND
+ VPWR VPWR _0439_ sky130_fd_sc_hd__and3_1
XFILLER_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1059_ clknet_2_2__leaf_clk _0008_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1128_ clknet_4_12_0_A_in_serial_clk _0076_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0628_ _0435_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__nor2_1
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0559_ net6 systolic_inst.ce_local VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__nor2_1
XFILLER_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer487 deser_B.bit_idx\[2\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_42_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_39_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer476 net491 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_48_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1393_ clknet_2_0__leaf_clk _0337_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0893_ deser_B.kept_shift_reg\[12\] deser_B.kept_shift_reg\[13\] net640 VGND VGND
+ VPWR VPWR _0208_ sky130_fd_sc_hd__mux2_4
X_0962_ deser_B.kept_shift_reg\[81\] deser_B.kept_shift_reg\[82\] net10 VGND VGND
+ VPWR VPWR _0277_ sky130_fd_sc_hd__mux2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1376_ clknet_4_13_0_B_in_serial_clk _0323_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1161_ clknet_4_13_0_A_in_serial_clk _0109_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_1230_ clknet_4_8_0_A_in_serial_clk _0178_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1092_ clknet_4_10_0_A_in_serial_clk _0041_ net14 VGND VGND VPWR VPWR deser_A.bit_idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0876_ deser_B.kept_bit_idx\[6\] _0348_ net43 VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a21o_1
X_0945_ deser_B.kept_shift_reg\[64\] deser_B.kept_shift_reg\[65\] net10 VGND VGND
+ VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1359_ clknet_4_5_0_B_in_serial_clk _0306_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload2 clknet_2_3__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xload_slew14 net15 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_29_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0661_ _0400_ _0435_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_12_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0730_ deser_A.kept_shift_reg\[21\] deser_A.kept_shift_reg\[22\] net740 VGND VGND
+ VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_2
X_0592_ systolic_inst.cycle_cnt\[8\] _0436_ _0448_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1213_ clknet_4_5_0_A_in_serial_clk _0161_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1075_ clknet_2_1__leaf_clk _0024_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1144_ clknet_4_6_0_A_in_serial_clk _0092_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0859_ _0426_ deser_B.kept_bit_idx\[0\] deser_B.kept_bit_idx\[1\] VGND VGND VPWR
+ VPWR _0360_ sky130_fd_sc_hd__a21oi_2
X_0928_ deser_B.kept_shift_reg\[47\] deser_B.kept_shift_reg\[48\] net11 VGND VGND
+ VPWR VPWR _0243_ sky130_fd_sc_hd__mux2_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0644_ systolic_inst.cycle_cnt\[24\] _0470_ _0482_ systolic_inst.cycle_cnt\[25\]
+ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a31o_1
X_0713_ deser_A.kept_shift_reg\[4\] deser_A.kept_shift_reg\[5\] net17 VGND VGND VPWR
+ VPWR _0056_ sky130_fd_sc_hd__mux2_1
X_0575_ systolic_inst.cycle_cnt\[2\] _0428_ _0433_ systolic_inst.cycle_cnt\[3\] VGND
+ VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_27_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1058_ clknet_2_2__leaf_clk _0007_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_11_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1127_ clknet_4_12_0_A_in_serial_clk _0075_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xrebuffer625 net644 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_8
XFILLER_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0558_ _0424_ _0425_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__nor2_1
X_0627_ _0448_ _0464_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__and3_1
XFILLER_38_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer488 deser_B.bit_idx\[2\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer477 deser_A.bit_idx\[2\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_59_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1392_ clknet_2_0__leaf_clk _0002_ net5 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_65_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0961_ deser_B.kept_shift_reg\[80\] deser_B.kept_shift_reg\[81\] net47 VGND VGND
+ VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
XFILLER_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0892_ deser_B.kept_shift_reg\[11\] deser_B.kept_shift_reg\[12\] net11 VGND VGND
+ VPWR VPWR _0207_ sky130_fd_sc_hd__mux2_1
X_1375_ clknet_4_7_0_B_in_serial_clk _0322_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1160_ clknet_4_13_0_A_in_serial_clk _0108_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_1091_ clknet_4_10_0_A_in_serial_clk _0040_ net14 VGND VGND VPWR VPWR deser_A.bit_idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclone712 net731 VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__clkbuf_16
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0944_ deser_B.kept_shift_reg\[63\] deser_B.kept_shift_reg\[64\] net47 VGND VGND
+ VPWR VPWR _0259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0875_ deser_B.kept_bit_idx\[6\] _0368_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__nand2_1
Xclkload20 clknet_4_6_0_B_in_serial_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__inv_6
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1358_ clknet_4_5_0_B_in_serial_clk _0305_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1289_ clknet_4_11_0_B_in_serial_clk _0236_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload3 clknet_4_1_0_A_in_serial_clk VGND VGND VPWR VPWR clkload3/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_21_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xload_slew15 net5 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_16
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0660_ _0494_ _0495_ _0496_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__a21oi_1
X_0591_ _0436_ _0445_ _0449_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__and3_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1212_ clknet_4_5_0_A_in_serial_clk _0160_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1074_ clknet_2_1__leaf_clk _0023_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1143_ clknet_4_3_0_A_in_serial_clk _0091_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_0927_ deser_B.kept_shift_reg\[46\] deser_B.kept_shift_reg\[47\] net11 VGND VGND
+ VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_1
X_0858_ net845 _0425_ deser_B.kept_bit_idx\[0\] VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_4
X_0789_ deser_A.kept_shift_reg\[80\] deser_A.kept_shift_reg\[81\] net732 VGND VGND
+ VPWR VPWR _0132_ sky130_fd_sc_hd__mux2_4
XFILLER_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0574_ _0434_ _0437_ systolic_inst.cycle_cnt\[2\] VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__mux2_1
X_0643_ systolic_inst.cycle_cnt\[24\] _0483_ _0484_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a21oi_1
X_0712_ deser_A.kept_shift_reg\[3\] deser_A.kept_shift_reg\[4\] net17 VGND VGND VPWR
+ VPWR _0055_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1126_ clknet_4_12_0_A_in_serial_clk _0074_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1057_ clknet_2_2__leaf_clk _0006_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0557_ net3 net34 VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or2_4
X_0626_ systolic_inst.cycle_cnt\[16\] systolic_inst.cycle_cnt\[17\] systolic_inst.cycle_cnt\[18\]
+ systolic_inst.cycle_cnt\[19\] VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1109_ clknet_4_9_0_A_in_serial_clk _0057_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer489 deser_B.bit_idx\[1\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer478 deser_A.bit_idx\[1\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_59_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1391_ clknet_4_14_0_B_in_serial_clk _0336_ net15 VGND VGND VPWR VPWR deser_B.kept_receiving
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0609_ _0460_ _0461_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__nor2_1
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0960_ deser_B.kept_shift_reg\[79\] deser_B.kept_shift_reg\[80\] net10 VGND VGND
+ VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
X_0891_ deser_B.kept_shift_reg\[10\] deser_B.kept_shift_reg\[11\] net643 VGND VGND
+ VPWR VPWR _0206_ sky130_fd_sc_hd__mux2_4
X_1374_ clknet_4_13_0_B_in_serial_clk _0321_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone724 net739 VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__clkbuf_16
XFILLER_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ clknet_4_8_0_A_in_serial_clk _0039_ net14 VGND VGND VPWR VPWR deser_A.bit_idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_0874_ net45 _0369_ _0370_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__and3_1
X_0943_ deser_B.kept_shift_reg\[62\] deser_B.kept_shift_reg\[63\] net47 VGND VGND
+ VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
Xclkload10 clknet_4_11_0_A_in_serial_clk VGND VGND VPWR VPWR clkload10/X sky130_fd_sc_hd__clkbuf_8
Xclkload21 clknet_4_7_0_B_in_serial_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__clkinvlp_4
X_1357_ clknet_4_5_0_B_in_serial_clk _0304_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1288_ clknet_4_11_0_B_in_serial_clk _0235_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload4 clknet_4_3_0_A_in_serial_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_21_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0590_ _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__inv_2
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1211_ clknet_4_5_0_A_in_serial_clk _0159_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_1142_ clknet_4_3_0_A_in_serial_clk _0090_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1073_ clknet_2_1__leaf_clk _0022_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_0857_ _0424_ _0359_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__or2_4
X_0926_ deser_B.kept_shift_reg\[45\] deser_B.kept_shift_reg\[46\] net642 VGND VGND
+ VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_4
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0788_ deser_A.kept_shift_reg\[79\] deser_A.kept_shift_reg\[80\] net730 VGND VGND
+ VPWR VPWR _0131_ sky130_fd_sc_hd__mux2_4
XFILLER_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0711_ deser_A.kept_shift_reg\[2\] deser_A.kept_shift_reg\[3\] net17 VGND VGND VPWR
+ VPWR _0054_ sky130_fd_sc_hd__mux2_1
X_0573_ _0432_ _0437_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__and2_1
X_0642_ systolic_inst.cycle_cnt\[24\] _0483_ _0436_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1125_ clknet_4_12_0_A_in_serial_clk _0073_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_1056_ clknet_2_2__leaf_clk _0005_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0909_ deser_B.kept_shift_reg\[28\] deser_B.kept_shift_reg\[29\] net642 VGND VGND
+ VPWR VPWR _0224_ sky130_fd_sc_hd__mux2_4
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSystolic4x4_serial_io_16 VGND VGND VPWR VPWR Systolic4x4_serial_io_16/HI C_out_serial_data
+ sky130_fd_sc_hd__conb_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_4_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_4_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0625_ systolic_inst.cycle_cnt\[16\] systolic_inst.cycle_cnt\[17\] systolic_inst.cycle_cnt\[18\]
+ _0470_ systolic_inst.cycle_cnt\[19\] VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__a41o_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0556_ net3 net38 VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__nor2_8
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1108_ clknet_4_8_0_A_in_serial_clk _0056_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1039_ ser_C.kept_bit_idx\[0\] net7 ser_C.kept_bit_idx\[1\] ser_C.kept_bit_idx\[2\]
+ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__a31o_1
XFILLER_42_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer479 net494 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_59_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1390_ clknet_2_0__leaf_clk _0335_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0608_ systolic_inst.cycle_cnt\[12\] systolic_inst.cycle_cnt\[13\] _0448_ _0455_
+ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_56_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ systolic_inst.cycle_cnt\[4\] systolic_inst.cycle_cnt\[5\] systolic_inst.cycle_cnt\[6\]
+ systolic_inst.cycle_cnt\[7\] VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_64_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_12_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0890_ deser_B.kept_shift_reg\[9\] deser_B.kept_shift_reg\[10\] net10 VGND VGND VPWR
+ VPWR _0205_ sky130_fd_sc_hd__mux2_1
X_1373_ clknet_4_7_0_B_in_serial_clk _0320_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_5_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone714 net731 VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__buf_12
XFILLER_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0873_ deser_B.kept_bit_idx\[3\] deser_B.kept_bit_idx\[4\] _0426_ _0362_ deser_B.kept_bit_idx\[5\]
+ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a41o_1
Xclkload22 clknet_4_8_0_B_in_serial_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__clkinvlp_4
X_0942_ deser_B.kept_shift_reg\[61\] deser_B.kept_shift_reg\[62\] net47 VGND VGND
+ VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
Xclkload11 clknet_4_12_0_A_in_serial_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__bufinv_16
X_1356_ clknet_4_5_0_B_in_serial_clk _0303_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1287_ clknet_4_11_0_B_in_serial_clk _0234_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload5 clknet_4_4_0_A_in_serial_clk VGND VGND VPWR VPWR clkload5/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_21_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_A_in_serial_clk A_in_serial_clk VGND VGND VPWR VPWR clknet_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1210_ clknet_4_5_0_A_in_serial_clk _0158_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_1072_ clknet_2_1__leaf_clk _0021_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1141_ clknet_4_3_0_A_in_serial_clk _0089_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_13_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0856_ _0348_ _0423_ deser_B.bit_idx\[7\] VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__and3_1
X_0925_ deser_B.kept_shift_reg\[44\] deser_B.kept_shift_reg\[45\] net11 VGND VGND
+ VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
X_0787_ deser_A.kept_shift_reg\[78\] deser_A.kept_shift_reg\[79\] net808 VGND VGND
+ VPWR VPWR _0130_ sky130_fd_sc_hd__mux2_4
X_1339_ clknet_4_7_0_B_in_serial_clk _0286_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0641_ systolic_inst.ce_local _0447_ _0464_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__and4_1
X_0710_ deser_A.kept_shift_reg\[1\] deser_A.kept_shift_reg\[2\] net17 VGND VGND VPWR
+ VPWR _0053_ sky130_fd_sc_hd__mux2_1
X_0572_ _0434_ _0435_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__nor2_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1124_ clknet_4_12_0_A_in_serial_clk _0072_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_1055_ ser_C.kept_bit_idx\[9\] _0397_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__xnor2_1
Xrebuffer628 net821 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_31_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0839_ net37 net3 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__nand2b_4
X_0908_ deser_B.kept_shift_reg\[27\] deser_B.kept_shift_reg\[28\] net11 VGND VGND
+ VPWR VPWR _0223_ sky130_fd_sc_hd__mux2_1
XFILLER_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0624_ _0468_ _0469_ systolic_inst.cycle_cnt\[18\] VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__mux2_1
X_0555_ _0423_ deser_B.bit_idx\[7\] VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ clknet_4_8_0_A_in_serial_clk _0055_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1038_ ser_C.kept_bit_idx\[0\] net7 ser_C.kept_bit_idx\[1\] ser_C.kept_bit_idx\[2\]
+ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_59_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0538_ systolic_inst.cycle_cnt\[8\] systolic_inst.cycle_cnt\[9\] systolic_inst.cycle_cnt\[10\]
+ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__or3_1
X_0607_ systolic_inst.cycle_cnt\[13\] _0436_ _0456_ systolic_inst.cycle_cnt\[12\]
+ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_56_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1372_ clknet_4_7_0_B_in_serial_clk _0319_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_63_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0941_ deser_B.kept_shift_reg\[60\] deser_B.kept_shift_reg\[61\] net47 VGND VGND
+ VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
X_0872_ net42 VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__inv_2
XFILLER_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload23 clknet_4_9_0_B_in_serial_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_9_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload12 clknet_4_13_0_A_in_serial_clk VGND VGND VPWR VPWR clkload12/X sky130_fd_sc_hd__clkbuf_4
X_1355_ clknet_4_5_0_B_in_serial_clk _0302_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1286_ clknet_4_11_0_B_in_serial_clk _0233_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload6 clknet_4_6_0_A_in_serial_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_2
XFILLER_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ clknet_2_1__leaf_clk _0020_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ clknet_4_3_0_A_in_serial_clk _0088_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ deser_B.kept_shift_reg\[43\] deser_B.kept_shift_reg\[44\] net643 VGND VGND
+ VPWR VPWR _0239_ sky130_fd_sc_hd__mux2_4
X_0855_ _0423_ _0358_ net45 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__and3_1
X_0786_ deser_A.kept_shift_reg\[77\] deser_A.kept_shift_reg\[78\] net40 VGND VGND
+ VPWR VPWR _0129_ sky130_fd_sc_hd__mux2_1
X_1338_ clknet_4_6_0_B_in_serial_clk _0285_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_1269_ clknet_4_10_0_B_in_serial_clk _0216_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0571_ systolic_inst.ce_local net6 VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__nand2b_4
X_0640_ systolic_inst.cycle_cnt\[23\] _0473_ _0479_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and3_1
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1123_ clknet_4_14_0_A_in_serial_clk _0071_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1054_ _0397_ _0398_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__and2_1
Xrebuffer629 deser_B.receiving VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__buf_2
X_0907_ deser_B.kept_shift_reg\[26\] deser_B.kept_shift_reg\[27\] net11 VGND VGND
+ VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0838_ net34 net3 VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__and2b_1
X_0769_ deser_A.kept_shift_reg\[60\] deser_A.kept_shift_reg\[61\] net40 VGND VGND
+ VPWR VPWR _0112_ sky130_fd_sc_hd__mux2_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0554_ _0422_ deser_B.bit_idx\[5\] deser_B.bit_idx\[6\] net34 VGND VGND VPWR VPWR
+ _0423_ sky130_fd_sc_hd__nand4_4
X_0623_ _0469_ _0471_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__and2_1
X_1106_ clknet_4_8_0_A_in_serial_clk _0054_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1037_ ser_C.kept_bit_idx\[1\] _0387_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0537_ systolic_inst.cycle_cnt\[1\] systolic_inst.cycle_cnt\[2\] systolic_inst.cycle_cnt\[3\]
+ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__o21a_1
X_0606_ _0459_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1371_ clknet_4_7_0_B_in_serial_clk _0318_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone716 net733 VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__buf_12
X_0940_ deser_B.kept_shift_reg\[59\] deser_B.kept_shift_reg\[60\] net47 VGND VGND
+ VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0871_ deser_B.kept_bit_idx\[3\] deser_B.kept_bit_idx\[4\] _0363_ deser_B.kept_bit_idx\[5\]
+ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__and4_1
Xclkload24 clknet_4_10_0_B_in_serial_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__bufinv_16
Xclkload13 clknet_4_14_0_A_in_serial_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinv_2
X_1354_ clknet_4_5_0_B_in_serial_clk _0301_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1285_ clknet_4_9_0_B_in_serial_clk _0232_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload7 clknet_4_8_0_A_in_serial_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinv_2
XFILLER_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ clknet_2_0__leaf_clk _0019_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0854_ _0426_ _0422_ deser_B.bit_idx\[5\] deser_B.bit_idx\[6\] VGND VGND VPWR VPWR
+ _0358_ sky130_fd_sc_hd__a31o_1
X_0923_ deser_B.kept_shift_reg\[42\] deser_B.kept_shift_reg\[43\] net640 VGND VGND
+ VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0785_ deser_A.kept_shift_reg\[76\] deser_A.kept_shift_reg\[77\] net18 VGND VGND
+ VPWR VPWR _0128_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1337_ clknet_4_12_0_B_in_serial_clk _0284_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_1268_ clknet_4_10_0_B_in_serial_clk _0215_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1199_ clknet_4_1_0_A_in_serial_clk _0147_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0570_ systolic_inst.ce_local net6 VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_40_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1122_ clknet_4_14_0_A_in_serial_clk _0070_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1053_ ser_C.kept_bit_idx\[8\] _0395_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or2_1
X_0837_ net845 _0425_ deser_B.bit_idx\[0\] VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_4
X_0906_ deser_B.kept_shift_reg\[25\] deser_B.kept_shift_reg\[26\] net11 VGND VGND
+ VPWR VPWR _0221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0768_ deser_A.kept_shift_reg\[59\] deser_A.kept_shift_reg\[60\] net40 VGND VGND
+ VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_1
X_0699_ _0520_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
XFILLER_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0553_ deser_B.bit_idx\[4\] _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__and2_4
X_0622_ systolic_inst.cycle_cnt\[16\] _0470_ systolic_inst.cycle_cnt\[17\] VGND VGND
+ VPWR VPWR _0471_ sky130_fd_sc_hd__a21o_1
X_1105_ clknet_4_8_0_A_in_serial_clk _0053_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1036_ _0387_ _0388_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0536_ systolic_inst.cycle_cnt\[28\] systolic_inst.cycle_cnt\[29\] systolic_inst.cycle_cnt\[30\]
+ systolic_inst.cycle_cnt\[31\] VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or4_1
X_0605_ _0458_ systolic_inst.cycle_cnt\[12\] _0456_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1019_ _0379_ _0380_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__nor2_1
XFILLER_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ clknet_4_7_0_B_in_serial_clk _0317_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0870_ _0367_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__inv_2
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload25 clknet_4_11_0_B_in_serial_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__clkinv_2
Xclkload14 clknet_4_15_0_A_in_serial_clk VGND VGND VPWR VPWR clkload14/X sky130_fd_sc_hd__clkbuf_4
X_1353_ clknet_4_5_0_B_in_serial_clk _0300_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1284_ clknet_4_9_0_B_in_serial_clk _0231_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0999_ deser_B.kept_shift_reg\[118\] deser_B.kept_shift_reg\[119\] net847 VGND VGND
+ VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_1
Xclkload8 clknet_4_9_0_A_in_serial_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__bufinv_16
XFILLER_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0853_ _0356_ _0357_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__nor2_1
XFILLER_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0922_ deser_B.kept_shift_reg\[41\] deser_B.kept_shift_reg\[42\] net640 VGND VGND
+ VPWR VPWR _0237_ sky130_fd_sc_hd__mux2_4
X_0784_ deser_A.kept_shift_reg\[75\] deser_A.kept_shift_reg\[76\] net18 VGND VGND
+ VPWR VPWR _0127_ sky130_fd_sc_hd__mux2_4
X_1336_ clknet_4_12_0_B_in_serial_clk _0283_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_1267_ clknet_4_10_0_B_in_serial_clk _0214_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1198_ clknet_4_1_0_A_in_serial_clk _0146_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 A_in_frame_sync VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_0_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_0_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_34_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1121_ clknet_4_14_0_A_in_serial_clk _0069_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1052_ ser_C.kept_bit_idx\[8\] _0395_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__nand2_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0905_ deser_B.kept_shift_reg\[24\] deser_B.kept_shift_reg\[25\] net642 VGND VGND
+ VPWR VPWR _0220_ sky130_fd_sc_hd__mux2_4
X_0767_ deser_A.kept_shift_reg\[58\] deser_A.kept_shift_reg\[59\] net40 VGND VGND
+ VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0836_ deser_A.kept_shift_reg\[127\] net2 net647 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux2_4
XFILLER_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0698_ deser_A.kept_bit_idx\[3\] deser_A.kept_bit_idx\[4\] net28 _0519_ VGND VGND
+ VPWR VPWR _0520_ sky130_fd_sc_hd__a31o_1
X_1319_ clknet_4_1_0_B_in_serial_clk _0266_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0621_ _0428_ _0447_ _0464_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__and3_1
X_0552_ deser_B.bit_idx\[0\] deser_B.bit_idx\[1\] deser_B.bit_idx\[3\] deser_B.bit_idx\[2\]
+ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__and4_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1104_ clknet_4_10_0_A_in_serial_clk _0000_ net14 VGND VGND VPWR VPWR deser_A.receiving
+ sky130_fd_sc_hd__dfrtp_4
X_1035_ ser_C.kept_bit_idx\[0\] net7 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or2_1
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0819_ deser_A.kept_shift_reg\[110\] deser_A.kept_shift_reg\[111\] net730 VGND VGND
+ VPWR VPWR _0162_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_42_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0604_ systolic_inst.cycle_cnt\[12\] _0436_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0535_ systolic_inst.cycle_cnt\[20\] systolic_inst.cycle_cnt\[21\] systolic_inst.cycle_cnt\[22\]
+ systolic_inst.cycle_cnt\[23\] VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or4_1
XFILLER_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1018_ ser_C.bit_idx\[2\] _0377_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone718 net733 VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__buf_12
XFILLER_57_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload26 clknet_4_12_0_B_in_serial_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__inv_6
Xclkload15 clknet_4_0_0_B_in_serial_clk VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__bufinv_16
XPHY_EDGE_ROW_41_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1352_ clknet_4_5_0_B_in_serial_clk _0299_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_50_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1283_ clknet_4_9_0_B_in_serial_clk _0230_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ deser_B.kept_shift_reg\[117\] deser_B.kept_shift_reg\[118\] net19 VGND VGND
+ VPWR VPWR _0313_ sky130_fd_sc_hd__mux2_1
Xclkload9 clknet_4_10_0_A_in_serial_clk VGND VGND VPWR VPWR clkload9/X sky130_fd_sc_hd__clkbuf_8
XFILLER_54_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0921_ deser_B.kept_shift_reg\[40\] deser_B.kept_shift_reg\[41\] net643 VGND VGND
+ VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_4
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0852_ deser_B.bit_idx\[5\] net811 _0426_ net499 VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a31o_1
XFILLER_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0783_ deser_A.kept_shift_reg\[74\] deser_A.kept_shift_reg\[75\] net740 VGND VGND
+ VPWR VPWR _0126_ sky130_fd_sc_hd__mux2_2
X_1335_ clknet_4_9_0_B_in_serial_clk _0282_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_1266_ clknet_4_10_0_B_in_serial_clk _0213_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 A_in_serial_data VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
X_1197_ clknet_4_1_0_A_in_serial_clk _0145_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1120_ clknet_4_14_0_A_in_serial_clk _0068_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1051_ _0395_ _0396_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__nor2_1
X_0904_ deser_B.kept_shift_reg\[23\] deser_B.kept_shift_reg\[24\] net642 VGND VGND
+ VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_4
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0766_ deser_A.kept_shift_reg\[57\] deser_A.kept_shift_reg\[58\] net40 VGND VGND
+ VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_1
X_0835_ deser_A.kept_shift_reg\[126\] deser_A.kept_shift_reg\[127\] net728 VGND VGND
+ VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_4
X_0697_ deser_A.kept_bit_idx\[4\] _0501_ net28 deser_A.kept_bit_idx\[3\] VGND VGND
+ VPWR VPWR _0519_ sky130_fd_sc_hd__a22oi_2
X_1318_ clknet_4_1_0_B_in_serial_clk _0265_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[69\]
+ sky130_fd_sc_hd__dfrtp_1
X_1249_ clknet_4_11_0_A_in_serial_clk _0196_ net14 VGND VGND VPWR VPWR deser_A.kept_receiving
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0620_ systolic_inst.cycle_cnt\[16\] systolic_inst.cycle_cnt\[17\] _0465_ _0435_
+ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__a31oi_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0551_ _0418_ _0419_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__nor2_1
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1103_ clknet_4_11_0_A_in_serial_clk _0052_ net14 VGND VGND VPWR VPWR deser_A.kept_bit_idx\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1034_ ser_C.kept_bit_idx\[0\] net7 VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__nand2_1
XFILLER_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0749_ deser_A.kept_shift_reg\[40\] deser_A.kept_shift_reg\[41\] net734 VGND VGND
+ VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_4
X_0818_ deser_A.kept_shift_reg\[109\] deser_A.kept_shift_reg\[110\] net12 VGND VGND
+ VPWR VPWR _0161_ sky130_fd_sc_hd__mux2_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0534_ systolic_inst.cycle_cnt\[24\] systolic_inst.cycle_cnt\[25\] systolic_inst.cycle_cnt\[26\]
+ systolic_inst.cycle_cnt\[27\] VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or4_1
X_0603_ _0436_ _0454_ _0457_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_7_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_7_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_64_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ ser_C.bit_idx\[0\] ser_C.bit_idx\[1\] ser_C.bit_idx\[2\] net7 VGND VGND VPWR
+ VPWR _0379_ sky130_fd_sc_hd__and4_1
XFILLER_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone719 net733 VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__clkbuf_16
XFILLER_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_15_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_15_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
Xclkload27 clknet_4_13_0_B_in_serial_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__bufinv_16
Xclkload16 clknet_4_1_0_B_in_serial_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_23_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1351_ clknet_4_5_0_B_in_serial_clk _0298_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_1282_ clknet_4_9_0_B_in_serial_clk _0229_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0997_ deser_B.kept_shift_reg\[116\] deser_B.kept_shift_reg\[117\] net847 VGND VGND
+ VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
XFILLER_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_8_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0920_ deser_B.kept_shift_reg\[39\] deser_B.kept_shift_reg\[40\] net11 VGND VGND
+ VPWR VPWR _0235_ sky130_fd_sc_hd__mux2_1
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_23_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0851_ net811 _0426_ deser_B.bit_idx\[5\] VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a21oi_1
X_0782_ deser_A.kept_shift_reg\[73\] deser_A.kept_shift_reg\[74\] net44 VGND VGND
+ VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_2
X_1334_ clknet_4_9_0_B_in_serial_clk _0281_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1265_ clknet_4_10_0_B_in_serial_clk _0212_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 B_in_frame_sync VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1196_ clknet_4_0_0_A_in_serial_clk _0144_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1050_ ser_C.kept_bit_idx\[6\] _0393_ ser_C.kept_bit_idx\[7\] VGND VGND VPWR VPWR
+ _0396_ sky130_fd_sc_hd__a21oi_1
X_0903_ deser_B.kept_shift_reg\[22\] deser_B.kept_shift_reg\[23\] net11 VGND VGND
+ VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0834_ deser_A.kept_shift_reg\[125\] deser_A.kept_shift_reg\[126\] net735 VGND VGND
+ VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_4
XFILLER_21_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0765_ deser_A.kept_shift_reg\[56\] deser_A.kept_shift_reg\[57\] net769 VGND VGND
+ VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_4
X_0696_ deser_A.kept_bit_idx\[3\] net28 _0518_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1248_ clknet_4_14_0_B_in_serial_clk _0001_ net15 VGND VGND VPWR VPWR deser_B.receiving
+ sky130_fd_sc_hd__dfrtp_4
X_1317_ clknet_4_1_0_B_in_serial_clk _0264_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1179_ clknet_4_6_0_A_in_serial_clk _0127_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap10 net11 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_12
XFILLER_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0550_ deser_A.receiving net1 VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__or2_4
X_1102_ clknet_4_11_0_A_in_serial_clk _0051_ net14 VGND VGND VPWR VPWR deser_A.kept_bit_idx\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1033_ _0404_ _0424_ net45 VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__o21ai_1
X_0817_ deser_A.kept_shift_reg\[108\] deser_A.kept_shift_reg\[109\] net728 VGND VGND
+ VPWR VPWR _0160_ sky130_fd_sc_hd__mux2_2
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0679_ _0508_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_10_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0748_ deser_A.kept_shift_reg\[39\] deser_A.kept_shift_reg\[40\] net12 VGND VGND
+ VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_1
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0533_ deser_B.kept_receiving VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__inv_2
X_0602_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1016_ _0377_ _0378_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone31 net11 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_16
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer794 _0514_ VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload28 clknet_4_14_0_B_in_serial_clk VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__inv_6
Xclkload17 clknet_4_2_0_B_in_serial_clk VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_23_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1350_ clknet_4_4_0_B_in_serial_clk _0297_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_1281_ clknet_4_3_0_B_in_serial_clk _0228_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0996_ deser_B.kept_shift_reg\[115\] deser_B.kept_shift_reg\[116\] net27 VGND VGND
+ VPWR VPWR _0311_ sky130_fd_sc_hd__mux2_1
XFILLER_8_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ _0355_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__inv_2
X_1402_ clknet_2_1__leaf_clk _0346_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_0781_ deser_A.kept_shift_reg\[72\] deser_A.kept_shift_reg\[73\] net740 VGND VGND
+ VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_2
Xinput4 B_in_serial_data VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_1333_ clknet_4_12_0_B_in_serial_clk _0280_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_1264_ clknet_4_11_0_B_in_serial_clk _0211_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1195_ clknet_4_0_0_A_in_serial_clk _0143_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_0979_ deser_B.kept_shift_reg\[98\] deser_B.kept_shift_reg\[99\] net10 VGND VGND
+ VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0902_ deser_B.kept_shift_reg\[21\] deser_B.kept_shift_reg\[22\] net11 VGND VGND
+ VPWR VPWR _0217_ sky130_fd_sc_hd__mux2_1
X_0833_ deser_A.kept_shift_reg\[124\] deser_A.kept_shift_reg\[125\] net12 VGND VGND
+ VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_47_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0764_ deser_A.kept_shift_reg\[55\] deser_A.kept_shift_reg\[56\] net40 VGND VGND
+ VPWR VPWR _0107_ sky130_fd_sc_hd__mux2_1
X_0695_ deser_A.kept_bit_idx\[3\] _0501_ net30 VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1247_ clknet_4_14_0_B_in_serial_clk _0195_ net15 VGND VGND VPWR VPWR deser_B.kept_bit_idx\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1316_ clknet_4_0_0_B_in_serial_clk _0263_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_1178_ clknet_4_12_0_A_in_serial_clk _0126_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_65_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap11 net645 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_12
XFILLER_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1032_ ser_C.bit_idx\[9\] _0385_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__xor2_1
X_1101_ clknet_4_11_0_A_in_serial_clk _0050_ net14 VGND VGND VPWR VPWR deser_A.kept_bit_idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_0816_ deser_A.kept_shift_reg\[107\] deser_A.kept_shift_reg\[108\] net728 VGND VGND
+ VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_2
X_0747_ deser_A.kept_shift_reg\[38\] deser_A.kept_shift_reg\[39\] net12 VGND VGND
+ VPWR VPWR _0090_ sky130_fd_sc_hd__mux2_1
X_0678_ deser_A.bit_idx\[4\] _0507_ _0506_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux2_4
XFILLER_52_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0601_ _0448_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__and2_1
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0532_ deser_A.kept_receiving VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1015_ ser_C.bit_idx\[0\] net7 ser_C.bit_idx\[1\] VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21oi_1
X_1917_ clknet_2_0__leaf_clk VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_4_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer795 _0422_ VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload29 clknet_4_15_0_B_in_serial_clk VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__clkinv_4
Xclkload18 clknet_4_3_0_B_in_serial_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__inv_6
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1280_ clknet_4_3_0_B_in_serial_clk _0227_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ deser_B.kept_shift_reg\[114\] deser_B.kept_shift_reg\[115\] net27 VGND VGND
+ VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_1
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0780_ deser_A.kept_shift_reg\[71\] deser_A.kept_shift_reg\[72\] net769 VGND VGND
+ VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_4
X_1401_ clknet_2_1__leaf_clk _0345_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput5 rst_n VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_12
X_1332_ clknet_4_9_0_B_in_serial_clk _0279_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_1263_ clknet_4_11_0_B_in_serial_clk _0210_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1194_ clknet_4_0_0_A_in_serial_clk _0142_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0978_ deser_B.kept_shift_reg\[97\] deser_B.kept_shift_reg\[98\] net10 VGND VGND
+ VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0901_ deser_B.kept_shift_reg\[20\] deser_B.kept_shift_reg\[21\] net643 VGND VGND
+ VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_4
X_0763_ deser_A.kept_shift_reg\[54\] deser_A.kept_shift_reg\[55\] net809 VGND VGND
+ VPWR VPWR _0106_ sky130_fd_sc_hd__mux2_4
X_0832_ deser_A.kept_shift_reg\[123\] deser_A.kept_shift_reg\[124\] net735 VGND VGND
+ VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_4
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1315_ clknet_4_0_0_B_in_serial_clk _0262_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_0694_ net29 _0517_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__nor2_1
XFILLER_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1246_ clknet_4_14_0_B_in_serial_clk _0194_ net15 VGND VGND VPWR VPWR deser_B.kept_bit_idx\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1177_ clknet_4_13_0_A_in_serial_clk _0125_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap12 net729 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_53_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1031_ _0385_ _0386_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__nor2_1
X_1100_ clknet_4_11_0_A_in_serial_clk _0049_ net14 VGND VGND VPWR VPWR deser_A.kept_bit_idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_0815_ deser_A.kept_shift_reg\[106\] deser_A.kept_shift_reg\[107\] net647 VGND VGND
+ VPWR VPWR _0158_ sky130_fd_sc_hd__mux2_4
X_0746_ deser_A.kept_shift_reg\[37\] deser_A.kept_shift_reg\[38\] net728 VGND VGND
+ VPWR VPWR _0089_ sky130_fd_sc_hd__mux2_4
X_0677_ deser_A.bit_idx\[4\] _0501_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__nand2_1
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1229_ clknet_4_2_0_A_in_serial_clk _0177_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0600_ systolic_inst.cycle_cnt\[8\] systolic_inst.cycle_cnt\[9\] systolic_inst.cycle_cnt\[10\]
+ systolic_inst.cycle_cnt\[11\] VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__and4_1
X_0531_ net7 VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__inv_2
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1014_ ser_C.bit_idx\[0\] ser_C.bit_idx\[1\] net7 VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__and3_1
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0729_ deser_A.kept_shift_reg\[20\] deser_A.kept_shift_reg\[21\] net740 VGND VGND
+ VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_4_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload19 clknet_4_4_0_B_in_serial_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__bufinv_16
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_2_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_2_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0994_ deser_B.kept_shift_reg\[113\] deser_B.kept_shift_reg\[114\] net19 VGND VGND
+ VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1331_ clknet_4_3_0_B_in_serial_clk _0278_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_1400_ clknet_2_1__leaf_clk _0344_ net5 VGND VGND VPWR VPWR ser_C.kept_bit_idx\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1262_ clknet_4_11_0_B_in_serial_clk _0209_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput6 start VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1193_ clknet_4_0_0_A_in_serial_clk _0141_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_0977_ deser_B.kept_shift_reg\[96\] deser_B.kept_shift_reg\[97\] net47 VGND VGND
+ VPWR VPWR _0292_ sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_10_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0900_ deser_B.kept_shift_reg\[19\] deser_B.kept_shift_reg\[20\] net643 VGND VGND
+ VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_4
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0762_ deser_A.kept_shift_reg\[53\] deser_A.kept_shift_reg\[54\] net18 VGND VGND
+ VPWR VPWR _0105_ sky130_fd_sc_hd__mux2_4
X_0831_ deser_A.kept_shift_reg\[122\] deser_A.kept_shift_reg\[123\] net735 VGND VGND
+ VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_4
X_0693_ deser_A.kept_bit_idx\[2\] _0501_ _0514_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ clknet_4_0_0_B_in_serial_clk _0261_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_1245_ clknet_4_15_0_B_in_serial_clk _0193_ net15 VGND VGND VPWR VPWR deser_B.kept_bit_idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1176_ clknet_4_13_0_A_in_serial_clk _0124_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_3_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_46_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap13 deser_A.receiving VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ ser_C.bit_idx\[7\] _0383_ ser_C.bit_idx\[8\] VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0814_ deser_A.kept_shift_reg\[105\] deser_A.kept_shift_reg\[106\] net732 VGND VGND
+ VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_4
X_0676_ _0505_ _0501_ _0506_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__and3_1
X_0745_ deser_A.kept_shift_reg\[36\] deser_A.kept_shift_reg\[37\] net12 VGND VGND
+ VPWR VPWR _0088_ sky130_fd_sc_hd__mux2_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ clknet_4_2_0_A_in_serial_clk _0176_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_1159_ clknet_4_13_0_A_in_serial_clk _0107_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0530_ systolic_inst.cycle_cnt\[31\] VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__inv_2
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_11_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_64_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ ser_C.bit_idx\[0\] net7 VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__xor2_1
X_0659_ systolic_inst.cycle_cnt\[28\] systolic_inst.cycle_cnt\[29\] _0492_ VGND VGND
+ VPWR VPWR _0496_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0728_ deser_A.kept_shift_reg\[19\] deser_A.kept_shift_reg\[20\] net808 VGND VGND
+ VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_4_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer720 _0500_ VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0993_ deser_B.kept_shift_reg\[112\] deser_B.kept_shift_reg\[113\] net36 VGND VGND
+ VPWR VPWR _0308_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_14_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1261_ clknet_4_14_0_B_in_serial_clk _0208_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1330_ clknet_4_3_0_B_in_serial_clk _0277_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1192_ clknet_4_0_0_A_in_serial_clk _0140_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_0976_ deser_B.kept_shift_reg\[95\] deser_B.kept_shift_reg\[96\] net10 VGND VGND
+ VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0830_ deser_A.kept_shift_reg\[121\] deser_A.kept_shift_reg\[122\] net728 VGND VGND
+ VPWR VPWR _0173_ sky130_fd_sc_hd__mux2_4
X_0761_ deser_A.kept_shift_reg\[52\] deser_A.kept_shift_reg\[53\] net809 VGND VGND
+ VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_4
X_0692_ net13 deser_A.kept_bit_idx\[0\] deser_A.kept_bit_idx\[1\] deser_A.kept_bit_idx\[2\]
+ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__and4_1
X_1244_ clknet_4_15_0_B_in_serial_clk _0192_ net15 VGND VGND VPWR VPWR deser_B.kept_bit_idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1313_ clknet_4_0_0_B_in_serial_clk _0260_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1175_ clknet_4_13_0_A_in_serial_clk _0123_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_0959_ deser_B.kept_shift_reg\[78\] deser_B.kept_shift_reg\[79\] net47 VGND VGND
+ VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_34_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0813_ deser_A.kept_shift_reg\[104\] deser_A.kept_shift_reg\[105\] net12 VGND VGND
+ VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0675_ net21 net497 VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__nand2_2
XFILLER_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0744_ deser_A.kept_shift_reg\[35\] deser_A.kept_shift_reg\[36\] net12 VGND VGND
+ VPWR VPWR _0087_ sky130_fd_sc_hd__mux2_1
X_1158_ clknet_4_13_0_A_in_serial_clk _0106_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_1227_ clknet_4_2_0_A_in_serial_clk _0175_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1089_ clknet_4_10_0_A_in_serial_clk _0038_ net14 VGND VGND VPWR VPWR deser_A.bit_idx\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1012_ deser_A.kept_shift_reg\[0\] _0419_ _0500_ net2 _0376_ VGND VGND VPWR VPWR
+ _0325_ sky130_fd_sc_hd__a221o_1
XFILLER_21_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0727_ deser_A.kept_shift_reg\[18\] deser_A.kept_shift_reg\[19\] net44 VGND VGND
+ VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_2
X_0658_ systolic_inst.cycle_cnt\[29\] _0436_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nand2_1
X_0589_ systolic_inst.ce_local _0433_ _0441_ _0446_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__and4_2
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer721 _0348_ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_6
Xclone24 net41 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer798 net818 VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_31_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0992_ deser_B.kept_shift_reg\[111\] deser_B.kept_shift_reg\[112\] net36 VGND VGND
+ VPWR VPWR _0307_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_14_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1260_ clknet_4_14_0_B_in_serial_clk _0207_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1191_ clknet_4_0_0_A_in_serial_clk _0139_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0975_ deser_B.kept_shift_reg\[94\] deser_B.kept_shift_reg\[95\] net47 VGND VGND
+ VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1389_ clknet_2_0__leaf_clk _0334_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0760_ deser_A.kept_shift_reg\[51\] deser_A.kept_shift_reg\[52\] net40 VGND VGND
+ VPWR VPWR _0103_ sky130_fd_sc_hd__mux2_1
X_0691_ deser_A.kept_bit_idx\[0\] deser_A.kept_bit_idx\[1\] deser_A.kept_bit_idx\[2\]
+ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__and3_1
X_1243_ clknet_4_15_0_B_in_serial_clk _0191_ net15 VGND VGND VPWR VPWR deser_B.kept_bit_idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1312_ clknet_4_0_0_B_in_serial_clk _0259_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_1174_ clknet_4_13_0_A_in_serial_clk _0122_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0889_ deser_B.kept_shift_reg\[8\] deser_B.kept_shift_reg\[9\] net10 VGND VGND VPWR
+ VPWR _0204_ sky130_fd_sc_hd__mux2_1
X_0958_ deser_B.kept_shift_reg\[77\] deser_B.kept_shift_reg\[78\] net10 VGND VGND
+ VPWR VPWR _0273_ sky130_fd_sc_hd__mux2_1
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0812_ deser_A.kept_shift_reg\[103\] deser_A.kept_shift_reg\[104\] net730 VGND VGND
+ VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_4
X_0743_ deser_A.kept_shift_reg\[34\] deser_A.kept_shift_reg\[35\] net647 VGND VGND
+ VPWR VPWR _0086_ sky130_fd_sc_hd__mux2_4
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0674_ _0420_ net490 deser_A.bit_idx\[2\] net496 deser_A.bit_idx\[3\] VGND VGND VPWR
+ VPWR _0505_ sky130_fd_sc_hd__a41o_1
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1226_ clknet_4_0_0_A_in_serial_clk _0174_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_1157_ clknet_4_13_0_A_in_serial_clk _0105_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1088_ clknet_4_10_0_A_in_serial_clk _0037_ net14 VGND VGND VPWR VPWR deser_A.bit_idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1011_ net17 deser_A.kept_shift_reg\[1\] VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_62_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0726_ deser_A.kept_shift_reg\[17\] deser_A.kept_shift_reg\[18\] net18 VGND VGND
+ VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_4
X_0657_ _0492_ _0493_ _0494_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__o21a_1
X_0588_ _0433_ _0441_ _0446_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__and3_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1209_ clknet_4_5_0_A_in_serial_clk _0157_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0709_ _0527_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__inv_2
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ deser_B.kept_shift_reg\[110\] deser_B.kept_shift_reg\[111\] net845 VGND VGND
+ VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ clknet_4_0_0_A_in_serial_clk _0138_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0974_ deser_B.kept_shift_reg\[93\] deser_B.kept_shift_reg\[94\] net10 VGND VGND
+ VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_1
XFILLER_59_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1388_ clknet_2_0__leaf_clk _0333_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0690_ net736 _0513_ net810 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__nor3_2
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1311_ clknet_4_0_0_B_in_serial_clk _0258_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_1242_ clknet_4_15_0_B_in_serial_clk _0190_ net15 VGND VGND VPWR VPWR deser_B.kept_bit_idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclone831 net848 VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__clkbuf_16
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ clknet_4_15_0_A_in_serial_clk _0121_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0957_ deser_B.kept_shift_reg\[76\] deser_B.kept_shift_reg\[77\] net47 VGND VGND
+ VPWR VPWR _0272_ sky130_fd_sc_hd__mux2_1
X_0888_ deser_B.kept_shift_reg\[7\] deser_B.kept_shift_reg\[8\] net47 VGND VGND VPWR
+ VPWR _0203_ sky130_fd_sc_hd__mux2_1
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0811_ deser_A.kept_shift_reg\[102\] deser_A.kept_shift_reg\[103\] net12 VGND VGND
+ VPWR VPWR _0154_ sky130_fd_sc_hd__mux2_1
X_0673_ _0502_ _0503_ net493 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux2_4
X_0742_ deser_A.kept_shift_reg\[33\] deser_A.kept_shift_reg\[34\] net647 VGND VGND
+ VPWR VPWR _0085_ sky130_fd_sc_hd__mux2_4
X_1087_ clknet_2_3__leaf_clk _0036_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1156_ clknet_4_7_0_A_in_serial_clk _0104_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_1225_ clknet_4_2_0_A_in_serial_clk _0173_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1010_ _0425_ deser_B.kept_shift_reg\[0\] net500 net4 _0375_ VGND VGND VPWR VPWR
+ _0324_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_6_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0656_ systolic_inst.cycle_cnt\[28\] _0492_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__nand2_1
X_0725_ deser_A.kept_shift_reg\[16\] deser_A.kept_shift_reg\[17\] net808 VGND VGND
+ VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_4
X_0587_ systolic_inst.cycle_cnt\[5\] systolic_inst.cycle_cnt\[6\] systolic_inst.cycle_cnt\[7\]
+ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__and3_1
X_1208_ clknet_4_5_0_A_in_serial_clk _0156_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1139_ clknet_4_2_0_A_in_serial_clk _0087_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer723 net13 VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_3_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0639_ _0399_ _0481_ _0480_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux2_1
X_0708_ deser_A.kept_bit_idx\[7\] _0526_ _0524_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__mux2_4
XFILLER_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0990_ deser_B.kept_shift_reg\[109\] deser_B.kept_shift_reg\[110\] net27 VGND VGND
+ VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0973_ deser_B.kept_shift_reg\[92\] deser_B.kept_shift_reg\[93\] net27 VGND VGND
+ VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
X_1387_ clknet_2_1__leaf_clk _0332_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1241_ clknet_4_15_0_B_in_serial_clk _0189_ net15 VGND VGND VPWR VPWR deser_B.kept_bit_idx\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1310_ clknet_4_0_0_B_in_serial_clk _0257_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ clknet_4_15_0_A_in_serial_clk _0120_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[68\]
+ sky130_fd_sc_hd__dfrtp_1
X_0956_ deser_B.kept_shift_reg\[75\] deser_B.kept_shift_reg\[76\] net10 VGND VGND
+ VPWR VPWR _0271_ sky130_fd_sc_hd__mux2_1
XFILLER_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0887_ deser_B.kept_shift_reg\[6\] deser_B.kept_shift_reg\[7\] net10 VGND VGND VPWR
+ VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0810_ deser_A.kept_shift_reg\[101\] deser_A.kept_shift_reg\[102\] net728 VGND VGND
+ VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_4
X_0672_ _0503_ _0504_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__and2_1
X_0741_ deser_A.kept_shift_reg\[32\] deser_A.kept_shift_reg\[33\] net728 VGND VGND
+ VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_4
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1224_ clknet_4_2_0_A_in_serial_clk _0172_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_1086_ clknet_2_3__leaf_clk _0035_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_1155_ clknet_4_7_0_A_in_serial_clk _0103_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_0939_ deser_B.kept_shift_reg\[58\] deser_B.kept_shift_reg\[59\] net47 VGND VGND
+ VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
XFILLER_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0655_ systolic_inst.cycle_cnt\[28\] _0436_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__and2_1
X_0586_ systolic_inst.cycle_cnt\[5\] systolic_inst.cycle_cnt\[6\] _0444_ systolic_inst.cycle_cnt\[7\]
+ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a31o_1
X_0724_ deser_A.kept_shift_reg\[15\] deser_A.kept_shift_reg\[16\] net740 VGND VGND
+ VPWR VPWR _0067_ sky130_fd_sc_hd__mux2_2
X_1207_ clknet_4_5_0_A_in_serial_clk _0155_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1069_ clknet_2_2__leaf_clk _0018_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1138_ clknet_4_2_0_A_in_serial_clk _0086_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer713 net22 VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__clkbuf_2
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0707_ deser_A.kept_bit_idx\[7\] _0501_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__nand2_1
X_0569_ systolic_inst.ce_local systolic_inst.cycle_cnt\[0\] systolic_inst.cycle_cnt\[1\]
+ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__and3_1
X_0638_ _0399_ _0435_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__nor2_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0972_ deser_B.kept_shift_reg\[91\] deser_B.kept_shift_reg\[92\] net27 VGND VGND
+ VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_5_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1386_ clknet_2_1__leaf_clk _0331_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1240_ clknet_4_15_0_B_in_serial_clk _0188_ net15 VGND VGND VPWR VPWR deser_B.kept_bit_idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1171_ clknet_4_14_0_A_in_serial_clk _0119_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_0886_ deser_B.kept_shift_reg\[5\] deser_B.kept_shift_reg\[6\] net47 VGND VGND VPWR
+ VPWR _0201_ sky130_fd_sc_hd__mux2_1
X_0955_ deser_B.kept_shift_reg\[74\] deser_B.kept_shift_reg\[75\] net47 VGND VGND
+ VPWR VPWR _0270_ sky130_fd_sc_hd__mux2_1
XFILLER_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1369_ clknet_4_5_0_B_in_serial_clk _0316_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_13_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0740_ deser_A.kept_shift_reg\[31\] deser_A.kept_shift_reg\[32\] net17 VGND VGND
+ VPWR VPWR _0083_ sky130_fd_sc_hd__mux2_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0671_ _0420_ net492 net495 VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__a21o_1
Xclone630 net641 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__clkbuf_16
X_1154_ clknet_4_7_0_A_in_serial_clk _0102_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_1223_ clknet_4_2_0_A_in_serial_clk _0171_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1085_ clknet_2_3__leaf_clk _0034_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_0869_ deser_B.kept_bit_idx\[3\] deser_B.kept_bit_idx\[4\] net31 _0366_ VGND VGND
+ VPWR VPWR _0367_ sky130_fd_sc_hd__a31o_1
X_0938_ deser_B.kept_shift_reg\[57\] deser_B.kept_shift_reg\[58\] net47 VGND VGND
+ VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
XFILLER_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_6_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_6_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0723_ deser_A.kept_shift_reg\[14\] deser_A.kept_shift_reg\[15\] net769 VGND VGND
+ VPWR VPWR _0066_ sky130_fd_sc_hd__mux2_4
X_0585_ _0442_ _0443_ systolic_inst.cycle_cnt\[6\] VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__mux2_1
X_0654_ _0489_ _0490_ _0492_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__o21ba_1
XFILLER_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1206_ clknet_4_5_0_A_in_serial_clk _0154_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_1137_ clknet_4_2_0_A_in_serial_clk _0085_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_25_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1068_ clknet_2_0__leaf_clk _0017_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_14_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0706_ _0524_ _0525_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__and2_4
X_0568_ systolic_inst.cycle_cnt\[0\] systolic_inst.cycle_cnt\[1\] VGND VGND VPWR VPWR
+ _0433_ sky130_fd_sc_hd__and2_1
X_0637_ _0477_ _0478_ _0480_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__a21boi_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0971_ deser_B.kept_shift_reg\[90\] deser_B.kept_shift_reg\[91\] net19 VGND VGND
+ VPWR VPWR _0286_ sky130_fd_sc_hd__mux2_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1385_ clknet_2_0__leaf_clk _0330_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ clknet_4_15_0_A_in_serial_clk _0118_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0885_ deser_B.kept_shift_reg\[4\] deser_B.kept_shift_reg\[5\] net47 VGND VGND VPWR
+ VPWR _0200_ sky130_fd_sc_hd__mux2_1
X_0954_ deser_B.kept_shift_reg\[73\] deser_B.kept_shift_reg\[74\] net10 VGND VGND
+ VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1368_ clknet_4_5_0_B_in_serial_clk _0315_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1299_ clknet_4_2_0_B_in_serial_clk _0246_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0670_ _0500_ _0502_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__nor2_1
XFILLER_42_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1084_ clknet_2_3__leaf_clk _0033_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1153_ clknet_4_13_0_A_in_serial_clk _0101_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_1222_ clknet_4_0_0_A_in_serial_clk _0170_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[118\]
+ sky130_fd_sc_hd__dfrtp_1
Xclone631 net733 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__clkbuf_16
X_0868_ _0348_ deser_B.kept_bit_idx\[4\] net31 deser_B.kept_bit_idx\[3\] VGND VGND
+ VPWR VPWR _0366_ sky130_fd_sc_hd__a22oi_2
X_0937_ deser_B.kept_shift_reg\[56\] deser_B.kept_shift_reg\[57\] net10 VGND VGND
+ VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
X_0799_ deser_A.kept_shift_reg\[90\] deser_A.kept_shift_reg\[91\] net647 VGND VGND
+ VPWR VPWR _0142_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_58_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0653_ _0448_ _0464_ _0482_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__and4_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0722_ deser_A.kept_shift_reg\[13\] deser_A.kept_shift_reg\[14\] net44 VGND VGND
+ VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_2
X_0584_ systolic_inst.cycle_cnt\[5\] _0444_ _0443_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__o21a_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1067_ clknet_2_2__leaf_clk _0016_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1136_ clknet_4_2_0_A_in_serial_clk _0084_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_1205_ clknet_4_5_0_A_in_serial_clk _0153_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[101\]
+ sky130_fd_sc_hd__dfrtp_1
Xclone29 net37 net3 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__nand2b_2
Xrebuffer715 net22 VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__buf_8
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0636_ _0474_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nand2_1
X_0705_ deser_A.kept_bit_idx\[6\] _0501_ _0521_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__a21o_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0567_ systolic_inst.ce_local systolic_inst.cycle_cnt\[0\] systolic_inst.cycle_cnt\[1\]
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a21o_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ clknet_4_11_0_A_in_serial_clk _0067_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0619_ systolic_inst.cycle_cnt\[16\] systolic_inst.cycle_cnt\[17\] _0465_ VGND VGND
+ VPWR VPWR _0468_ sky130_fd_sc_hd__and3_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0970_ deser_B.kept_shift_reg\[89\] deser_B.kept_shift_reg\[90\] net47 VGND VGND
+ VPWR VPWR _0285_ sky130_fd_sc_hd__mux2_1
X_1384_ clknet_2_0__leaf_clk _0329_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0884_ deser_B.kept_shift_reg\[3\] deser_B.kept_shift_reg\[4\] net27 VGND VGND VPWR
+ VPWR _0199_ sky130_fd_sc_hd__mux2_1
X_0953_ deser_B.kept_shift_reg\[72\] deser_B.kept_shift_reg\[73\] net10 VGND VGND
+ VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1367_ clknet_4_5_0_B_in_serial_clk _0314_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1298_ clknet_4_2_0_B_in_serial_clk _0245_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1221_ clknet_4_1_0_A_in_serial_clk _0169_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1083_ clknet_2_3__leaf_clk _0032_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1152_ clknet_4_7_0_A_in_serial_clk _0100_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0936_ deser_B.kept_shift_reg\[55\] deser_B.kept_shift_reg\[56\] net47 VGND VGND
+ VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
X_0867_ deser_B.kept_bit_idx\[3\] net33 _0365_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a21oi_1
X_0798_ deser_A.kept_shift_reg\[89\] deser_A.kept_shift_reg\[90\] net735 VGND VGND
+ VPWR VPWR _0141_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_58_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0583_ _0428_ _0433_ _0441_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__and3_1
X_0652_ systolic_inst.cycle_cnt\[26\] systolic_inst.cycle_cnt\[27\] _0486_ VGND VGND
+ VPWR VPWR _0491_ sky130_fd_sc_hd__and3_1
X_0721_ deser_A.kept_shift_reg\[12\] deser_A.kept_shift_reg\[13\] net18 VGND VGND
+ VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1204_ clknet_4_5_0_A_in_serial_clk _0152_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1066_ clknet_2_2__leaf_clk _0015_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1135_ clknet_4_3_0_A_in_serial_clk _0083_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_0919_ deser_B.kept_shift_reg\[38\] deser_B.kept_shift_reg\[39\] net11 VGND VGND
+ VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0566_ systolic_inst.ce_local _0427_ systolic_inst.cycle_cnt\[0\] VGND VGND VPWR
+ VPWR _0005_ sky130_fd_sc_hd__mux2_1
X_0635_ systolic_inst.cycle_cnt\[20\] systolic_inst.cycle_cnt\[21\] systolic_inst.cycle_cnt\[22\]
+ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and3_1
X_0704_ deser_A.kept_bit_idx\[6\] _0521_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nand2_2
XFILLER_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1118_ clknet_4_11_0_A_in_serial_clk _0066_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1049_ ser_C.kept_bit_idx\[6\] ser_C.kept_bit_idx\[7\] _0393_ VGND VGND VPWR VPWR
+ _0395_ sky130_fd_sc_hd__and3_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0618_ _0465_ _0466_ systolic_inst.cycle_cnt\[16\] VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__mux2_1
X_0549_ net1 net22 VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__nor2_1
XFILLER_65_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_46_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_55_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1383_ clknet_2_0__leaf_clk _0328_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0952_ deser_B.kept_shift_reg\[71\] deser_B.kept_shift_reg\[72\] net10 VGND VGND
+ VPWR VPWR _0267_ sky130_fd_sc_hd__mux2_1
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0883_ deser_B.kept_shift_reg\[2\] deser_B.kept_shift_reg\[3\] net27 VGND VGND VPWR
+ VPWR _0198_ sky130_fd_sc_hd__mux2_1
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1366_ clknet_4_7_0_B_in_serial_clk _0313_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1297_ clknet_4_8_0_B_in_serial_clk _0244_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_0_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1151_ clknet_4_7_0_A_in_serial_clk _0099_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_1220_ clknet_4_1_0_A_in_serial_clk _0168_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1082_ clknet_2_3__leaf_clk _0031_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_0866_ deser_B.kept_bit_idx\[3\] _0348_ net32 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__a21oi_1
X_0935_ deser_B.kept_shift_reg\[54\] deser_B.kept_shift_reg\[55\] net646 VGND VGND
+ VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_4
X_0797_ deser_A.kept_shift_reg\[88\] deser_A.kept_shift_reg\[89\] net732 VGND VGND
+ VPWR VPWR _0140_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_58_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1349_ clknet_4_4_0_B_in_serial_clk _0296_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0720_ deser_A.kept_shift_reg\[11\] deser_A.kept_shift_reg\[12\] net769 VGND VGND
+ VPWR VPWR _0063_ sky130_fd_sc_hd__mux2_4
X_0582_ _0435_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__nor2_1
X_0651_ systolic_inst.cycle_cnt\[27\] _0436_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__and2_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1134_ clknet_4_3_0_A_in_serial_clk _0082_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_1203_ clknet_4_4_0_A_in_serial_clk _0151_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1065_ clknet_2_2__leaf_clk _0014_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_0849_ deser_B.bit_idx\[4\] _0354_ _0353_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_4
X_0918_ deser_B.kept_shift_reg\[37\] deser_B.kept_shift_reg\[38\] net11 VGND VGND
+ VPWR VPWR _0233_ sky130_fd_sc_hd__mux2_1
Xrebuffer717 net22 VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__buf_8
XFILLER_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone2 net24 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_16
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0703_ _0501_ _0522_ _0523_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_29_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0634_ systolic_inst.cycle_cnt\[22\] _0436_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_13_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0565_ _0431_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__inv_2
XFILLER_65_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ clknet_4_14_0_A_in_serial_clk _0065_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_1_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1048_ ser_C.kept_bit_idx\[6\] _0393_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__xor2_1
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xsplit11 net820 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_12
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0617_ systolic_inst.cycle_cnt\[15\] _0466_ _0467_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a21o_1
X_0548_ deser_A.bit_idx\[7\] net509 VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_36_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1382_ clknet_2_0__leaf_clk _0327_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0882_ deser_B.kept_shift_reg\[1\] deser_B.kept_shift_reg\[2\] net19 VGND VGND VPWR
+ VPWR _0197_ sky130_fd_sc_hd__mux2_2
X_0951_ deser_B.kept_shift_reg\[70\] deser_B.kept_shift_reg\[71\] net10 VGND VGND
+ VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1365_ clknet_4_7_0_B_in_serial_clk _0312_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_1296_ clknet_4_8_0_B_in_serial_clk _0243_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1150_ clknet_4_7_0_A_in_serial_clk _0098_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1081_ clknet_2_3__leaf_clk _0030_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_0865_ _0363_ _0364_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__nor2_1
X_0934_ deser_B.kept_shift_reg\[53\] deser_B.kept_shift_reg\[54\] net646 VGND VGND
+ VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_4
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0796_ deser_A.kept_shift_reg\[87\] deser_A.kept_shift_reg\[88\] net735 VGND VGND
+ VPWR VPWR _0139_ sky130_fd_sc_hd__mux2_4
X_1348_ clknet_4_4_0_B_in_serial_clk _0295_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_1279_ clknet_4_2_0_B_in_serial_clk _0226_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0581_ systolic_inst.cycle_cnt\[5\] _0434_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__and3_1
X_0650_ _0487_ _0488_ _0489_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1064_ clknet_2_3__leaf_clk _0013_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1133_ clknet_4_3_0_A_in_serial_clk _0081_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1202_ clknet_4_4_0_A_in_serial_clk _0150_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0848_ net737 deser_B.bit_idx\[4\] VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__nand2_2
X_0917_ deser_B.kept_shift_reg\[36\] deser_B.kept_shift_reg\[37\] net11 VGND VGND
+ VPWR VPWR _0232_ sky130_fd_sc_hd__mux2_1
X_0779_ deser_A.kept_shift_reg\[70\] deser_A.kept_shift_reg\[71\] net769 VGND VGND
+ VPWR VPWR _0122_ sky130_fd_sc_hd__mux2_4
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0633_ _0436_ _0476_ _0477_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__and3_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0702_ deser_A.kept_bit_idx\[3\] deser_A.kept_bit_idx\[4\] _0420_ _0515_ deser_A.kept_bit_idx\[5\]
+ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__a41o_1
X_0564_ ser_C.bit_idx\[5\] ser_C.bit_idx\[4\] _0429_ _0430_ _0402_ VGND VGND VPWR
+ VPWR _0431_ sky130_fd_sc_hd__a41o_1
XFILLER_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1116_ clknet_4_14_0_A_in_serial_clk _0064_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1047_ _0393_ _0394_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__and2b_1
XFILLER_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0616_ _0465_ _0463_ _0456_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__and3b_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0547_ _0416_ deser_A.bit_idx\[5\] deser_A.bit_idx\[6\] net20 VGND VGND VPWR VPWR
+ _0417_ sky130_fd_sc_hd__nand4_4
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1381_ clknet_2_0__leaf_clk _0326_ net5 VGND VGND VPWR VPWR ser_C.bit_idx\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0950_ deser_B.kept_shift_reg\[69\] deser_B.kept_shift_reg\[70\] net10 VGND VGND
+ VPWR VPWR _0265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0881_ _0403_ _0418_ _0501_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1364_ clknet_4_6_0_B_in_serial_clk _0311_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_1295_ clknet_4_8_0_B_in_serial_clk _0242_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_8_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_8_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1080_ clknet_2_3__leaf_clk _0029_ net5 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xclone624 net641 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkbuf_16
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0864_ deser_B.kept_bit_idx\[2\] net45 _0361_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__a21oi_1
X_0933_ deser_B.kept_shift_reg\[52\] deser_B.kept_shift_reg\[53\] net642 VGND VGND
+ VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_4
X_0795_ deser_A.kept_shift_reg\[86\] deser_A.kept_shift_reg\[87\] net735 VGND VGND
+ VPWR VPWR _0138_ sky130_fd_sc_hd__mux2_4
X_1347_ clknet_4_4_0_B_in_serial_clk _0294_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ clknet_4_2_0_B_in_serial_clk _0225_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0580_ systolic_inst.cycle_cnt\[2\] systolic_inst.cycle_cnt\[3\] systolic_inst.cycle_cnt\[4\]
+ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__and3_1
X_1201_ clknet_4_4_0_A_in_serial_clk _0149_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1063_ clknet_2_3__leaf_clk _0012_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1132_ clknet_4_3_0_A_in_serial_clk _0080_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_0916_ deser_B.kept_shift_reg\[35\] deser_B.kept_shift_reg\[36\] net11 VGND VGND
+ VPWR VPWR _0231_ sky130_fd_sc_hd__mux2_1
X_0847_ _0352_ net45 _0353_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__and3_1
X_0778_ deser_A.kept_shift_reg\[69\] deser_A.kept_shift_reg\[70\] net40 VGND VGND
+ VPWR VPWR _0121_ sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_9_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0632_ systolic_inst.cycle_cnt\[20\] systolic_inst.cycle_cnt\[21\] _0474_ VGND VGND
+ VPWR VPWR _0477_ sky130_fd_sc_hd__nand3_1
X_0701_ net39 VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__inv_2
X_0563_ ser_C.bit_idx\[0\] ser_C.bit_idx\[1\] ser_C.bit_idx\[2\] ser_C.bit_idx\[3\]
+ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__and4_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1115_ clknet_4_11_0_A_in_serial_clk _0063_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1046_ ser_C.kept_bit_idx\[3\] ser_C.kept_bit_idx\[4\] _0389_ ser_C.kept_bit_idx\[5\]
+ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__a31o_1
XFILLER_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_35_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0615_ _0435_ _0465_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__nor2_1
X_0546_ _0415_ deser_A.bit_idx\[4\] VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__and2_4
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1029_ ser_C.bit_idx\[7\] ser_C.bit_idx\[8\] _0383_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__and3_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1380_ clknet_2_2__leaf_clk _0003_ net5 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ systolic_inst.cycle_cnt\[30\] VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__inv_2
Xrebuffer20 net34 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_6
XFILLER_26_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0880_ _0374_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1363_ clknet_4_6_0_B_in_serial_clk _0310_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1294_ clknet_4_8_0_B_in_serial_clk _0241_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0932_ deser_B.kept_shift_reg\[51\] deser_B.kept_shift_reg\[52\] net646 VGND VGND
+ VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_4
X_0863_ deser_B.kept_bit_idx\[1\] deser_B.kept_bit_idx\[0\] deser_B.receiving deser_B.kept_bit_idx\[2\]
+ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__and4_1
XFILLER_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0794_ deser_A.kept_shift_reg\[85\] deser_A.kept_shift_reg\[86\] net647 VGND VGND
+ VPWR VPWR _0137_ sky130_fd_sc_hd__mux2_4
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1346_ clknet_4_4_0_B_in_serial_clk _0293_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1277_ clknet_4_8_0_B_in_serial_clk _0224_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1200_ clknet_4_4_0_A_in_serial_clk _0148_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_1062_ clknet_2_3__leaf_clk _0011_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1131_ clknet_4_6_0_A_in_serial_clk _0079_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_0915_ deser_B.kept_shift_reg\[34\] deser_B.kept_shift_reg\[35\] net11 VGND VGND
+ VPWR VPWR _0230_ sky130_fd_sc_hd__mux2_1
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0846_ net35 net506 VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__nand2_2
X_0777_ deser_A.kept_shift_reg\[68\] deser_A.kept_shift_reg\[69\] net808 VGND VGND
+ VPWR VPWR _0120_ sky130_fd_sc_hd__mux2_4
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1329_ clknet_4_3_0_B_in_serial_clk _0276_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0700_ deser_A.kept_bit_idx\[3\] deser_A.kept_bit_idx\[4\] _0516_ deser_A.kept_bit_idx\[5\]
+ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and4_1
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0631_ systolic_inst.cycle_cnt\[20\] _0470_ _0473_ systolic_inst.cycle_cnt\[21\]
+ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__a31o_1
X_0562_ ser_C.bit_idx\[9\] ser_C.bit_idx\[8\] ser_C.bit_idx\[7\] ser_C.bit_idx\[6\]
+ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__and4b_1
X_1114_ clknet_4_11_0_A_in_serial_clk _0062_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ ser_C.kept_bit_idx\[3\] ser_C.kept_bit_idx\[4\] ser_C.kept_bit_idx\[5\] _0389_
+ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__and4_1
X_0829_ deser_A.kept_shift_reg\[120\] deser_A.kept_shift_reg\[121\] net12 VGND VGND
+ VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0614_ _0448_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__and2_1
X_0545_ deser_A.bit_idx\[2\] deser_A.bit_idx\[0\] deser_A.bit_idx\[3\] deser_A.bit_idx\[1\]
+ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1028_ ser_C.bit_idx\[7\] _0383_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__xor2_1
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xsplit1 net814 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_33_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0528_ systolic_inst.cycle_cnt\[23\] VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__inv_2
Xrebuffer21 net34 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_6
Xrebuffer10 net22 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone829 net846 VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__clkbuf_16
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1362_ clknet_4_5_0_B_in_serial_clk _0309_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_1293_ clknet_4_8_0_B_in_serial_clk _0240_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_52_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone626 net641 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__buf_8
X_0862_ deser_B.kept_bit_idx\[0\] deser_B.kept_bit_idx\[1\] deser_B.kept_bit_idx\[2\]
+ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ deser_B.kept_shift_reg\[50\] deser_B.kept_shift_reg\[51\] net643 VGND VGND
+ VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_4
XFILLER_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0793_ deser_A.kept_shift_reg\[84\] deser_A.kept_shift_reg\[85\] net732 VGND VGND
+ VPWR VPWR _0136_ sky130_fd_sc_hd__mux2_4
X_1345_ clknet_4_4_0_B_in_serial_clk _0292_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_1276_ clknet_4_8_0_B_in_serial_clk _0223_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1130_ clknet_4_6_0_A_in_serial_clk _0078_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1061_ clknet_2_2__leaf_clk _0010_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0845_ _0426_ deser_B.bit_idx\[0\] net504 net505 deser_B.bit_idx\[3\] VGND VGND VPWR
+ VPWR _0352_ sky130_fd_sc_hd__a41o_1
X_0914_ deser_B.kept_shift_reg\[33\] deser_B.kept_shift_reg\[34\] net11 VGND VGND
+ VPWR VPWR _0229_ sky130_fd_sc_hd__mux2_1
X_0776_ deser_A.kept_shift_reg\[67\] deser_A.kept_shift_reg\[68\] net18 VGND VGND
+ VPWR VPWR _0119_ sky130_fd_sc_hd__mux2_4
X_1259_ clknet_4_11_0_B_in_serial_clk _0206_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1328_ clknet_4_3_0_B_in_serial_clk _0275_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0561_ _0003_ _0427_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__nor2_1
X_0630_ _0474_ _0475_ systolic_inst.cycle_cnt\[20\] VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__mux2_1
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1113_ clknet_4_9_0_A_in_serial_clk _0061_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1044_ ser_C.kept_bit_idx\[4\] _0391_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__xnor2_1
X_0759_ deser_A.kept_shift_reg\[50\] deser_A.kept_shift_reg\[51\] net40 VGND VGND
+ VPWR VPWR _0102_ sky130_fd_sc_hd__mux2_1
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0828_ deser_A.kept_shift_reg\[119\] deser_A.kept_shift_reg\[120\] net732 VGND VGND
+ VPWR VPWR _0171_ sky130_fd_sc_hd__mux2_4
XFILLER_28_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0613_ systolic_inst.cycle_cnt\[15\] _0455_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__and3_1
XFILLER_7_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0544_ systolic_inst.cycle_cnt\[11\] _0413_ _0414_ systolic_inst.ce_local VGND VGND
+ VPWR VPWR _0003_ sky130_fd_sc_hd__o31a_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1027_ _0383_ _0384_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer22 net37 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_6
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1361_ clknet_4_4_0_B_in_serial_clk _0308_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_1292_ clknet_4_10_0_B_in_serial_clk _0239_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone627 net641 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_9_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0861_ net499 _0360_ _0361_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__nor3_1
X_0930_ deser_B.kept_shift_reg\[49\] deser_B.kept_shift_reg\[50\] net646 VGND VGND
+ VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
X_0792_ deser_A.kept_shift_reg\[83\] deser_A.kept_shift_reg\[84\] net12 VGND VGND
+ VPWR VPWR _0135_ sky130_fd_sc_hd__mux2_1
XFILLER_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1344_ clknet_4_6_0_B_in_serial_clk _0291_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_1275_ clknet_4_9_0_B_in_serial_clk _0222_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1060_ clknet_2_2__leaf_clk _0009_ net15 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_3_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_3_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0844_ _0349_ _0350_ net503 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux2_4
X_0913_ deser_B.kept_shift_reg\[32\] deser_B.kept_shift_reg\[33\] net11 VGND VGND
+ VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_1
X_0775_ deser_A.kept_shift_reg\[66\] deser_A.kept_shift_reg\[67\] net40 VGND VGND
+ VPWR VPWR _0118_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1258_ clknet_4_11_0_B_in_serial_clk _0205_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1327_ clknet_4_3_0_B_in_serial_clk _0274_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_1189_ clknet_4_0_0_A_in_serial_clk _0137_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0560_ net6 systolic_inst.ce_local VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__or2_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1112_ clknet_4_9_0_A_in_serial_clk _0060_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1043_ _0391_ _0392_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__and2_1
X_0758_ deser_A.kept_shift_reg\[49\] deser_A.kept_shift_reg\[50\] net809 VGND VGND
+ VPWR VPWR _0101_ sky130_fd_sc_hd__mux2_4
X_0827_ deser_A.kept_shift_reg\[118\] deser_A.kept_shift_reg\[119\] net734 VGND VGND
+ VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_24_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0689_ net809 deser_A.kept_bit_idx\[0\] deser_A.kept_bit_idx\[1\] VGND VGND VPWR
+ VPWR _0514_ sky130_fd_sc_hd__and3_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_4_11_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0612_ systolic_inst.cycle_cnt\[14\] _0461_ _0462_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0543_ _0408_ _0409_ _0410_ _0411_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or4_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1026_ ser_C.bit_idx\[5\] _0381_ ser_C.bit_idx\[6\] VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_4_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xsplit3 deser_B.receiving VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_12
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer23 _0521_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
Xrebuffer12 _0516_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_6
X_1009_ net19 deser_B.kept_shift_reg\[1\] VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__and2_1
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ clknet_4_5_0_B_in_serial_clk _0307_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1291_ clknet_4_10_0_B_in_serial_clk _0238_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_12_0_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_4_12_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_46_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0860_ net845 deser_B.kept_bit_idx\[0\] deser_B.kept_bit_idx\[1\] VGND VGND VPWR
+ VPWR _0361_ sky130_fd_sc_hd__and3_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0791_ deser_A.kept_shift_reg\[82\] deser_A.kept_shift_reg\[83\] net734 VGND VGND
+ VPWR VPWR _0134_ sky130_fd_sc_hd__mux2_4
X_1343_ clknet_4_6_0_B_in_serial_clk _0290_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1274_ clknet_4_8_0_B_in_serial_clk _0221_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_0989_ deser_B.kept_shift_reg\[108\] deser_B.kept_shift_reg\[109\] net847 VGND VGND
+ VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0912_ deser_B.kept_shift_reg\[31\] deser_B.kept_shift_reg\[32\] net11 VGND VGND
+ VPWR VPWR _0227_ sky130_fd_sc_hd__mux2_1
X_0843_ _0350_ _0351_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__and2_4
X_0774_ deser_A.kept_shift_reg\[65\] deser_A.kept_shift_reg\[66\] net44 VGND VGND
+ VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_2
XFILLER_56_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_B_in_serial_clk B_in_serial_clk VGND VGND VPWR VPWR clknet_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
X_1326_ clknet_4_1_0_B_in_serial_clk _0273_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_1257_ clknet_4_11_0_B_in_serial_clk _0204_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1188_ clknet_4_0_0_A_in_serial_clk _0136_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1111_ clknet_4_9_0_A_in_serial_clk _0059_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1042_ ser_C.kept_bit_idx\[3\] _0389_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or2_1
XFILLER_61_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0757_ deser_A.kept_shift_reg\[48\] deser_A.kept_shift_reg\[49\] net809 VGND VGND
+ VPWR VPWR _0100_ sky130_fd_sc_hd__mux2_4
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0688_ deser_A.kept_bit_idx\[0\] _0420_ deser_A.kept_bit_idx\[1\] VGND VGND VPWR
+ VPWR _0513_ sky130_fd_sc_hd__a21oi_1
X_0826_ deser_A.kept_shift_reg\[117\] deser_A.kept_shift_reg\[118\] net12 VGND VGND
+ VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1309_ clknet_4_2_0_B_in_serial_clk _0256_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0542_ _0405_ _0406_ _0407_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__or4_1
X_0611_ systolic_inst.cycle_cnt\[12\] systolic_inst.cycle_cnt\[13\] systolic_inst.cycle_cnt\[14\]
+ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__and3_1
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1025_ ser_C.bit_idx\[5\] ser_C.bit_idx\[6\] _0381_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__and3_1
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0809_ deser_A.kept_shift_reg\[100\] deser_A.kept_shift_reg\[101\] net12 VGND VGND
+ VPWR VPWR _0152_ sky130_fd_sc_hd__mux2_1
XFILLER_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer13 net28 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s4s_1
X_1008_ deser_B.kept_shift_reg\[127\] net4 net845 VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ clknet_4_11_0_B_in_serial_clk _0237_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer4 net814 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
X_0790_ deser_A.kept_shift_reg\[81\] deser_A.kept_shift_reg\[82\] net732 VGND VGND
+ VPWR VPWR _0133_ sky130_fd_sc_hd__mux2_4
X_1342_ clknet_4_6_0_B_in_serial_clk _0289_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[93\]
+ sky130_fd_sc_hd__dfrtp_1
X_1273_ clknet_4_8_0_B_in_serial_clk _0220_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0988_ deser_B.kept_shift_reg\[107\] deser_B.kept_shift_reg\[108\] net845 VGND VGND
+ VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
XFILLER_47_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0842_ _0426_ net502 deser_B.bit_idx\[1\] VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a21o_1
X_0911_ deser_B.kept_shift_reg\[30\] deser_B.kept_shift_reg\[31\] net640 VGND VGND
+ VPWR VPWR _0226_ sky130_fd_sc_hd__mux2_4
XFILLER_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0773_ deser_A.kept_shift_reg\[64\] deser_A.kept_shift_reg\[65\] net44 VGND VGND
+ VPWR VPWR _0116_ sky130_fd_sc_hd__mux2_2
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1325_ clknet_4_4_0_B_in_serial_clk _0272_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_1256_ clknet_4_9_0_B_in_serial_clk _0203_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1187_ clknet_4_1_0_A_in_serial_clk _0135_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ clknet_4_9_0_A_in_serial_clk _0058_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1041_ ser_C.kept_bit_idx\[3\] _0389_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__nand2_1
X_0825_ deser_A.kept_shift_reg\[116\] deser_A.kept_shift_reg\[117\] net647 VGND VGND
+ VPWR VPWR _0168_ sky130_fd_sc_hd__mux2_4
X_0756_ deser_A.kept_shift_reg\[47\] deser_A.kept_shift_reg\[48\] net40 VGND VGND
+ VPWR VPWR _0099_ sky130_fd_sc_hd__mux2_1
X_0687_ net17 _0419_ deser_A.kept_bit_idx\[0\] VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux2_1
XFILLER_56_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1239_ clknet_4_14_0_B_in_serial_clk _0187_ net15 VGND VGND VPWR VPWR deser_B.bit_idx\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1308_ clknet_4_0_0_B_in_serial_clk _0255_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0610_ systolic_inst.cycle_cnt\[14\] _0436_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a21oi_1
X_0541_ systolic_inst.cycle_cnt\[16\] systolic_inst.cycle_cnt\[17\] systolic_inst.cycle_cnt\[18\]
+ systolic_inst.cycle_cnt\[19\] VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or4_1
X_1024_ ser_C.bit_idx\[5\] _0381_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__xor2_1
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0808_ deser_A.kept_shift_reg\[99\] deser_A.kept_shift_reg\[100\] net732 VGND VGND
+ VPWR VPWR _0151_ sky130_fd_sc_hd__mux2_4
XFILLER_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0739_ deser_A.kept_shift_reg\[30\] deser_A.kept_shift_reg\[31\] net17 VGND VGND
+ VPWR VPWR _0082_ sky130_fd_sc_hd__mux2_1
XFILLER_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer830 deser_B.receiving VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_35_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_2 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ deser_B.kept_shift_reg\[126\] deser_B.kept_shift_reg\[127\] net27 VGND VGND
+ VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer25 deser_A.receiving VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xrebuffer14 net28 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer490 _0421_ VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer5 net20 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
X_1341_ clknet_4_6_0_B_in_serial_clk _0288_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[92\]
+ sky130_fd_sc_hd__dfrtp_1
X_1272_ clknet_4_10_0_B_in_serial_clk _0219_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0987_ deser_B.kept_shift_reg\[106\] deser_B.kept_shift_reg\[107\] net845 VGND VGND
+ VPWR VPWR _0302_ sky130_fd_sc_hd__mux2_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0841_ _0349_ _0347_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__nor2_2
X_0910_ deser_B.kept_shift_reg\[29\] deser_B.kept_shift_reg\[30\] net646 VGND VGND
+ VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_4
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0772_ deser_A.kept_shift_reg\[63\] deser_A.kept_shift_reg\[64\] net769 VGND VGND
+ VPWR VPWR _0115_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ clknet_4_12_0_B_in_serial_clk _0202_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1324_ clknet_4_1_0_B_in_serial_clk _0271_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ clknet_4_1_0_A_in_serial_clk _0134_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1040_ _0389_ _0390_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__and2b_1
XFILLER_14_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0755_ deser_A.kept_shift_reg\[46\] deser_A.kept_shift_reg\[47\] net730 VGND VGND
+ VPWR VPWR _0098_ sky130_fd_sc_hd__mux2_4
X_0824_ deser_A.kept_shift_reg\[115\] deser_A.kept_shift_reg\[116\] net734 VGND VGND
+ VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_4
X_0686_ _0418_ _0512_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__or2_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1238_ clknet_4_15_0_B_in_serial_clk _0186_ net15 VGND VGND VPWR VPWR deser_B.bit_idx\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1307_ clknet_4_0_0_B_in_serial_clk _0254_ net14 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_1169_ clknet_4_15_0_A_in_serial_clk _0117_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0540_ systolic_inst.cycle_cnt\[12\] systolic_inst.cycle_cnt\[13\] systolic_inst.cycle_cnt\[14\]
+ systolic_inst.cycle_cnt\[15\] VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_28_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1023_ _0381_ _0382_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nor2_1
XFILLER_61_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0738_ deser_A.kept_shift_reg\[29\] deser_A.kept_shift_reg\[30\] net17 VGND VGND
+ VPWR VPWR _0081_ sky130_fd_sc_hd__mux2_1
X_0807_ deser_A.kept_shift_reg\[98\] deser_A.kept_shift_reg\[99\] net647 VGND VGND
+ VPWR VPWR _0150_ sky130_fd_sc_hd__mux2_4
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0669_ net26 net494 net491 VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_3 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1006_ deser_B.kept_shift_reg\[125\] deser_B.kept_shift_reg\[126\] net27 VGND VGND
+ VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
Xrebuffer15 net816 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_6
Xrebuffer26 _0368_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1340_ clknet_4_7_0_B_in_serial_clk _0287_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer480 deser_A.bit_idx\[1\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer6 deser_A.receiving VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_8
X_1271_ clknet_4_10_0_B_in_serial_clk _0218_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0986_ deser_B.kept_shift_reg\[105\] deser_B.kept_shift_reg\[106\] net845 VGND VGND
+ VPWR VPWR _0301_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ net34 deser_B.bit_idx\[1\] net501 VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__and3_1
X_0771_ deser_A.kept_shift_reg\[62\] deser_A.kept_shift_reg\[63\] net809 VGND VGND
+ VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_4
X_1323_ clknet_4_4_0_B_in_serial_clk _0270_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1254_ clknet_4_12_0_B_in_serial_clk _0201_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1185_ clknet_4_1_0_A_in_serial_clk _0133_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0969_ deser_B.kept_shift_reg\[88\] deser_B.kept_shift_reg\[89\] net47 VGND VGND
+ VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0754_ deser_A.kept_shift_reg\[45\] deser_A.kept_shift_reg\[46\] net734 VGND VGND
+ VPWR VPWR _0097_ sky130_fd_sc_hd__mux2_4
X_0685_ _0417_ deser_A.bit_idx\[7\] _0501_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__and3_1
X_0823_ deser_A.kept_shift_reg\[114\] deser_A.kept_shift_reg\[115\] net734 VGND VGND
+ VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_4
X_1306_ clknet_4_1_0_B_in_serial_clk _0253_ net15 VGND VGND VPWR VPWR deser_B.kept_shift_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_1237_ clknet_4_15_0_B_in_serial_clk _0185_ net15 VGND VGND VPWR VPWR deser_B.bit_idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1168_ clknet_4_14_0_A_in_serial_clk _0116_ net14 VGND VGND VPWR VPWR deser_A.kept_shift_reg\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_1099_ clknet_4_9_0_A_in_serial_clk _0048_ net14 VGND VGND VPWR VPWR deser_A.kept_bit_idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclone792 net24 VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__buf_8
XFILLER_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1022_ ser_C.bit_idx\[3\] _0379_ ser_C.bit_idx\[4\] VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0668_ deser_A.receiving net1 VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__nand2b_4
X_0737_ deser_A.kept_shift_reg\[28\] deser_A.kept_shift_reg\[29\] net17 VGND VGND
+ VPWR VPWR _0080_ sky130_fd_sc_hd__mux2_1
X_0806_ deser_A.kept_shift_reg\[97\] deser_A.kept_shift_reg\[98\] net734 VGND VGND
+ VPWR VPWR _0149_ sky130_fd_sc_hd__mux2_4
XFILLER_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0599_ systolic_inst.cycle_cnt\[9\] systolic_inst.cycle_cnt\[10\] _0453_ systolic_inst.cycle_cnt\[11\]
+ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__a31o_1
XFILLER_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer832 deser_B.receiving VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_4_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_4 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer16 net31 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
Xrebuffer27 _0368_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1005_ deser_B.kept_shift_reg\[124\] deser_B.kept_shift_reg\[125\] net19 VGND VGND
+ VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

