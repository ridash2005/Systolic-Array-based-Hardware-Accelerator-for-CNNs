module Systolic4x4_serial_io (A_in_frame_sync,
    A_in_serial_clk,
    A_in_serial_data,
    B_in_frame_sync,
    B_in_serial_clk,
    B_in_serial_data,
    C_out_frame_sync,
    C_out_serial_clk,
    C_out_serial_data,
    clk,
    done,
    rst_n,
    start);
 input A_in_frame_sync;
 input A_in_serial_clk;
 input A_in_serial_data;
 input B_in_frame_sync;
 input B_in_serial_clk;
 input B_in_serial_data;
 output C_out_frame_sync;
 output C_out_serial_clk;
 output C_out_serial_data;
 input clk;
 output done;
 input rst_n;
 input start;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire \deser_A.bit_idx[0] ;
 wire \deser_A.bit_idx[1] ;
 wire \deser_A.bit_idx[2] ;
 wire \deser_A.bit_idx[3] ;
 wire \deser_A.bit_idx[4] ;
 wire \deser_A.bit_idx[5] ;
 wire \deser_A.bit_idx[6] ;
 wire \deser_A.bit_idx[7] ;
 wire \deser_A.kept_bit_idx[0] ;
 wire \deser_A.kept_bit_idx[1] ;
 wire \deser_A.kept_bit_idx[2] ;
 wire \deser_A.kept_bit_idx[3] ;
 wire \deser_A.kept_bit_idx[4] ;
 wire \deser_A.kept_bit_idx[5] ;
 wire \deser_A.kept_bit_idx[6] ;
 wire \deser_A.kept_bit_idx[7] ;
 wire \deser_A.kept_receiving ;
 wire \deser_A.kept_shift_reg[0] ;
 wire \deser_A.kept_shift_reg[100] ;
 wire \deser_A.kept_shift_reg[101] ;
 wire \deser_A.kept_shift_reg[102] ;
 wire \deser_A.kept_shift_reg[103] ;
 wire \deser_A.kept_shift_reg[104] ;
 wire \deser_A.kept_shift_reg[105] ;
 wire \deser_A.kept_shift_reg[106] ;
 wire \deser_A.kept_shift_reg[107] ;
 wire \deser_A.kept_shift_reg[108] ;
 wire \deser_A.kept_shift_reg[109] ;
 wire \deser_A.kept_shift_reg[10] ;
 wire \deser_A.kept_shift_reg[110] ;
 wire \deser_A.kept_shift_reg[111] ;
 wire \deser_A.kept_shift_reg[112] ;
 wire \deser_A.kept_shift_reg[113] ;
 wire \deser_A.kept_shift_reg[114] ;
 wire \deser_A.kept_shift_reg[115] ;
 wire \deser_A.kept_shift_reg[116] ;
 wire \deser_A.kept_shift_reg[117] ;
 wire \deser_A.kept_shift_reg[118] ;
 wire \deser_A.kept_shift_reg[119] ;
 wire \deser_A.kept_shift_reg[11] ;
 wire \deser_A.kept_shift_reg[120] ;
 wire \deser_A.kept_shift_reg[121] ;
 wire \deser_A.kept_shift_reg[122] ;
 wire \deser_A.kept_shift_reg[123] ;
 wire \deser_A.kept_shift_reg[124] ;
 wire \deser_A.kept_shift_reg[125] ;
 wire \deser_A.kept_shift_reg[126] ;
 wire \deser_A.kept_shift_reg[127] ;
 wire \deser_A.kept_shift_reg[12] ;
 wire \deser_A.kept_shift_reg[13] ;
 wire \deser_A.kept_shift_reg[14] ;
 wire \deser_A.kept_shift_reg[15] ;
 wire \deser_A.kept_shift_reg[16] ;
 wire \deser_A.kept_shift_reg[17] ;
 wire \deser_A.kept_shift_reg[18] ;
 wire \deser_A.kept_shift_reg[19] ;
 wire \deser_A.kept_shift_reg[1] ;
 wire \deser_A.kept_shift_reg[20] ;
 wire \deser_A.kept_shift_reg[21] ;
 wire \deser_A.kept_shift_reg[22] ;
 wire \deser_A.kept_shift_reg[23] ;
 wire \deser_A.kept_shift_reg[24] ;
 wire \deser_A.kept_shift_reg[25] ;
 wire \deser_A.kept_shift_reg[26] ;
 wire \deser_A.kept_shift_reg[27] ;
 wire \deser_A.kept_shift_reg[28] ;
 wire \deser_A.kept_shift_reg[29] ;
 wire \deser_A.kept_shift_reg[2] ;
 wire \deser_A.kept_shift_reg[30] ;
 wire \deser_A.kept_shift_reg[31] ;
 wire \deser_A.kept_shift_reg[32] ;
 wire \deser_A.kept_shift_reg[33] ;
 wire \deser_A.kept_shift_reg[34] ;
 wire \deser_A.kept_shift_reg[35] ;
 wire \deser_A.kept_shift_reg[36] ;
 wire \deser_A.kept_shift_reg[37] ;
 wire \deser_A.kept_shift_reg[38] ;
 wire \deser_A.kept_shift_reg[39] ;
 wire \deser_A.kept_shift_reg[3] ;
 wire \deser_A.kept_shift_reg[40] ;
 wire \deser_A.kept_shift_reg[41] ;
 wire \deser_A.kept_shift_reg[42] ;
 wire \deser_A.kept_shift_reg[43] ;
 wire \deser_A.kept_shift_reg[44] ;
 wire \deser_A.kept_shift_reg[45] ;
 wire \deser_A.kept_shift_reg[46] ;
 wire \deser_A.kept_shift_reg[47] ;
 wire \deser_A.kept_shift_reg[48] ;
 wire \deser_A.kept_shift_reg[49] ;
 wire \deser_A.kept_shift_reg[4] ;
 wire \deser_A.kept_shift_reg[50] ;
 wire \deser_A.kept_shift_reg[51] ;
 wire \deser_A.kept_shift_reg[52] ;
 wire \deser_A.kept_shift_reg[53] ;
 wire \deser_A.kept_shift_reg[54] ;
 wire \deser_A.kept_shift_reg[55] ;
 wire \deser_A.kept_shift_reg[56] ;
 wire \deser_A.kept_shift_reg[57] ;
 wire \deser_A.kept_shift_reg[58] ;
 wire \deser_A.kept_shift_reg[59] ;
 wire \deser_A.kept_shift_reg[5] ;
 wire \deser_A.kept_shift_reg[60] ;
 wire \deser_A.kept_shift_reg[61] ;
 wire \deser_A.kept_shift_reg[62] ;
 wire \deser_A.kept_shift_reg[63] ;
 wire \deser_A.kept_shift_reg[64] ;
 wire \deser_A.kept_shift_reg[65] ;
 wire \deser_A.kept_shift_reg[66] ;
 wire \deser_A.kept_shift_reg[67] ;
 wire \deser_A.kept_shift_reg[68] ;
 wire \deser_A.kept_shift_reg[69] ;
 wire \deser_A.kept_shift_reg[6] ;
 wire \deser_A.kept_shift_reg[70] ;
 wire \deser_A.kept_shift_reg[71] ;
 wire \deser_A.kept_shift_reg[72] ;
 wire \deser_A.kept_shift_reg[73] ;
 wire \deser_A.kept_shift_reg[74] ;
 wire \deser_A.kept_shift_reg[75] ;
 wire \deser_A.kept_shift_reg[76] ;
 wire \deser_A.kept_shift_reg[77] ;
 wire \deser_A.kept_shift_reg[78] ;
 wire \deser_A.kept_shift_reg[79] ;
 wire \deser_A.kept_shift_reg[7] ;
 wire \deser_A.kept_shift_reg[80] ;
 wire \deser_A.kept_shift_reg[81] ;
 wire \deser_A.kept_shift_reg[82] ;
 wire \deser_A.kept_shift_reg[83] ;
 wire \deser_A.kept_shift_reg[84] ;
 wire \deser_A.kept_shift_reg[85] ;
 wire \deser_A.kept_shift_reg[86] ;
 wire \deser_A.kept_shift_reg[87] ;
 wire \deser_A.kept_shift_reg[88] ;
 wire \deser_A.kept_shift_reg[89] ;
 wire \deser_A.kept_shift_reg[8] ;
 wire \deser_A.kept_shift_reg[90] ;
 wire \deser_A.kept_shift_reg[91] ;
 wire \deser_A.kept_shift_reg[92] ;
 wire \deser_A.kept_shift_reg[93] ;
 wire \deser_A.kept_shift_reg[94] ;
 wire \deser_A.kept_shift_reg[95] ;
 wire \deser_A.kept_shift_reg[96] ;
 wire \deser_A.kept_shift_reg[97] ;
 wire \deser_A.kept_shift_reg[98] ;
 wire \deser_A.kept_shift_reg[99] ;
 wire \deser_A.kept_shift_reg[9] ;
 wire \deser_A.receiving ;
 wire \deser_B.bit_idx[0] ;
 wire \deser_B.bit_idx[1] ;
 wire \deser_B.bit_idx[2] ;
 wire \deser_B.bit_idx[3] ;
 wire \deser_B.bit_idx[4] ;
 wire \deser_B.bit_idx[5] ;
 wire \deser_B.bit_idx[6] ;
 wire \deser_B.bit_idx[7] ;
 wire \deser_B.kept_bit_idx[0] ;
 wire \deser_B.kept_bit_idx[1] ;
 wire \deser_B.kept_bit_idx[2] ;
 wire \deser_B.kept_bit_idx[3] ;
 wire \deser_B.kept_bit_idx[4] ;
 wire \deser_B.kept_bit_idx[5] ;
 wire \deser_B.kept_bit_idx[6] ;
 wire \deser_B.kept_bit_idx[7] ;
 wire \deser_B.kept_receiving ;
 wire \deser_B.kept_shift_reg[0] ;
 wire \deser_B.kept_shift_reg[100] ;
 wire \deser_B.kept_shift_reg[101] ;
 wire \deser_B.kept_shift_reg[102] ;
 wire \deser_B.kept_shift_reg[103] ;
 wire \deser_B.kept_shift_reg[104] ;
 wire \deser_B.kept_shift_reg[105] ;
 wire \deser_B.kept_shift_reg[106] ;
 wire \deser_B.kept_shift_reg[107] ;
 wire \deser_B.kept_shift_reg[108] ;
 wire \deser_B.kept_shift_reg[109] ;
 wire \deser_B.kept_shift_reg[10] ;
 wire \deser_B.kept_shift_reg[110] ;
 wire \deser_B.kept_shift_reg[111] ;
 wire \deser_B.kept_shift_reg[112] ;
 wire \deser_B.kept_shift_reg[113] ;
 wire \deser_B.kept_shift_reg[114] ;
 wire \deser_B.kept_shift_reg[115] ;
 wire \deser_B.kept_shift_reg[116] ;
 wire \deser_B.kept_shift_reg[117] ;
 wire \deser_B.kept_shift_reg[118] ;
 wire \deser_B.kept_shift_reg[119] ;
 wire \deser_B.kept_shift_reg[11] ;
 wire \deser_B.kept_shift_reg[120] ;
 wire \deser_B.kept_shift_reg[121] ;
 wire \deser_B.kept_shift_reg[122] ;
 wire \deser_B.kept_shift_reg[123] ;
 wire \deser_B.kept_shift_reg[124] ;
 wire \deser_B.kept_shift_reg[125] ;
 wire \deser_B.kept_shift_reg[126] ;
 wire \deser_B.kept_shift_reg[127] ;
 wire \deser_B.kept_shift_reg[12] ;
 wire \deser_B.kept_shift_reg[13] ;
 wire \deser_B.kept_shift_reg[14] ;
 wire \deser_B.kept_shift_reg[15] ;
 wire \deser_B.kept_shift_reg[16] ;
 wire \deser_B.kept_shift_reg[17] ;
 wire \deser_B.kept_shift_reg[18] ;
 wire \deser_B.kept_shift_reg[19] ;
 wire \deser_B.kept_shift_reg[1] ;
 wire \deser_B.kept_shift_reg[20] ;
 wire \deser_B.kept_shift_reg[21] ;
 wire \deser_B.kept_shift_reg[22] ;
 wire \deser_B.kept_shift_reg[23] ;
 wire \deser_B.kept_shift_reg[24] ;
 wire \deser_B.kept_shift_reg[25] ;
 wire \deser_B.kept_shift_reg[26] ;
 wire \deser_B.kept_shift_reg[27] ;
 wire \deser_B.kept_shift_reg[28] ;
 wire \deser_B.kept_shift_reg[29] ;
 wire \deser_B.kept_shift_reg[2] ;
 wire \deser_B.kept_shift_reg[30] ;
 wire \deser_B.kept_shift_reg[31] ;
 wire \deser_B.kept_shift_reg[32] ;
 wire \deser_B.kept_shift_reg[33] ;
 wire \deser_B.kept_shift_reg[34] ;
 wire \deser_B.kept_shift_reg[35] ;
 wire \deser_B.kept_shift_reg[36] ;
 wire \deser_B.kept_shift_reg[37] ;
 wire \deser_B.kept_shift_reg[38] ;
 wire \deser_B.kept_shift_reg[39] ;
 wire \deser_B.kept_shift_reg[3] ;
 wire \deser_B.kept_shift_reg[40] ;
 wire \deser_B.kept_shift_reg[41] ;
 wire \deser_B.kept_shift_reg[42] ;
 wire \deser_B.kept_shift_reg[43] ;
 wire \deser_B.kept_shift_reg[44] ;
 wire \deser_B.kept_shift_reg[45] ;
 wire \deser_B.kept_shift_reg[46] ;
 wire \deser_B.kept_shift_reg[47] ;
 wire \deser_B.kept_shift_reg[48] ;
 wire \deser_B.kept_shift_reg[49] ;
 wire \deser_B.kept_shift_reg[4] ;
 wire \deser_B.kept_shift_reg[50] ;
 wire \deser_B.kept_shift_reg[51] ;
 wire \deser_B.kept_shift_reg[52] ;
 wire \deser_B.kept_shift_reg[53] ;
 wire \deser_B.kept_shift_reg[54] ;
 wire \deser_B.kept_shift_reg[55] ;
 wire \deser_B.kept_shift_reg[56] ;
 wire \deser_B.kept_shift_reg[57] ;
 wire \deser_B.kept_shift_reg[58] ;
 wire \deser_B.kept_shift_reg[59] ;
 wire \deser_B.kept_shift_reg[5] ;
 wire \deser_B.kept_shift_reg[60] ;
 wire \deser_B.kept_shift_reg[61] ;
 wire \deser_B.kept_shift_reg[62] ;
 wire \deser_B.kept_shift_reg[63] ;
 wire \deser_B.kept_shift_reg[64] ;
 wire \deser_B.kept_shift_reg[65] ;
 wire \deser_B.kept_shift_reg[66] ;
 wire \deser_B.kept_shift_reg[67] ;
 wire \deser_B.kept_shift_reg[68] ;
 wire \deser_B.kept_shift_reg[69] ;
 wire \deser_B.kept_shift_reg[6] ;
 wire \deser_B.kept_shift_reg[70] ;
 wire \deser_B.kept_shift_reg[71] ;
 wire \deser_B.kept_shift_reg[72] ;
 wire \deser_B.kept_shift_reg[73] ;
 wire \deser_B.kept_shift_reg[74] ;
 wire \deser_B.kept_shift_reg[75] ;
 wire \deser_B.kept_shift_reg[76] ;
 wire \deser_B.kept_shift_reg[77] ;
 wire \deser_B.kept_shift_reg[78] ;
 wire \deser_B.kept_shift_reg[79] ;
 wire \deser_B.kept_shift_reg[7] ;
 wire \deser_B.kept_shift_reg[80] ;
 wire \deser_B.kept_shift_reg[81] ;
 wire \deser_B.kept_shift_reg[82] ;
 wire \deser_B.kept_shift_reg[83] ;
 wire \deser_B.kept_shift_reg[84] ;
 wire \deser_B.kept_shift_reg[85] ;
 wire \deser_B.kept_shift_reg[86] ;
 wire \deser_B.kept_shift_reg[87] ;
 wire \deser_B.kept_shift_reg[88] ;
 wire \deser_B.kept_shift_reg[89] ;
 wire \deser_B.kept_shift_reg[8] ;
 wire \deser_B.kept_shift_reg[90] ;
 wire \deser_B.kept_shift_reg[91] ;
 wire \deser_B.kept_shift_reg[92] ;
 wire \deser_B.kept_shift_reg[93] ;
 wire \deser_B.kept_shift_reg[94] ;
 wire \deser_B.kept_shift_reg[95] ;
 wire \deser_B.kept_shift_reg[96] ;
 wire \deser_B.kept_shift_reg[97] ;
 wire \deser_B.kept_shift_reg[98] ;
 wire \deser_B.kept_shift_reg[99] ;
 wire \deser_B.kept_shift_reg[9] ;
 wire \deser_B.receiving ;
 wire \ser_C.bit_idx[0] ;
 wire \ser_C.bit_idx[1] ;
 wire \ser_C.bit_idx[2] ;
 wire \ser_C.bit_idx[3] ;
 wire \ser_C.bit_idx[4] ;
 wire \ser_C.bit_idx[5] ;
 wire \ser_C.bit_idx[6] ;
 wire \ser_C.bit_idx[7] ;
 wire \ser_C.bit_idx[8] ;
 wire \ser_C.bit_idx[9] ;
 wire \ser_C.kept_bit_idx[0] ;
 wire \ser_C.kept_bit_idx[1] ;
 wire \ser_C.kept_bit_idx[2] ;
 wire \ser_C.kept_bit_idx[3] ;
 wire \ser_C.kept_bit_idx[4] ;
 wire \ser_C.kept_bit_idx[5] ;
 wire \ser_C.kept_bit_idx[6] ;
 wire \ser_C.kept_bit_idx[7] ;
 wire \ser_C.kept_bit_idx[8] ;
 wire \ser_C.kept_bit_idx[9] ;
 wire clknet_4_15_0_B_in_serial_clk;
 wire clknet_4_14_0_B_in_serial_clk;
 wire clknet_4_13_0_B_in_serial_clk;
 wire clknet_4_12_0_B_in_serial_clk;
 wire clknet_4_11_0_B_in_serial_clk;
 wire clknet_4_10_0_B_in_serial_clk;
 wire clknet_4_9_0_B_in_serial_clk;
 wire clknet_4_8_0_B_in_serial_clk;
 wire clknet_4_7_0_B_in_serial_clk;
 wire clknet_4_6_0_B_in_serial_clk;
 wire clknet_4_5_0_B_in_serial_clk;
 wire clknet_4_4_0_B_in_serial_clk;
 wire clknet_4_3_0_B_in_serial_clk;
 wire clknet_4_2_0_B_in_serial_clk;
 wire clknet_4_1_0_B_in_serial_clk;
 wire clknet_4_0_0_B_in_serial_clk;
 wire clknet_0_B_in_serial_clk;
 wire clknet_4_15_0_A_in_serial_clk;
 wire clknet_4_14_0_A_in_serial_clk;
 wire clknet_4_13_0_A_in_serial_clk;
 wire clknet_4_12_0_A_in_serial_clk;
 wire clknet_4_11_0_A_in_serial_clk;
 wire clknet_4_10_0_A_in_serial_clk;
 wire clknet_4_9_0_A_in_serial_clk;
 wire clknet_4_8_0_A_in_serial_clk;
 wire clknet_4_7_0_A_in_serial_clk;
 wire clknet_4_6_0_A_in_serial_clk;
 wire clknet_4_5_0_A_in_serial_clk;
 wire clknet_4_4_0_A_in_serial_clk;
 wire clknet_4_3_0_A_in_serial_clk;
 wire clknet_4_2_0_A_in_serial_clk;
 wire clknet_4_1_0_A_in_serial_clk;
 wire clknet_4_0_0_A_in_serial_clk;
 wire clknet_0_A_in_serial_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_0_clk;
 wire \systolic_inst.ce_local ;
 wire \systolic_inst.cycle_cnt[0] ;
 wire \systolic_inst.cycle_cnt[10] ;
 wire \systolic_inst.cycle_cnt[11] ;
 wire \systolic_inst.cycle_cnt[12] ;
 wire \systolic_inst.cycle_cnt[13] ;
 wire \systolic_inst.cycle_cnt[14] ;
 wire \systolic_inst.cycle_cnt[15] ;
 wire \systolic_inst.cycle_cnt[16] ;
 wire \systolic_inst.cycle_cnt[17] ;
 wire \systolic_inst.cycle_cnt[18] ;
 wire \systolic_inst.cycle_cnt[19] ;
 wire \systolic_inst.cycle_cnt[1] ;
 wire \systolic_inst.cycle_cnt[20] ;
 wire \systolic_inst.cycle_cnt[21] ;
 wire \systolic_inst.cycle_cnt[22] ;
 wire \systolic_inst.cycle_cnt[23] ;
 wire \systolic_inst.cycle_cnt[24] ;
 wire \systolic_inst.cycle_cnt[25] ;
 wire \systolic_inst.cycle_cnt[26] ;
 wire \systolic_inst.cycle_cnt[27] ;
 wire \systolic_inst.cycle_cnt[28] ;
 wire \systolic_inst.cycle_cnt[29] ;
 wire \systolic_inst.cycle_cnt[2] ;
 wire \systolic_inst.cycle_cnt[30] ;
 wire \systolic_inst.cycle_cnt[31] ;
 wire \systolic_inst.cycle_cnt[3] ;
 wire \systolic_inst.cycle_cnt[4] ;
 wire \systolic_inst.cycle_cnt[5] ;
 wire \systolic_inst.cycle_cnt[6] ;
 wire \systolic_inst.cycle_cnt[7] ;
 wire \systolic_inst.cycle_cnt[8] ;
 wire \systolic_inst.cycle_cnt[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;

 sky130_fd_sc_hd__inv_2 _0528_ (.A(\systolic_inst.cycle_cnt[23] ),
    .Y(_0399_));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(\systolic_inst.cycle_cnt[30] ),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(\systolic_inst.cycle_cnt[31] ),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_2 _0531_ (.A(net7),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(\deser_A.kept_receiving ),
    .Y(_0403_));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(\deser_B.kept_receiving ),
    .Y(_0404_));
 sky130_fd_sc_hd__or4_1 _0534_ (.A(\systolic_inst.cycle_cnt[24] ),
    .B(\systolic_inst.cycle_cnt[25] ),
    .C(\systolic_inst.cycle_cnt[26] ),
    .D(\systolic_inst.cycle_cnt[27] ),
    .X(_0405_));
 sky130_fd_sc_hd__or4_1 _0535_ (.A(\systolic_inst.cycle_cnt[20] ),
    .B(\systolic_inst.cycle_cnt[21] ),
    .C(\systolic_inst.cycle_cnt[22] ),
    .D(\systolic_inst.cycle_cnt[23] ),
    .X(_0406_));
 sky130_fd_sc_hd__or4_1 _0536_ (.A(\systolic_inst.cycle_cnt[28] ),
    .B(\systolic_inst.cycle_cnt[29] ),
    .C(\systolic_inst.cycle_cnt[30] ),
    .D(\systolic_inst.cycle_cnt[31] ),
    .X(_0407_));
 sky130_fd_sc_hd__o21a_1 _0537_ (.A1(\systolic_inst.cycle_cnt[1] ),
    .A2(\systolic_inst.cycle_cnt[2] ),
    .B1(\systolic_inst.cycle_cnt[3] ),
    .X(_0408_));
 sky130_fd_sc_hd__or3_1 _0538_ (.A(\systolic_inst.cycle_cnt[8] ),
    .B(\systolic_inst.cycle_cnt[9] ),
    .C(\systolic_inst.cycle_cnt[10] ),
    .X(_0409_));
 sky130_fd_sc_hd__or4_1 _0539_ (.A(\systolic_inst.cycle_cnt[4] ),
    .B(\systolic_inst.cycle_cnt[5] ),
    .C(\systolic_inst.cycle_cnt[6] ),
    .D(\systolic_inst.cycle_cnt[7] ),
    .X(_0410_));
 sky130_fd_sc_hd__or4_1 _0540_ (.A(\systolic_inst.cycle_cnt[12] ),
    .B(\systolic_inst.cycle_cnt[13] ),
    .C(\systolic_inst.cycle_cnt[14] ),
    .D(\systolic_inst.cycle_cnt[15] ),
    .X(_0411_));
 sky130_fd_sc_hd__or4_1 _0541_ (.A(\systolic_inst.cycle_cnt[16] ),
    .B(\systolic_inst.cycle_cnt[17] ),
    .C(\systolic_inst.cycle_cnt[18] ),
    .D(\systolic_inst.cycle_cnt[19] ),
    .X(_0412_));
 sky130_fd_sc_hd__or4_1 _0542_ (.A(_0405_),
    .B(_0406_),
    .C(_0407_),
    .D(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__or4_1 _0543_ (.A(_0408_),
    .B(_0409_),
    .C(_0410_),
    .D(_0411_),
    .X(_0414_));
 sky130_fd_sc_hd__o31a_1 _0544_ (.A1(\systolic_inst.cycle_cnt[11] ),
    .A2(_0413_),
    .A3(_0414_),
    .B1(\systolic_inst.ce_local ),
    .X(_0003_));
 sky130_fd_sc_hd__and4_1 _0545_ (.A(\deser_A.bit_idx[1] ),
    .B(\deser_A.bit_idx[0] ),
    .C(\deser_A.bit_idx[3] ),
    .D(\deser_A.bit_idx[2] ),
    .X(_0415_));
 sky130_fd_sc_hd__and2_1 _0546_ (.A(\deser_A.bit_idx[4] ),
    .B(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__nand4_1 _0547_ (.A(\deser_A.receiving ),
    .B(\deser_A.bit_idx[5] ),
    .C(\deser_A.bit_idx[6] ),
    .D(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__nor2_1 _0548_ (.A(\deser_A.bit_idx[7] ),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_1 _0549_ (.A(net1),
    .B(\deser_A.receiving ),
    .Y(_0419_));
 sky130_fd_sc_hd__or2_2 _0550_ (.A(net1),
    .B(\deser_A.receiving ),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_1 _0551_ (.A(_0418_),
    .B(_0419_),
    .Y(_0000_));
 sky130_fd_sc_hd__and4_1 _0552_ (.A(\deser_B.bit_idx[1] ),
    .B(\deser_B.bit_idx[0] ),
    .C(\deser_B.bit_idx[3] ),
    .D(\deser_B.bit_idx[2] ),
    .X(_0421_));
 sky130_fd_sc_hd__and2_1 _0553_ (.A(\deser_B.bit_idx[4] ),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__nand4_1 _0554_ (.A(\deser_B.receiving ),
    .B(\deser_B.bit_idx[5] ),
    .C(\deser_B.bit_idx[6] ),
    .D(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__nor2_1 _0555_ (.A(\deser_B.bit_idx[7] ),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nor2_1 _0556_ (.A(net3),
    .B(\deser_B.receiving ),
    .Y(_0425_));
 sky130_fd_sc_hd__or2_2 _0557_ (.A(net3),
    .B(\deser_B.receiving ),
    .X(_0426_));
 sky130_fd_sc_hd__nor2_1 _0558_ (.A(_0424_),
    .B(_0425_),
    .Y(_0001_));
 sky130_fd_sc_hd__nor2_1 _0559_ (.A(net6),
    .B(\systolic_inst.ce_local ),
    .Y(_0427_));
 sky130_fd_sc_hd__or2_1 _0560_ (.A(net6),
    .B(\systolic_inst.ce_local ),
    .X(_0428_));
 sky130_fd_sc_hd__nor2_1 _0561_ (.A(_0003_),
    .B(_0427_),
    .Y(_0004_));
 sky130_fd_sc_hd__and4b_1 _0562_ (.A_N(\ser_C.bit_idx[9] ),
    .B(\ser_C.bit_idx[8] ),
    .C(\ser_C.bit_idx[7] ),
    .D(\ser_C.bit_idx[6] ),
    .X(_0429_));
 sky130_fd_sc_hd__and4_1 _0563_ (.A(\ser_C.bit_idx[0] ),
    .B(\ser_C.bit_idx[1] ),
    .C(\ser_C.bit_idx[2] ),
    .D(\ser_C.bit_idx[3] ),
    .X(_0430_));
 sky130_fd_sc_hd__a41o_1 _0564_ (.A1(\ser_C.bit_idx[5] ),
    .A2(\ser_C.bit_idx[4] ),
    .A3(_0429_),
    .A4(_0430_),
    .B1(_0402_),
    .X(_0431_));
 sky130_fd_sc_hd__inv_2 _0565_ (.A(_0431_),
    .Y(_0002_));
 sky130_fd_sc_hd__mux2_1 _0566_ (.A0(\systolic_inst.ce_local ),
    .A1(_0427_),
    .S(\systolic_inst.cycle_cnt[0] ),
    .X(_0005_));
 sky130_fd_sc_hd__a21o_1 _0567_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.cycle_cnt[0] ),
    .B1(\systolic_inst.cycle_cnt[1] ),
    .X(_0432_));
 sky130_fd_sc_hd__and2_1 _0568_ (.A(\systolic_inst.cycle_cnt[0] ),
    .B(\systolic_inst.cycle_cnt[1] ),
    .X(_0433_));
 sky130_fd_sc_hd__and3_1 _0569_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.cycle_cnt[0] ),
    .C(\systolic_inst.cycle_cnt[1] ),
    .X(_0434_));
 sky130_fd_sc_hd__and2b_2 _0570_ (.A_N(\systolic_inst.ce_local ),
    .B(net6),
    .X(_0435_));
 sky130_fd_sc_hd__nand2b_4 _0571_ (.A_N(\systolic_inst.ce_local ),
    .B(net6),
    .Y(_0436_));
 sky130_fd_sc_hd__nor2_1 _0572_ (.A(_0434_),
    .B(_0435_),
    .Y(_0437_));
 sky130_fd_sc_hd__and2_1 _0573_ (.A(_0432_),
    .B(_0437_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0574_ (.A0(_0434_),
    .A1(_0437_),
    .S(\systolic_inst.cycle_cnt[2] ),
    .X(_0007_));
 sky130_fd_sc_hd__a31o_1 _0575_ (.A1(\systolic_inst.cycle_cnt[2] ),
    .A2(_0428_),
    .A3(_0433_),
    .B1(\systolic_inst.cycle_cnt[3] ),
    .X(_0438_));
 sky130_fd_sc_hd__and3_1 _0576_ (.A(\systolic_inst.cycle_cnt[2] ),
    .B(\systolic_inst.cycle_cnt[3] ),
    .C(_0434_),
    .X(_0439_));
 sky130_fd_sc_hd__nor2_1 _0577_ (.A(_0435_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__and2_1 _0578_ (.A(_0438_),
    .B(_0440_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0579_ (.A0(_0439_),
    .A1(_0440_),
    .S(\systolic_inst.cycle_cnt[4] ),
    .X(_0009_));
 sky130_fd_sc_hd__and3_1 _0580_ (.A(\systolic_inst.cycle_cnt[2] ),
    .B(\systolic_inst.cycle_cnt[3] ),
    .C(\systolic_inst.cycle_cnt[4] ),
    .X(_0441_));
 sky130_fd_sc_hd__and3_1 _0581_ (.A(\systolic_inst.cycle_cnt[5] ),
    .B(_0434_),
    .C(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__nor2_1 _0582_ (.A(_0435_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__and3_1 _0583_ (.A(_0428_),
    .B(_0433_),
    .C(_0441_),
    .X(_0444_));
 sky130_fd_sc_hd__o21a_1 _0584_ (.A1(\systolic_inst.cycle_cnt[5] ),
    .A2(_0444_),
    .B1(_0443_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(_0442_),
    .A1(_0443_),
    .S(\systolic_inst.cycle_cnt[6] ),
    .X(_0011_));
 sky130_fd_sc_hd__a31o_1 _0586_ (.A1(\systolic_inst.cycle_cnt[5] ),
    .A2(\systolic_inst.cycle_cnt[6] ),
    .A3(_0444_),
    .B1(\systolic_inst.cycle_cnt[7] ),
    .X(_0445_));
 sky130_fd_sc_hd__and3_1 _0587_ (.A(\systolic_inst.cycle_cnt[5] ),
    .B(\systolic_inst.cycle_cnt[6] ),
    .C(\systolic_inst.cycle_cnt[7] ),
    .X(_0446_));
 sky130_fd_sc_hd__and3_1 _0588_ (.A(_0433_),
    .B(_0441_),
    .C(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__and4_2 _0589_ (.A(\systolic_inst.ce_local ),
    .B(_0433_),
    .C(_0441_),
    .D(_0446_),
    .X(_0448_));
 sky130_fd_sc_hd__inv_2 _0590_ (.A(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__and3_1 _0591_ (.A(_0436_),
    .B(_0445_),
    .C(_0449_),
    .X(_0012_));
 sky130_fd_sc_hd__a21oi_1 _0592_ (.A1(\systolic_inst.cycle_cnt[8] ),
    .A2(_0436_),
    .B1(_0448_),
    .Y(_0450_));
 sky130_fd_sc_hd__a21oi_1 _0593_ (.A1(\systolic_inst.cycle_cnt[8] ),
    .A2(_0448_),
    .B1(_0450_),
    .Y(_0013_));
 sky130_fd_sc_hd__and3_1 _0594_ (.A(\systolic_inst.cycle_cnt[8] ),
    .B(\systolic_inst.cycle_cnt[9] ),
    .C(_0448_),
    .X(_0451_));
 sky130_fd_sc_hd__nor2_1 _0595_ (.A(_0435_),
    .B(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__and3_1 _0596_ (.A(\systolic_inst.cycle_cnt[8] ),
    .B(_0428_),
    .C(_0447_),
    .X(_0453_));
 sky130_fd_sc_hd__o21a_1 _0597_ (.A1(\systolic_inst.cycle_cnt[9] ),
    .A2(_0453_),
    .B1(_0452_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0598_ (.A0(_0451_),
    .A1(_0452_),
    .S(\systolic_inst.cycle_cnt[10] ),
    .X(_0015_));
 sky130_fd_sc_hd__a31o_1 _0599_ (.A1(\systolic_inst.cycle_cnt[9] ),
    .A2(\systolic_inst.cycle_cnt[10] ),
    .A3(_0453_),
    .B1(\systolic_inst.cycle_cnt[11] ),
    .X(_0454_));
 sky130_fd_sc_hd__and4_1 _0600_ (.A(\systolic_inst.cycle_cnt[8] ),
    .B(\systolic_inst.cycle_cnt[9] ),
    .C(\systolic_inst.cycle_cnt[10] ),
    .D(\systolic_inst.cycle_cnt[11] ),
    .X(_0455_));
 sky130_fd_sc_hd__and2_1 _0601_ (.A(_0448_),
    .B(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__inv_2 _0602_ (.A(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__and3_1 _0603_ (.A(_0436_),
    .B(_0454_),
    .C(_0457_),
    .X(_0016_));
 sky130_fd_sc_hd__nand2_1 _0604_ (.A(\systolic_inst.cycle_cnt[12] ),
    .B(_0436_),
    .Y(_0458_));
 sky130_fd_sc_hd__mux2_1 _0605_ (.A0(_0458_),
    .A1(\systolic_inst.cycle_cnt[12] ),
    .S(_0456_),
    .X(_0459_));
 sky130_fd_sc_hd__inv_2 _0606_ (.A(_0459_),
    .Y(_0017_));
 sky130_fd_sc_hd__a22oi_1 _0607_ (.A1(\systolic_inst.cycle_cnt[13] ),
    .A2(_0436_),
    .B1(_0456_),
    .B2(\systolic_inst.cycle_cnt[12] ),
    .Y(_0460_));
 sky130_fd_sc_hd__and4_1 _0608_ (.A(\systolic_inst.cycle_cnt[12] ),
    .B(\systolic_inst.cycle_cnt[13] ),
    .C(_0448_),
    .D(_0455_),
    .X(_0461_));
 sky130_fd_sc_hd__nor2_1 _0609_ (.A(_0460_),
    .B(_0461_),
    .Y(_0018_));
 sky130_fd_sc_hd__a21oi_1 _0610_ (.A1(\systolic_inst.cycle_cnt[14] ),
    .A2(_0436_),
    .B1(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__and3_1 _0611_ (.A(\systolic_inst.cycle_cnt[12] ),
    .B(\systolic_inst.cycle_cnt[13] ),
    .C(\systolic_inst.cycle_cnt[14] ),
    .X(_0463_));
 sky130_fd_sc_hd__a21oi_1 _0612_ (.A1(\systolic_inst.cycle_cnt[14] ),
    .A2(_0461_),
    .B1(_0462_),
    .Y(_0019_));
 sky130_fd_sc_hd__and3_1 _0613_ (.A(\systolic_inst.cycle_cnt[15] ),
    .B(_0455_),
    .C(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__and2_1 _0614_ (.A(_0448_),
    .B(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__nor2_1 _0615_ (.A(_0435_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__and3b_1 _0616_ (.A_N(_0465_),
    .B(_0463_),
    .C(_0456_),
    .X(_0467_));
 sky130_fd_sc_hd__a21o_1 _0617_ (.A1(\systolic_inst.cycle_cnt[15] ),
    .A2(_0466_),
    .B1(_0467_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0618_ (.A0(_0465_),
    .A1(_0466_),
    .S(\systolic_inst.cycle_cnt[16] ),
    .X(_0021_));
 sky130_fd_sc_hd__and3_1 _0619_ (.A(\systolic_inst.cycle_cnt[16] ),
    .B(\systolic_inst.cycle_cnt[17] ),
    .C(_0465_),
    .X(_0468_));
 sky130_fd_sc_hd__a31oi_1 _0620_ (.A1(\systolic_inst.cycle_cnt[16] ),
    .A2(\systolic_inst.cycle_cnt[17] ),
    .A3(_0465_),
    .B1(_0435_),
    .Y(_0469_));
 sky130_fd_sc_hd__and3_1 _0621_ (.A(_0428_),
    .B(_0447_),
    .C(_0464_),
    .X(_0470_));
 sky130_fd_sc_hd__a21o_1 _0622_ (.A1(\systolic_inst.cycle_cnt[16] ),
    .A2(_0470_),
    .B1(\systolic_inst.cycle_cnt[17] ),
    .X(_0471_));
 sky130_fd_sc_hd__and2_1 _0623_ (.A(_0469_),
    .B(_0471_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0624_ (.A0(_0468_),
    .A1(_0469_),
    .S(\systolic_inst.cycle_cnt[18] ),
    .X(_0023_));
 sky130_fd_sc_hd__a41o_1 _0625_ (.A1(\systolic_inst.cycle_cnt[16] ),
    .A2(\systolic_inst.cycle_cnt[17] ),
    .A3(\systolic_inst.cycle_cnt[18] ),
    .A4(_0470_),
    .B1(\systolic_inst.cycle_cnt[19] ),
    .X(_0472_));
 sky130_fd_sc_hd__and4_1 _0626_ (.A(\systolic_inst.cycle_cnt[16] ),
    .B(\systolic_inst.cycle_cnt[17] ),
    .C(\systolic_inst.cycle_cnt[18] ),
    .D(\systolic_inst.cycle_cnt[19] ),
    .X(_0473_));
 sky130_fd_sc_hd__and3_1 _0627_ (.A(_0448_),
    .B(_0464_),
    .C(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_1 _0628_ (.A(_0435_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__and2_1 _0629_ (.A(_0472_),
    .B(_0475_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(_0474_),
    .A1(_0475_),
    .S(\systolic_inst.cycle_cnt[20] ),
    .X(_0025_));
 sky130_fd_sc_hd__a31o_1 _0631_ (.A1(\systolic_inst.cycle_cnt[20] ),
    .A2(_0470_),
    .A3(_0473_),
    .B1(\systolic_inst.cycle_cnt[21] ),
    .X(_0476_));
 sky130_fd_sc_hd__nand3_1 _0632_ (.A(\systolic_inst.cycle_cnt[20] ),
    .B(\systolic_inst.cycle_cnt[21] ),
    .C(_0474_),
    .Y(_0477_));
 sky130_fd_sc_hd__and3_1 _0633_ (.A(_0436_),
    .B(_0476_),
    .C(_0477_),
    .X(_0026_));
 sky130_fd_sc_hd__nand2_1 _0634_ (.A(\systolic_inst.cycle_cnt[22] ),
    .B(_0436_),
    .Y(_0478_));
 sky130_fd_sc_hd__and3_1 _0635_ (.A(\systolic_inst.cycle_cnt[20] ),
    .B(\systolic_inst.cycle_cnt[21] ),
    .C(\systolic_inst.cycle_cnt[22] ),
    .X(_0479_));
 sky130_fd_sc_hd__nand2_1 _0636_ (.A(_0474_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a21boi_1 _0637_ (.A1(_0477_),
    .A2(_0478_),
    .B1_N(_0480_),
    .Y(_0027_));
 sky130_fd_sc_hd__nor2_1 _0638_ (.A(_0399_),
    .B(_0435_),
    .Y(_0481_));
 sky130_fd_sc_hd__mux2_1 _0639_ (.A0(_0399_),
    .A1(_0481_),
    .S(_0480_),
    .X(_0028_));
 sky130_fd_sc_hd__and3_1 _0640_ (.A(\systolic_inst.cycle_cnt[23] ),
    .B(_0473_),
    .C(_0479_),
    .X(_0482_));
 sky130_fd_sc_hd__and4_1 _0641_ (.A(\systolic_inst.ce_local ),
    .B(_0447_),
    .C(_0464_),
    .D(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__o21ai_1 _0642_ (.A1(\systolic_inst.cycle_cnt[24] ),
    .A2(_0483_),
    .B1(_0436_),
    .Y(_0484_));
 sky130_fd_sc_hd__a21oi_1 _0643_ (.A1(\systolic_inst.cycle_cnt[24] ),
    .A2(_0483_),
    .B1(_0484_),
    .Y(_0029_));
 sky130_fd_sc_hd__a31o_1 _0644_ (.A1(\systolic_inst.cycle_cnt[24] ),
    .A2(_0470_),
    .A3(_0482_),
    .B1(\systolic_inst.cycle_cnt[25] ),
    .X(_0485_));
 sky130_fd_sc_hd__and2_1 _0645_ (.A(\systolic_inst.cycle_cnt[24] ),
    .B(\systolic_inst.cycle_cnt[25] ),
    .X(_0486_));
 sky130_fd_sc_hd__nand2_1 _0646_ (.A(_0483_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__and3_1 _0647_ (.A(_0436_),
    .B(_0485_),
    .C(_0487_),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_1 _0648_ (.A(\systolic_inst.cycle_cnt[26] ),
    .B(_0436_),
    .Y(_0488_));
 sky130_fd_sc_hd__and3_1 _0649_ (.A(\systolic_inst.cycle_cnt[26] ),
    .B(_0483_),
    .C(_0486_),
    .X(_0489_));
 sky130_fd_sc_hd__a21oi_1 _0650_ (.A1(_0487_),
    .A2(_0488_),
    .B1(_0489_),
    .Y(_0031_));
 sky130_fd_sc_hd__and2_1 _0651_ (.A(\systolic_inst.cycle_cnt[27] ),
    .B(_0436_),
    .X(_0490_));
 sky130_fd_sc_hd__and3_1 _0652_ (.A(\systolic_inst.cycle_cnt[26] ),
    .B(\systolic_inst.cycle_cnt[27] ),
    .C(_0486_),
    .X(_0491_));
 sky130_fd_sc_hd__and4_1 _0653_ (.A(_0448_),
    .B(_0464_),
    .C(_0482_),
    .D(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__o21ba_1 _0654_ (.A1(_0489_),
    .A2(_0490_),
    .B1_N(_0492_),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _0655_ (.A(\systolic_inst.cycle_cnt[28] ),
    .B(_0436_),
    .X(_0493_));
 sky130_fd_sc_hd__nand2_1 _0656_ (.A(\systolic_inst.cycle_cnt[28] ),
    .B(_0492_),
    .Y(_0494_));
 sky130_fd_sc_hd__o21a_1 _0657_ (.A1(_0492_),
    .A2(_0493_),
    .B1(_0494_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _0658_ (.A(\systolic_inst.cycle_cnt[29] ),
    .B(_0436_),
    .Y(_0495_));
 sky130_fd_sc_hd__and3_1 _0659_ (.A(\systolic_inst.cycle_cnt[28] ),
    .B(\systolic_inst.cycle_cnt[29] ),
    .C(_0492_),
    .X(_0496_));
 sky130_fd_sc_hd__a21oi_1 _0660_ (.A1(_0494_),
    .A2(_0495_),
    .B1(_0496_),
    .Y(_0034_));
 sky130_fd_sc_hd__nor2_1 _0661_ (.A(_0400_),
    .B(_0435_),
    .Y(_0497_));
 sky130_fd_sc_hd__and4_1 _0662_ (.A(\systolic_inst.cycle_cnt[28] ),
    .B(\systolic_inst.cycle_cnt[29] ),
    .C(\systolic_inst.cycle_cnt[30] ),
    .D(_0492_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _0663_ (.A0(_0497_),
    .A1(_0400_),
    .S(_0496_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_1 _0664_ (.A(_0401_),
    .B(_0435_),
    .Y(_0499_));
 sky130_fd_sc_hd__mux2_1 _0665_ (.A0(_0499_),
    .A1(_0401_),
    .S(_0498_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0666_ (.A0(\deser_A.receiving ),
    .A1(_0419_),
    .S(\deser_A.bit_idx[0] ),
    .X(_0037_));
 sky130_fd_sc_hd__and2b_1 _0667_ (.A_N(\deser_A.receiving ),
    .B(net1),
    .X(_0500_));
 sky130_fd_sc_hd__nand2b_4 _0668_ (.A_N(\deser_A.receiving ),
    .B(net1),
    .Y(_0501_));
 sky130_fd_sc_hd__and3_1 _0669_ (.A(\deser_A.receiving ),
    .B(\deser_A.bit_idx[1] ),
    .C(\deser_A.bit_idx[0] ),
    .X(_0502_));
 sky130_fd_sc_hd__nor2_1 _0670_ (.A(_0500_),
    .B(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__a21o_1 _0671_ (.A1(\deser_A.bit_idx[0] ),
    .A2(_0420_),
    .B1(\deser_A.bit_idx[1] ),
    .X(_0504_));
 sky130_fd_sc_hd__and2_1 _0672_ (.A(_0503_),
    .B(_0504_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0673_ (.A0(_0502_),
    .A1(_0503_),
    .S(\deser_A.bit_idx[2] ),
    .X(_0039_));
 sky130_fd_sc_hd__a41o_1 _0674_ (.A1(\deser_A.bit_idx[1] ),
    .A2(\deser_A.bit_idx[0] ),
    .A3(\deser_A.bit_idx[2] ),
    .A4(_0420_),
    .B1(\deser_A.bit_idx[3] ),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_1 _0675_ (.A(\deser_A.receiving ),
    .B(_0415_),
    .Y(_0506_));
 sky130_fd_sc_hd__and3_1 _0676_ (.A(_0501_),
    .B(_0505_),
    .C(_0506_),
    .X(_0040_));
 sky130_fd_sc_hd__nand2_1 _0677_ (.A(\deser_A.bit_idx[4] ),
    .B(_0501_),
    .Y(_0507_));
 sky130_fd_sc_hd__mux2_1 _0678_ (.A0(\deser_A.bit_idx[4] ),
    .A1(_0507_),
    .S(_0506_),
    .X(_0508_));
 sky130_fd_sc_hd__inv_2 _0679_ (.A(_0508_),
    .Y(_0041_));
 sky130_fd_sc_hd__nand3_1 _0680_ (.A(\deser_A.bit_idx[5] ),
    .B(_0416_),
    .C(_0420_),
    .Y(_0509_));
 sky130_fd_sc_hd__a31o_1 _0681_ (.A1(\deser_A.bit_idx[4] ),
    .A2(_0415_),
    .A3(_0420_),
    .B1(\deser_A.bit_idx[5] ),
    .X(_0510_));
 sky130_fd_sc_hd__and3_1 _0682_ (.A(_0501_),
    .B(_0509_),
    .C(_0510_),
    .X(_0042_));
 sky130_fd_sc_hd__a31o_1 _0683_ (.A1(\deser_A.bit_idx[5] ),
    .A2(_0416_),
    .A3(_0420_),
    .B1(\deser_A.bit_idx[6] ),
    .X(_0511_));
 sky130_fd_sc_hd__and3_1 _0684_ (.A(_0417_),
    .B(_0501_),
    .C(_0511_),
    .X(_0043_));
 sky130_fd_sc_hd__and3_1 _0685_ (.A(\deser_A.bit_idx[7] ),
    .B(_0417_),
    .C(_0501_),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _0686_ (.A(_0418_),
    .B(_0512_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(\deser_A.receiving ),
    .A1(_0419_),
    .S(\deser_A.kept_bit_idx[0] ),
    .X(_0045_));
 sky130_fd_sc_hd__a21oi_1 _0688_ (.A1(\deser_A.kept_bit_idx[0] ),
    .A2(_0420_),
    .B1(\deser_A.kept_bit_idx[1] ),
    .Y(_0513_));
 sky130_fd_sc_hd__and3_1 _0689_ (.A(net13),
    .B(\deser_A.kept_bit_idx[0] ),
    .C(\deser_A.kept_bit_idx[1] ),
    .X(_0514_));
 sky130_fd_sc_hd__nor3_1 _0690_ (.A(_0500_),
    .B(_0513_),
    .C(_0514_),
    .Y(_0046_));
 sky130_fd_sc_hd__and3_1 _0691_ (.A(\deser_A.kept_bit_idx[0] ),
    .B(\deser_A.kept_bit_idx[1] ),
    .C(\deser_A.kept_bit_idx[2] ),
    .X(_0515_));
 sky130_fd_sc_hd__and4_1 _0692_ (.A(net13),
    .B(\deser_A.kept_bit_idx[0] ),
    .C(\deser_A.kept_bit_idx[1] ),
    .D(\deser_A.kept_bit_idx[2] ),
    .X(_0516_));
 sky130_fd_sc_hd__a21oi_1 _0693_ (.A1(\deser_A.kept_bit_idx[2] ),
    .A2(_0501_),
    .B1(_0514_),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2_1 _0694_ (.A(_0516_),
    .B(_0517_),
    .Y(_0047_));
 sky130_fd_sc_hd__a21oi_1 _0695_ (.A1(\deser_A.kept_bit_idx[3] ),
    .A2(_0501_),
    .B1(_0516_),
    .Y(_0518_));
 sky130_fd_sc_hd__a21oi_1 _0696_ (.A1(\deser_A.kept_bit_idx[3] ),
    .A2(_0516_),
    .B1(_0518_),
    .Y(_0048_));
 sky130_fd_sc_hd__a22oi_1 _0697_ (.A1(\deser_A.kept_bit_idx[4] ),
    .A2(_0501_),
    .B1(_0516_),
    .B2(\deser_A.kept_bit_idx[3] ),
    .Y(_0519_));
 sky130_fd_sc_hd__a31o_1 _0698_ (.A1(\deser_A.kept_bit_idx[3] ),
    .A2(\deser_A.kept_bit_idx[4] ),
    .A3(_0516_),
    .B1(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(_0520_),
    .Y(_0049_));
 sky130_fd_sc_hd__and4_1 _0700_ (.A(\deser_A.kept_bit_idx[3] ),
    .B(\deser_A.kept_bit_idx[4] ),
    .C(\deser_A.kept_bit_idx[5] ),
    .D(_0516_),
    .X(_0521_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__a41o_1 _0702_ (.A1(\deser_A.kept_bit_idx[3] ),
    .A2(\deser_A.kept_bit_idx[4] ),
    .A3(_0420_),
    .A4(_0515_),
    .B1(\deser_A.kept_bit_idx[5] ),
    .X(_0523_));
 sky130_fd_sc_hd__and3_1 _0703_ (.A(_0501_),
    .B(_0522_),
    .C(_0523_),
    .X(_0050_));
 sky130_fd_sc_hd__nand2_1 _0704_ (.A(\deser_A.kept_bit_idx[6] ),
    .B(_0521_),
    .Y(_0524_));
 sky130_fd_sc_hd__a21o_1 _0705_ (.A1(\deser_A.kept_bit_idx[6] ),
    .A2(_0501_),
    .B1(_0521_),
    .X(_0525_));
 sky130_fd_sc_hd__and2_1 _0706_ (.A(_0524_),
    .B(_0525_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_1 _0707_ (.A(\deser_A.kept_bit_idx[7] ),
    .B(_0501_),
    .Y(_0526_));
 sky130_fd_sc_hd__mux2_1 _0708_ (.A0(\deser_A.kept_bit_idx[7] ),
    .A1(_0526_),
    .S(_0524_),
    .X(_0527_));
 sky130_fd_sc_hd__inv_2 _0709_ (.A(_0527_),
    .Y(_0052_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(\deser_A.kept_shift_reg[1] ),
    .A1(\deser_A.kept_shift_reg[2] ),
    .S(\deser_A.receiving ),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0711_ (.A0(\deser_A.kept_shift_reg[2] ),
    .A1(\deser_A.kept_shift_reg[3] ),
    .S(\deser_A.receiving ),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0712_ (.A0(\deser_A.kept_shift_reg[3] ),
    .A1(\deser_A.kept_shift_reg[4] ),
    .S(\deser_A.receiving ),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(\deser_A.kept_shift_reg[4] ),
    .A1(\deser_A.kept_shift_reg[5] ),
    .S(\deser_A.receiving ),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0714_ (.A0(\deser_A.kept_shift_reg[5] ),
    .A1(\deser_A.kept_shift_reg[6] ),
    .S(\deser_A.receiving ),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0715_ (.A0(\deser_A.kept_shift_reg[6] ),
    .A1(\deser_A.kept_shift_reg[7] ),
    .S(\deser_A.receiving ),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0716_ (.A0(\deser_A.kept_shift_reg[7] ),
    .A1(\deser_A.kept_shift_reg[8] ),
    .S(\deser_A.receiving ),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0717_ (.A0(\deser_A.kept_shift_reg[8] ),
    .A1(\deser_A.kept_shift_reg[9] ),
    .S(\deser_A.receiving ),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0718_ (.A0(\deser_A.kept_shift_reg[9] ),
    .A1(\deser_A.kept_shift_reg[10] ),
    .S(\deser_A.receiving ),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0719_ (.A0(\deser_A.kept_shift_reg[10] ),
    .A1(\deser_A.kept_shift_reg[11] ),
    .S(net13),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0720_ (.A0(\deser_A.kept_shift_reg[11] ),
    .A1(\deser_A.kept_shift_reg[12] ),
    .S(net13),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0721_ (.A0(\deser_A.kept_shift_reg[12] ),
    .A1(\deser_A.kept_shift_reg[13] ),
    .S(net13),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0722_ (.A0(\deser_A.kept_shift_reg[13] ),
    .A1(\deser_A.kept_shift_reg[14] ),
    .S(net13),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(\deser_A.kept_shift_reg[14] ),
    .A1(\deser_A.kept_shift_reg[15] ),
    .S(net13),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0724_ (.A0(\deser_A.kept_shift_reg[15] ),
    .A1(\deser_A.kept_shift_reg[16] ),
    .S(net13),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0725_ (.A0(\deser_A.kept_shift_reg[16] ),
    .A1(\deser_A.kept_shift_reg[17] ),
    .S(net13),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(\deser_A.kept_shift_reg[17] ),
    .A1(\deser_A.kept_shift_reg[18] ),
    .S(net13),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0727_ (.A0(\deser_A.kept_shift_reg[18] ),
    .A1(\deser_A.kept_shift_reg[19] ),
    .S(net13),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0728_ (.A0(\deser_A.kept_shift_reg[19] ),
    .A1(\deser_A.kept_shift_reg[20] ),
    .S(net13),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0729_ (.A0(\deser_A.kept_shift_reg[20] ),
    .A1(\deser_A.kept_shift_reg[21] ),
    .S(net13),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _0730_ (.A0(\deser_A.kept_shift_reg[21] ),
    .A1(\deser_A.kept_shift_reg[22] ),
    .S(net13),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0731_ (.A0(\deser_A.kept_shift_reg[22] ),
    .A1(\deser_A.kept_shift_reg[23] ),
    .S(net13),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(\deser_A.kept_shift_reg[23] ),
    .A1(\deser_A.kept_shift_reg[24] ),
    .S(net13),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0733_ (.A0(\deser_A.kept_shift_reg[24] ),
    .A1(\deser_A.kept_shift_reg[25] ),
    .S(net13),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _0734_ (.A0(\deser_A.kept_shift_reg[25] ),
    .A1(\deser_A.kept_shift_reg[26] ),
    .S(net13),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(\deser_A.kept_shift_reg[26] ),
    .A1(\deser_A.kept_shift_reg[27] ),
    .S(net13),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(\deser_A.kept_shift_reg[27] ),
    .A1(\deser_A.kept_shift_reg[28] ),
    .S(\deser_A.receiving ),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0737_ (.A0(\deser_A.kept_shift_reg[28] ),
    .A1(\deser_A.kept_shift_reg[29] ),
    .S(\deser_A.receiving ),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0738_ (.A0(\deser_A.kept_shift_reg[29] ),
    .A1(\deser_A.kept_shift_reg[30] ),
    .S(\deser_A.receiving ),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0739_ (.A0(\deser_A.kept_shift_reg[30] ),
    .A1(\deser_A.kept_shift_reg[31] ),
    .S(\deser_A.receiving ),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(\deser_A.kept_shift_reg[31] ),
    .A1(\deser_A.kept_shift_reg[32] ),
    .S(\deser_A.receiving ),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0741_ (.A0(\deser_A.kept_shift_reg[32] ),
    .A1(\deser_A.kept_shift_reg[33] ),
    .S(net12),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(\deser_A.kept_shift_reg[33] ),
    .A1(\deser_A.kept_shift_reg[34] ),
    .S(net12),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0743_ (.A0(\deser_A.kept_shift_reg[34] ),
    .A1(\deser_A.kept_shift_reg[35] ),
    .S(net12),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0744_ (.A0(\deser_A.kept_shift_reg[35] ),
    .A1(\deser_A.kept_shift_reg[36] ),
    .S(net12),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0745_ (.A0(\deser_A.kept_shift_reg[36] ),
    .A1(\deser_A.kept_shift_reg[37] ),
    .S(net12),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0746_ (.A0(\deser_A.kept_shift_reg[37] ),
    .A1(\deser_A.kept_shift_reg[38] ),
    .S(net12),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0747_ (.A0(\deser_A.kept_shift_reg[38] ),
    .A1(\deser_A.kept_shift_reg[39] ),
    .S(net12),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(\deser_A.kept_shift_reg[39] ),
    .A1(\deser_A.kept_shift_reg[40] ),
    .S(net12),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0749_ (.A0(\deser_A.kept_shift_reg[40] ),
    .A1(\deser_A.kept_shift_reg[41] ),
    .S(net12),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0750_ (.A0(\deser_A.kept_shift_reg[41] ),
    .A1(\deser_A.kept_shift_reg[42] ),
    .S(net12),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0751_ (.A0(\deser_A.kept_shift_reg[42] ),
    .A1(\deser_A.kept_shift_reg[43] ),
    .S(net12),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(\deser_A.kept_shift_reg[43] ),
    .A1(\deser_A.kept_shift_reg[44] ),
    .S(net12),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0753_ (.A0(\deser_A.kept_shift_reg[44] ),
    .A1(\deser_A.kept_shift_reg[45] ),
    .S(net12),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0754_ (.A0(\deser_A.kept_shift_reg[45] ),
    .A1(\deser_A.kept_shift_reg[46] ),
    .S(net12),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0755_ (.A0(\deser_A.kept_shift_reg[46] ),
    .A1(\deser_A.kept_shift_reg[47] ),
    .S(net12),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(\deser_A.kept_shift_reg[47] ),
    .A1(\deser_A.kept_shift_reg[48] ),
    .S(net13),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0757_ (.A0(\deser_A.kept_shift_reg[48] ),
    .A1(\deser_A.kept_shift_reg[49] ),
    .S(net13),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(\deser_A.kept_shift_reg[49] ),
    .A1(\deser_A.kept_shift_reg[50] ),
    .S(net13),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0759_ (.A0(\deser_A.kept_shift_reg[50] ),
    .A1(\deser_A.kept_shift_reg[51] ),
    .S(net13),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(\deser_A.kept_shift_reg[51] ),
    .A1(\deser_A.kept_shift_reg[52] ),
    .S(net13),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0761_ (.A0(\deser_A.kept_shift_reg[52] ),
    .A1(\deser_A.kept_shift_reg[53] ),
    .S(net13),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0762_ (.A0(\deser_A.kept_shift_reg[53] ),
    .A1(\deser_A.kept_shift_reg[54] ),
    .S(net13),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0763_ (.A0(\deser_A.kept_shift_reg[54] ),
    .A1(\deser_A.kept_shift_reg[55] ),
    .S(net13),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(\deser_A.kept_shift_reg[55] ),
    .A1(\deser_A.kept_shift_reg[56] ),
    .S(net13),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(\deser_A.kept_shift_reg[56] ),
    .A1(\deser_A.kept_shift_reg[57] ),
    .S(net13),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0766_ (.A0(\deser_A.kept_shift_reg[57] ),
    .A1(\deser_A.kept_shift_reg[58] ),
    .S(net13),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(\deser_A.kept_shift_reg[58] ),
    .A1(\deser_A.kept_shift_reg[59] ),
    .S(net13),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0768_ (.A0(\deser_A.kept_shift_reg[59] ),
    .A1(\deser_A.kept_shift_reg[60] ),
    .S(net13),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0769_ (.A0(\deser_A.kept_shift_reg[60] ),
    .A1(\deser_A.kept_shift_reg[61] ),
    .S(net13),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0770_ (.A0(\deser_A.kept_shift_reg[61] ),
    .A1(\deser_A.kept_shift_reg[62] ),
    .S(net13),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(\deser_A.kept_shift_reg[62] ),
    .A1(\deser_A.kept_shift_reg[63] ),
    .S(net13),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(\deser_A.kept_shift_reg[63] ),
    .A1(\deser_A.kept_shift_reg[64] ),
    .S(net13),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(\deser_A.kept_shift_reg[64] ),
    .A1(\deser_A.kept_shift_reg[65] ),
    .S(net13),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0774_ (.A0(\deser_A.kept_shift_reg[65] ),
    .A1(\deser_A.kept_shift_reg[66] ),
    .S(net13),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _0775_ (.A0(\deser_A.kept_shift_reg[66] ),
    .A1(\deser_A.kept_shift_reg[67] ),
    .S(net13),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0776_ (.A0(\deser_A.kept_shift_reg[67] ),
    .A1(\deser_A.kept_shift_reg[68] ),
    .S(net13),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(\deser_A.kept_shift_reg[68] ),
    .A1(\deser_A.kept_shift_reg[69] ),
    .S(net13),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0778_ (.A0(\deser_A.kept_shift_reg[69] ),
    .A1(\deser_A.kept_shift_reg[70] ),
    .S(net13),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(\deser_A.kept_shift_reg[70] ),
    .A1(\deser_A.kept_shift_reg[71] ),
    .S(net13),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _0780_ (.A0(\deser_A.kept_shift_reg[71] ),
    .A1(\deser_A.kept_shift_reg[72] ),
    .S(net13),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0781_ (.A0(\deser_A.kept_shift_reg[72] ),
    .A1(\deser_A.kept_shift_reg[73] ),
    .S(net13),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _0782_ (.A0(\deser_A.kept_shift_reg[73] ),
    .A1(\deser_A.kept_shift_reg[74] ),
    .S(net13),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(\deser_A.kept_shift_reg[74] ),
    .A1(\deser_A.kept_shift_reg[75] ),
    .S(net13),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _0784_ (.A0(\deser_A.kept_shift_reg[75] ),
    .A1(\deser_A.kept_shift_reg[76] ),
    .S(net13),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(\deser_A.kept_shift_reg[76] ),
    .A1(\deser_A.kept_shift_reg[77] ),
    .S(net13),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0786_ (.A0(\deser_A.kept_shift_reg[77] ),
    .A1(\deser_A.kept_shift_reg[78] ),
    .S(net13),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(\deser_A.kept_shift_reg[78] ),
    .A1(\deser_A.kept_shift_reg[79] ),
    .S(net13),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _0788_ (.A0(\deser_A.kept_shift_reg[79] ),
    .A1(\deser_A.kept_shift_reg[80] ),
    .S(net12),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(\deser_A.kept_shift_reg[80] ),
    .A1(\deser_A.kept_shift_reg[81] ),
    .S(net12),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _0790_ (.A0(\deser_A.kept_shift_reg[81] ),
    .A1(\deser_A.kept_shift_reg[82] ),
    .S(net12),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(\deser_A.kept_shift_reg[82] ),
    .A1(\deser_A.kept_shift_reg[83] ),
    .S(net12),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _0792_ (.A0(\deser_A.kept_shift_reg[83] ),
    .A1(\deser_A.kept_shift_reg[84] ),
    .S(net12),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(\deser_A.kept_shift_reg[84] ),
    .A1(\deser_A.kept_shift_reg[85] ),
    .S(net12),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _0794_ (.A0(\deser_A.kept_shift_reg[85] ),
    .A1(\deser_A.kept_shift_reg[86] ),
    .S(net12),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0795_ (.A0(\deser_A.kept_shift_reg[86] ),
    .A1(\deser_A.kept_shift_reg[87] ),
    .S(net12),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _0796_ (.A0(\deser_A.kept_shift_reg[87] ),
    .A1(\deser_A.kept_shift_reg[88] ),
    .S(net12),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0797_ (.A0(\deser_A.kept_shift_reg[88] ),
    .A1(\deser_A.kept_shift_reg[89] ),
    .S(net12),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _0798_ (.A0(\deser_A.kept_shift_reg[89] ),
    .A1(\deser_A.kept_shift_reg[90] ),
    .S(net12),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _0799_ (.A0(\deser_A.kept_shift_reg[90] ),
    .A1(\deser_A.kept_shift_reg[91] ),
    .S(net12),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0800_ (.A0(\deser_A.kept_shift_reg[91] ),
    .A1(\deser_A.kept_shift_reg[92] ),
    .S(net12),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(\deser_A.kept_shift_reg[92] ),
    .A1(\deser_A.kept_shift_reg[93] ),
    .S(net12),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0802_ (.A0(\deser_A.kept_shift_reg[93] ),
    .A1(\deser_A.kept_shift_reg[94] ),
    .S(net12),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0803_ (.A0(\deser_A.kept_shift_reg[94] ),
    .A1(\deser_A.kept_shift_reg[95] ),
    .S(net12),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _0804_ (.A0(\deser_A.kept_shift_reg[95] ),
    .A1(\deser_A.kept_shift_reg[96] ),
    .S(net12),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(\deser_A.kept_shift_reg[96] ),
    .A1(\deser_A.kept_shift_reg[97] ),
    .S(net12),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0806_ (.A0(\deser_A.kept_shift_reg[97] ),
    .A1(\deser_A.kept_shift_reg[98] ),
    .S(net12),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0807_ (.A0(\deser_A.kept_shift_reg[98] ),
    .A1(\deser_A.kept_shift_reg[99] ),
    .S(net12),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0808_ (.A0(\deser_A.kept_shift_reg[99] ),
    .A1(\deser_A.kept_shift_reg[100] ),
    .S(net12),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(\deser_A.kept_shift_reg[100] ),
    .A1(\deser_A.kept_shift_reg[101] ),
    .S(net12),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0810_ (.A0(\deser_A.kept_shift_reg[101] ),
    .A1(\deser_A.kept_shift_reg[102] ),
    .S(net12),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0811_ (.A0(\deser_A.kept_shift_reg[102] ),
    .A1(\deser_A.kept_shift_reg[103] ),
    .S(net12),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _0812_ (.A0(\deser_A.kept_shift_reg[103] ),
    .A1(\deser_A.kept_shift_reg[104] ),
    .S(net12),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(\deser_A.kept_shift_reg[104] ),
    .A1(\deser_A.kept_shift_reg[105] ),
    .S(net12),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _0814_ (.A0(\deser_A.kept_shift_reg[105] ),
    .A1(\deser_A.kept_shift_reg[106] ),
    .S(net12),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _0815_ (.A0(\deser_A.kept_shift_reg[106] ),
    .A1(\deser_A.kept_shift_reg[107] ),
    .S(net12),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _0816_ (.A0(\deser_A.kept_shift_reg[107] ),
    .A1(\deser_A.kept_shift_reg[108] ),
    .S(net12),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _0817_ (.A0(\deser_A.kept_shift_reg[108] ),
    .A1(\deser_A.kept_shift_reg[109] ),
    .S(net12),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _0818_ (.A0(\deser_A.kept_shift_reg[109] ),
    .A1(\deser_A.kept_shift_reg[110] ),
    .S(net12),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _0819_ (.A0(\deser_A.kept_shift_reg[110] ),
    .A1(\deser_A.kept_shift_reg[111] ),
    .S(net12),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _0820_ (.A0(\deser_A.kept_shift_reg[111] ),
    .A1(\deser_A.kept_shift_reg[112] ),
    .S(net12),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _0821_ (.A0(\deser_A.kept_shift_reg[112] ),
    .A1(\deser_A.kept_shift_reg[113] ),
    .S(net12),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _0822_ (.A0(\deser_A.kept_shift_reg[113] ),
    .A1(\deser_A.kept_shift_reg[114] ),
    .S(net12),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _0823_ (.A0(\deser_A.kept_shift_reg[114] ),
    .A1(\deser_A.kept_shift_reg[115] ),
    .S(net12),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _0824_ (.A0(\deser_A.kept_shift_reg[115] ),
    .A1(\deser_A.kept_shift_reg[116] ),
    .S(net12),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _0825_ (.A0(\deser_A.kept_shift_reg[116] ),
    .A1(\deser_A.kept_shift_reg[117] ),
    .S(net12),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _0826_ (.A0(\deser_A.kept_shift_reg[117] ),
    .A1(\deser_A.kept_shift_reg[118] ),
    .S(net12),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _0827_ (.A0(\deser_A.kept_shift_reg[118] ),
    .A1(\deser_A.kept_shift_reg[119] ),
    .S(net12),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(\deser_A.kept_shift_reg[119] ),
    .A1(\deser_A.kept_shift_reg[120] ),
    .S(net12),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0829_ (.A0(\deser_A.kept_shift_reg[120] ),
    .A1(\deser_A.kept_shift_reg[121] ),
    .S(net12),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _0830_ (.A0(\deser_A.kept_shift_reg[121] ),
    .A1(\deser_A.kept_shift_reg[122] ),
    .S(net12),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _0831_ (.A0(\deser_A.kept_shift_reg[122] ),
    .A1(\deser_A.kept_shift_reg[123] ),
    .S(net12),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _0832_ (.A0(\deser_A.kept_shift_reg[123] ),
    .A1(\deser_A.kept_shift_reg[124] ),
    .S(net12),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _0833_ (.A0(\deser_A.kept_shift_reg[124] ),
    .A1(\deser_A.kept_shift_reg[125] ),
    .S(net12),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _0834_ (.A0(\deser_A.kept_shift_reg[125] ),
    .A1(\deser_A.kept_shift_reg[126] ),
    .S(net12),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _0835_ (.A0(\deser_A.kept_shift_reg[126] ),
    .A1(\deser_A.kept_shift_reg[127] ),
    .S(net12),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _0836_ (.A0(\deser_A.kept_shift_reg[127] ),
    .A1(net2),
    .S(net12),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _0837_ (.A0(\deser_B.receiving ),
    .A1(_0425_),
    .S(\deser_B.bit_idx[0] ),
    .X(_0180_));
 sky130_fd_sc_hd__and2b_1 _0838_ (.A_N(\deser_B.receiving ),
    .B(net3),
    .X(_0347_));
 sky130_fd_sc_hd__nand2b_4 _0839_ (.A_N(\deser_B.receiving ),
    .B(net3),
    .Y(_0348_));
 sky130_fd_sc_hd__and3_1 _0840_ (.A(\deser_B.receiving ),
    .B(\deser_B.bit_idx[1] ),
    .C(\deser_B.bit_idx[0] ),
    .X(_0349_));
 sky130_fd_sc_hd__nor2_1 _0841_ (.A(_0347_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__a21o_1 _0842_ (.A1(\deser_B.bit_idx[0] ),
    .A2(_0426_),
    .B1(\deser_B.bit_idx[1] ),
    .X(_0351_));
 sky130_fd_sc_hd__and2_1 _0843_ (.A(_0350_),
    .B(_0351_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(_0349_),
    .A1(_0350_),
    .S(\deser_B.bit_idx[2] ),
    .X(_0182_));
 sky130_fd_sc_hd__a41o_1 _0845_ (.A1(\deser_B.bit_idx[1] ),
    .A2(\deser_B.bit_idx[0] ),
    .A3(\deser_B.bit_idx[2] ),
    .A4(_0426_),
    .B1(\deser_B.bit_idx[3] ),
    .X(_0352_));
 sky130_fd_sc_hd__nand2_1 _0846_ (.A(\deser_B.receiving ),
    .B(_0421_),
    .Y(_0353_));
 sky130_fd_sc_hd__and3_1 _0847_ (.A(_0348_),
    .B(_0352_),
    .C(_0353_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_1 _0848_ (.A(\deser_B.bit_idx[4] ),
    .B(_0348_),
    .Y(_0354_));
 sky130_fd_sc_hd__mux2_1 _0849_ (.A0(\deser_B.bit_idx[4] ),
    .A1(_0354_),
    .S(_0353_),
    .X(_0355_));
 sky130_fd_sc_hd__inv_2 _0850_ (.A(_0355_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21oi_1 _0851_ (.A1(_0422_),
    .A2(_0426_),
    .B1(\deser_B.bit_idx[5] ),
    .Y(_0356_));
 sky130_fd_sc_hd__a31o_1 _0852_ (.A1(\deser_B.bit_idx[5] ),
    .A2(_0422_),
    .A3(_0426_),
    .B1(_0347_),
    .X(_0357_));
 sky130_fd_sc_hd__nor2_1 _0853_ (.A(_0356_),
    .B(_0357_),
    .Y(_0185_));
 sky130_fd_sc_hd__a31o_1 _0854_ (.A1(\deser_B.bit_idx[5] ),
    .A2(_0422_),
    .A3(_0426_),
    .B1(\deser_B.bit_idx[6] ),
    .X(_0358_));
 sky130_fd_sc_hd__and3_1 _0855_ (.A(_0423_),
    .B(_0348_),
    .C(_0358_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _0856_ (.A(\deser_B.bit_idx[7] ),
    .B(_0423_),
    .C(_0348_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _0857_ (.A(_0424_),
    .B(_0359_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _0858_ (.A0(\deser_B.receiving ),
    .A1(_0425_),
    .S(\deser_B.kept_bit_idx[0] ),
    .X(_0188_));
 sky130_fd_sc_hd__a21oi_1 _0859_ (.A1(\deser_B.kept_bit_idx[0] ),
    .A2(_0426_),
    .B1(\deser_B.kept_bit_idx[1] ),
    .Y(_0360_));
 sky130_fd_sc_hd__and3_1 _0860_ (.A(\deser_B.receiving ),
    .B(\deser_B.kept_bit_idx[0] ),
    .C(\deser_B.kept_bit_idx[1] ),
    .X(_0361_));
 sky130_fd_sc_hd__nor3_1 _0861_ (.A(_0347_),
    .B(_0360_),
    .C(_0361_),
    .Y(_0189_));
 sky130_fd_sc_hd__and3_1 _0862_ (.A(\deser_B.kept_bit_idx[0] ),
    .B(\deser_B.kept_bit_idx[1] ),
    .C(\deser_B.kept_bit_idx[2] ),
    .X(_0362_));
 sky130_fd_sc_hd__and4_1 _0863_ (.A(\deser_B.receiving ),
    .B(\deser_B.kept_bit_idx[0] ),
    .C(\deser_B.kept_bit_idx[1] ),
    .D(\deser_B.kept_bit_idx[2] ),
    .X(_0363_));
 sky130_fd_sc_hd__a21oi_1 _0864_ (.A1(\deser_B.kept_bit_idx[2] ),
    .A2(_0348_),
    .B1(_0361_),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _0865_ (.A(_0363_),
    .B(_0364_),
    .Y(_0190_));
 sky130_fd_sc_hd__a21oi_1 _0866_ (.A1(\deser_B.kept_bit_idx[3] ),
    .A2(_0348_),
    .B1(_0363_),
    .Y(_0365_));
 sky130_fd_sc_hd__a21oi_1 _0867_ (.A1(\deser_B.kept_bit_idx[3] ),
    .A2(_0363_),
    .B1(_0365_),
    .Y(_0191_));
 sky130_fd_sc_hd__a22oi_1 _0868_ (.A1(\deser_B.kept_bit_idx[4] ),
    .A2(_0348_),
    .B1(_0363_),
    .B2(\deser_B.kept_bit_idx[3] ),
    .Y(_0366_));
 sky130_fd_sc_hd__a31o_1 _0869_ (.A1(\deser_B.kept_bit_idx[3] ),
    .A2(\deser_B.kept_bit_idx[4] ),
    .A3(_0363_),
    .B1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__inv_2 _0870_ (.A(_0367_),
    .Y(_0192_));
 sky130_fd_sc_hd__and4_1 _0871_ (.A(\deser_B.kept_bit_idx[3] ),
    .B(\deser_B.kept_bit_idx[4] ),
    .C(\deser_B.kept_bit_idx[5] ),
    .D(_0363_),
    .X(_0368_));
 sky130_fd_sc_hd__inv_2 _0872_ (.A(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__a41o_1 _0873_ (.A1(\deser_B.kept_bit_idx[3] ),
    .A2(\deser_B.kept_bit_idx[4] ),
    .A3(_0426_),
    .A4(_0362_),
    .B1(\deser_B.kept_bit_idx[5] ),
    .X(_0370_));
 sky130_fd_sc_hd__and3_1 _0874_ (.A(_0348_),
    .B(_0369_),
    .C(_0370_),
    .X(_0193_));
 sky130_fd_sc_hd__nand2_1 _0875_ (.A(\deser_B.kept_bit_idx[6] ),
    .B(_0368_),
    .Y(_0371_));
 sky130_fd_sc_hd__a21o_1 _0876_ (.A1(\deser_B.kept_bit_idx[6] ),
    .A2(_0348_),
    .B1(_0368_),
    .X(_0372_));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(_0371_),
    .B(_0372_),
    .X(_0194_));
 sky130_fd_sc_hd__nand2_1 _0878_ (.A(\deser_B.kept_bit_idx[7] ),
    .B(_0348_),
    .Y(_0373_));
 sky130_fd_sc_hd__mux2_1 _0879_ (.A0(\deser_B.kept_bit_idx[7] ),
    .A1(_0373_),
    .S(_0371_),
    .X(_0374_));
 sky130_fd_sc_hd__inv_2 _0880_ (.A(_0374_),
    .Y(_0195_));
 sky130_fd_sc_hd__o21ai_1 _0881_ (.A1(_0403_),
    .A2(_0418_),
    .B1(_0501_),
    .Y(_0196_));
 sky130_fd_sc_hd__mux2_1 _0882_ (.A0(\deser_B.kept_shift_reg[1] ),
    .A1(\deser_B.kept_shift_reg[2] ),
    .S(\deser_B.receiving ),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _0883_ (.A0(\deser_B.kept_shift_reg[2] ),
    .A1(\deser_B.kept_shift_reg[3] ),
    .S(\deser_B.receiving ),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _0884_ (.A0(\deser_B.kept_shift_reg[3] ),
    .A1(\deser_B.kept_shift_reg[4] ),
    .S(\deser_B.receiving ),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _0885_ (.A0(\deser_B.kept_shift_reg[4] ),
    .A1(\deser_B.kept_shift_reg[5] ),
    .S(net10),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _0886_ (.A0(\deser_B.kept_shift_reg[5] ),
    .A1(\deser_B.kept_shift_reg[6] ),
    .S(net10),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _0887_ (.A0(\deser_B.kept_shift_reg[6] ),
    .A1(\deser_B.kept_shift_reg[7] ),
    .S(net10),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(\deser_B.kept_shift_reg[7] ),
    .A1(\deser_B.kept_shift_reg[8] ),
    .S(net10),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _0889_ (.A0(\deser_B.kept_shift_reg[8] ),
    .A1(\deser_B.kept_shift_reg[9] ),
    .S(net10),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _0890_ (.A0(\deser_B.kept_shift_reg[9] ),
    .A1(\deser_B.kept_shift_reg[10] ),
    .S(net10),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _0891_ (.A0(\deser_B.kept_shift_reg[10] ),
    .A1(\deser_B.kept_shift_reg[11] ),
    .S(net11),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _0892_ (.A0(\deser_B.kept_shift_reg[11] ),
    .A1(\deser_B.kept_shift_reg[12] ),
    .S(net11),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _0893_ (.A0(\deser_B.kept_shift_reg[12] ),
    .A1(\deser_B.kept_shift_reg[13] ),
    .S(net11),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _0894_ (.A0(\deser_B.kept_shift_reg[13] ),
    .A1(\deser_B.kept_shift_reg[14] ),
    .S(net11),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _0895_ (.A0(\deser_B.kept_shift_reg[14] ),
    .A1(\deser_B.kept_shift_reg[15] ),
    .S(net11),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(\deser_B.kept_shift_reg[15] ),
    .A1(\deser_B.kept_shift_reg[16] ),
    .S(net11),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _0897_ (.A0(\deser_B.kept_shift_reg[16] ),
    .A1(\deser_B.kept_shift_reg[17] ),
    .S(net11),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(\deser_B.kept_shift_reg[17] ),
    .A1(\deser_B.kept_shift_reg[18] ),
    .S(net11),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _0899_ (.A0(\deser_B.kept_shift_reg[18] ),
    .A1(\deser_B.kept_shift_reg[19] ),
    .S(net11),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(\deser_B.kept_shift_reg[19] ),
    .A1(\deser_B.kept_shift_reg[20] ),
    .S(net11),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _0901_ (.A0(\deser_B.kept_shift_reg[20] ),
    .A1(\deser_B.kept_shift_reg[21] ),
    .S(net11),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _0902_ (.A0(\deser_B.kept_shift_reg[21] ),
    .A1(\deser_B.kept_shift_reg[22] ),
    .S(net11),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _0903_ (.A0(\deser_B.kept_shift_reg[22] ),
    .A1(\deser_B.kept_shift_reg[23] ),
    .S(net11),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(\deser_B.kept_shift_reg[23] ),
    .A1(\deser_B.kept_shift_reg[24] ),
    .S(net11),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _0905_ (.A0(\deser_B.kept_shift_reg[24] ),
    .A1(\deser_B.kept_shift_reg[25] ),
    .S(net11),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _0906_ (.A0(\deser_B.kept_shift_reg[25] ),
    .A1(\deser_B.kept_shift_reg[26] ),
    .S(net11),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _0907_ (.A0(\deser_B.kept_shift_reg[26] ),
    .A1(\deser_B.kept_shift_reg[27] ),
    .S(net11),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _0908_ (.A0(\deser_B.kept_shift_reg[27] ),
    .A1(\deser_B.kept_shift_reg[28] ),
    .S(net11),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _0909_ (.A0(\deser_B.kept_shift_reg[28] ),
    .A1(\deser_B.kept_shift_reg[29] ),
    .S(net11),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(\deser_B.kept_shift_reg[29] ),
    .A1(\deser_B.kept_shift_reg[30] ),
    .S(net11),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _0911_ (.A0(\deser_B.kept_shift_reg[30] ),
    .A1(\deser_B.kept_shift_reg[31] ),
    .S(net11),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(\deser_B.kept_shift_reg[31] ),
    .A1(\deser_B.kept_shift_reg[32] ),
    .S(net11),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _0913_ (.A0(\deser_B.kept_shift_reg[32] ),
    .A1(\deser_B.kept_shift_reg[33] ),
    .S(net11),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(\deser_B.kept_shift_reg[33] ),
    .A1(\deser_B.kept_shift_reg[34] ),
    .S(net11),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _0915_ (.A0(\deser_B.kept_shift_reg[34] ),
    .A1(\deser_B.kept_shift_reg[35] ),
    .S(net11),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(\deser_B.kept_shift_reg[35] ),
    .A1(\deser_B.kept_shift_reg[36] ),
    .S(net11),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _0917_ (.A0(\deser_B.kept_shift_reg[36] ),
    .A1(\deser_B.kept_shift_reg[37] ),
    .S(net11),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(\deser_B.kept_shift_reg[37] ),
    .A1(\deser_B.kept_shift_reg[38] ),
    .S(net11),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _0919_ (.A0(\deser_B.kept_shift_reg[38] ),
    .A1(\deser_B.kept_shift_reg[39] ),
    .S(net11),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(\deser_B.kept_shift_reg[39] ),
    .A1(\deser_B.kept_shift_reg[40] ),
    .S(net11),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _0921_ (.A0(\deser_B.kept_shift_reg[40] ),
    .A1(\deser_B.kept_shift_reg[41] ),
    .S(net11),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _0922_ (.A0(\deser_B.kept_shift_reg[41] ),
    .A1(\deser_B.kept_shift_reg[42] ),
    .S(net11),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0923_ (.A0(\deser_B.kept_shift_reg[42] ),
    .A1(\deser_B.kept_shift_reg[43] ),
    .S(net11),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _0924_ (.A0(\deser_B.kept_shift_reg[43] ),
    .A1(\deser_B.kept_shift_reg[44] ),
    .S(net11),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0925_ (.A0(\deser_B.kept_shift_reg[44] ),
    .A1(\deser_B.kept_shift_reg[45] ),
    .S(net11),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _0926_ (.A0(\deser_B.kept_shift_reg[45] ),
    .A1(\deser_B.kept_shift_reg[46] ),
    .S(net11),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _0927_ (.A0(\deser_B.kept_shift_reg[46] ),
    .A1(\deser_B.kept_shift_reg[47] ),
    .S(net11),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(\deser_B.kept_shift_reg[47] ),
    .A1(\deser_B.kept_shift_reg[48] ),
    .S(net11),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _0929_ (.A0(\deser_B.kept_shift_reg[48] ),
    .A1(\deser_B.kept_shift_reg[49] ),
    .S(net11),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0930_ (.A0(\deser_B.kept_shift_reg[49] ),
    .A1(\deser_B.kept_shift_reg[50] ),
    .S(net11),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _0931_ (.A0(\deser_B.kept_shift_reg[50] ),
    .A1(\deser_B.kept_shift_reg[51] ),
    .S(net11),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(\deser_B.kept_shift_reg[51] ),
    .A1(\deser_B.kept_shift_reg[52] ),
    .S(net11),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(\deser_B.kept_shift_reg[52] ),
    .A1(\deser_B.kept_shift_reg[53] ),
    .S(net11),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(\deser_B.kept_shift_reg[53] ),
    .A1(\deser_B.kept_shift_reg[54] ),
    .S(net11),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _0935_ (.A0(\deser_B.kept_shift_reg[54] ),
    .A1(\deser_B.kept_shift_reg[55] ),
    .S(net11),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(\deser_B.kept_shift_reg[55] ),
    .A1(\deser_B.kept_shift_reg[56] ),
    .S(net10),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0937_ (.A0(\deser_B.kept_shift_reg[56] ),
    .A1(\deser_B.kept_shift_reg[57] ),
    .S(net10),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(\deser_B.kept_shift_reg[57] ),
    .A1(\deser_B.kept_shift_reg[58] ),
    .S(net10),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0939_ (.A0(\deser_B.kept_shift_reg[58] ),
    .A1(\deser_B.kept_shift_reg[59] ),
    .S(net10),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(\deser_B.kept_shift_reg[59] ),
    .A1(\deser_B.kept_shift_reg[60] ),
    .S(net10),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0941_ (.A0(\deser_B.kept_shift_reg[60] ),
    .A1(\deser_B.kept_shift_reg[61] ),
    .S(net10),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(\deser_B.kept_shift_reg[61] ),
    .A1(\deser_B.kept_shift_reg[62] ),
    .S(net10),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _0943_ (.A0(\deser_B.kept_shift_reg[62] ),
    .A1(\deser_B.kept_shift_reg[63] ),
    .S(net10),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(\deser_B.kept_shift_reg[63] ),
    .A1(\deser_B.kept_shift_reg[64] ),
    .S(net10),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _0945_ (.A0(\deser_B.kept_shift_reg[64] ),
    .A1(\deser_B.kept_shift_reg[65] ),
    .S(net10),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(\deser_B.kept_shift_reg[65] ),
    .A1(\deser_B.kept_shift_reg[66] ),
    .S(net10),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _0947_ (.A0(\deser_B.kept_shift_reg[66] ),
    .A1(\deser_B.kept_shift_reg[67] ),
    .S(net10),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(\deser_B.kept_shift_reg[67] ),
    .A1(\deser_B.kept_shift_reg[68] ),
    .S(net10),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _0949_ (.A0(\deser_B.kept_shift_reg[68] ),
    .A1(\deser_B.kept_shift_reg[69] ),
    .S(net10),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(\deser_B.kept_shift_reg[69] ),
    .A1(\deser_B.kept_shift_reg[70] ),
    .S(net10),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _0951_ (.A0(\deser_B.kept_shift_reg[70] ),
    .A1(\deser_B.kept_shift_reg[71] ),
    .S(net10),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(\deser_B.kept_shift_reg[71] ),
    .A1(\deser_B.kept_shift_reg[72] ),
    .S(net10),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(\deser_B.kept_shift_reg[72] ),
    .A1(\deser_B.kept_shift_reg[73] ),
    .S(net10),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(\deser_B.kept_shift_reg[73] ),
    .A1(\deser_B.kept_shift_reg[74] ),
    .S(net10),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _0955_ (.A0(\deser_B.kept_shift_reg[74] ),
    .A1(\deser_B.kept_shift_reg[75] ),
    .S(net10),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(\deser_B.kept_shift_reg[75] ),
    .A1(\deser_B.kept_shift_reg[76] ),
    .S(net10),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _0957_ (.A0(\deser_B.kept_shift_reg[76] ),
    .A1(\deser_B.kept_shift_reg[77] ),
    .S(net10),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(\deser_B.kept_shift_reg[77] ),
    .A1(\deser_B.kept_shift_reg[78] ),
    .S(net10),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _0959_ (.A0(\deser_B.kept_shift_reg[78] ),
    .A1(\deser_B.kept_shift_reg[79] ),
    .S(net10),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(\deser_B.kept_shift_reg[79] ),
    .A1(\deser_B.kept_shift_reg[80] ),
    .S(net10),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(\deser_B.kept_shift_reg[80] ),
    .A1(\deser_B.kept_shift_reg[81] ),
    .S(net10),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _0962_ (.A0(\deser_B.kept_shift_reg[81] ),
    .A1(\deser_B.kept_shift_reg[82] ),
    .S(net10),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _0963_ (.A0(\deser_B.kept_shift_reg[82] ),
    .A1(\deser_B.kept_shift_reg[83] ),
    .S(net10),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(\deser_B.kept_shift_reg[83] ),
    .A1(\deser_B.kept_shift_reg[84] ),
    .S(net10),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _0965_ (.A0(\deser_B.kept_shift_reg[84] ),
    .A1(\deser_B.kept_shift_reg[85] ),
    .S(net10),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _0966_ (.A0(\deser_B.kept_shift_reg[85] ),
    .A1(\deser_B.kept_shift_reg[86] ),
    .S(net10),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _0967_ (.A0(\deser_B.kept_shift_reg[86] ),
    .A1(\deser_B.kept_shift_reg[87] ),
    .S(net10),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(\deser_B.kept_shift_reg[87] ),
    .A1(\deser_B.kept_shift_reg[88] ),
    .S(net10),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _0969_ (.A0(\deser_B.kept_shift_reg[88] ),
    .A1(\deser_B.kept_shift_reg[89] ),
    .S(net10),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _0970_ (.A0(\deser_B.kept_shift_reg[89] ),
    .A1(\deser_B.kept_shift_reg[90] ),
    .S(net10),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _0971_ (.A0(\deser_B.kept_shift_reg[90] ),
    .A1(\deser_B.kept_shift_reg[91] ),
    .S(\deser_B.receiving ),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _0972_ (.A0(\deser_B.kept_shift_reg[91] ),
    .A1(\deser_B.kept_shift_reg[92] ),
    .S(\deser_B.receiving ),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(\deser_B.kept_shift_reg[92] ),
    .A1(\deser_B.kept_shift_reg[93] ),
    .S(\deser_B.receiving ),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _0974_ (.A0(\deser_B.kept_shift_reg[93] ),
    .A1(\deser_B.kept_shift_reg[94] ),
    .S(net10),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _0975_ (.A0(\deser_B.kept_shift_reg[94] ),
    .A1(\deser_B.kept_shift_reg[95] ),
    .S(net10),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _0976_ (.A0(\deser_B.kept_shift_reg[95] ),
    .A1(\deser_B.kept_shift_reg[96] ),
    .S(net10),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _0977_ (.A0(\deser_B.kept_shift_reg[96] ),
    .A1(\deser_B.kept_shift_reg[97] ),
    .S(net10),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _0978_ (.A0(\deser_B.kept_shift_reg[97] ),
    .A1(\deser_B.kept_shift_reg[98] ),
    .S(net10),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _0979_ (.A0(\deser_B.kept_shift_reg[98] ),
    .A1(\deser_B.kept_shift_reg[99] ),
    .S(net10),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _0980_ (.A0(\deser_B.kept_shift_reg[99] ),
    .A1(\deser_B.kept_shift_reg[100] ),
    .S(net10),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _0981_ (.A0(\deser_B.kept_shift_reg[100] ),
    .A1(\deser_B.kept_shift_reg[101] ),
    .S(net10),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _0982_ (.A0(\deser_B.kept_shift_reg[101] ),
    .A1(\deser_B.kept_shift_reg[102] ),
    .S(net10),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _0983_ (.A0(\deser_B.kept_shift_reg[102] ),
    .A1(\deser_B.kept_shift_reg[103] ),
    .S(net10),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(\deser_B.kept_shift_reg[103] ),
    .A1(\deser_B.kept_shift_reg[104] ),
    .S(net10),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _0985_ (.A0(\deser_B.kept_shift_reg[104] ),
    .A1(\deser_B.kept_shift_reg[105] ),
    .S(\deser_B.receiving ),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(\deser_B.kept_shift_reg[105] ),
    .A1(\deser_B.kept_shift_reg[106] ),
    .S(\deser_B.receiving ),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _0987_ (.A0(\deser_B.kept_shift_reg[106] ),
    .A1(\deser_B.kept_shift_reg[107] ),
    .S(\deser_B.receiving ),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _0988_ (.A0(\deser_B.kept_shift_reg[107] ),
    .A1(\deser_B.kept_shift_reg[108] ),
    .S(\deser_B.receiving ),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _0989_ (.A0(\deser_B.kept_shift_reg[108] ),
    .A1(\deser_B.kept_shift_reg[109] ),
    .S(\deser_B.receiving ),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(\deser_B.kept_shift_reg[109] ),
    .A1(\deser_B.kept_shift_reg[110] ),
    .S(\deser_B.receiving ),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(\deser_B.kept_shift_reg[110] ),
    .A1(\deser_B.kept_shift_reg[111] ),
    .S(\deser_B.receiving ),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _0992_ (.A0(\deser_B.kept_shift_reg[111] ),
    .A1(\deser_B.kept_shift_reg[112] ),
    .S(\deser_B.receiving ),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(\deser_B.kept_shift_reg[112] ),
    .A1(\deser_B.kept_shift_reg[113] ),
    .S(\deser_B.receiving ),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(\deser_B.kept_shift_reg[113] ),
    .A1(\deser_B.kept_shift_reg[114] ),
    .S(\deser_B.receiving ),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _0995_ (.A0(\deser_B.kept_shift_reg[114] ),
    .A1(\deser_B.kept_shift_reg[115] ),
    .S(\deser_B.receiving ),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(\deser_B.kept_shift_reg[115] ),
    .A1(\deser_B.kept_shift_reg[116] ),
    .S(\deser_B.receiving ),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(\deser_B.kept_shift_reg[116] ),
    .A1(\deser_B.kept_shift_reg[117] ),
    .S(\deser_B.receiving ),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _0998_ (.A0(\deser_B.kept_shift_reg[117] ),
    .A1(\deser_B.kept_shift_reg[118] ),
    .S(\deser_B.receiving ),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(\deser_B.kept_shift_reg[118] ),
    .A1(\deser_B.kept_shift_reg[119] ),
    .S(\deser_B.receiving ),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(\deser_B.kept_shift_reg[119] ),
    .A1(\deser_B.kept_shift_reg[120] ),
    .S(\deser_B.receiving ),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(\deser_B.kept_shift_reg[120] ),
    .A1(\deser_B.kept_shift_reg[121] ),
    .S(\deser_B.receiving ),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(\deser_B.kept_shift_reg[121] ),
    .A1(\deser_B.kept_shift_reg[122] ),
    .S(\deser_B.receiving ),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(\deser_B.kept_shift_reg[122] ),
    .A1(\deser_B.kept_shift_reg[123] ),
    .S(\deser_B.receiving ),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(\deser_B.kept_shift_reg[123] ),
    .A1(\deser_B.kept_shift_reg[124] ),
    .S(\deser_B.receiving ),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(\deser_B.kept_shift_reg[124] ),
    .A1(\deser_B.kept_shift_reg[125] ),
    .S(\deser_B.receiving ),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(\deser_B.kept_shift_reg[125] ),
    .A1(\deser_B.kept_shift_reg[126] ),
    .S(\deser_B.receiving ),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _1007_ (.A0(\deser_B.kept_shift_reg[126] ),
    .A1(\deser_B.kept_shift_reg[127] ),
    .S(\deser_B.receiving ),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(\deser_B.kept_shift_reg[127] ),
    .A1(net4),
    .S(\deser_B.receiving ),
    .X(_0323_));
 sky130_fd_sc_hd__and2_1 _1009_ (.A(\deser_B.receiving ),
    .B(\deser_B.kept_shift_reg[1] ),
    .X(_0375_));
 sky130_fd_sc_hd__a221o_1 _1010_ (.A1(\deser_B.kept_shift_reg[0] ),
    .A2(_0425_),
    .B1(_0347_),
    .B2(net4),
    .C1(_0375_),
    .X(_0324_));
 sky130_fd_sc_hd__and2_1 _1011_ (.A(\deser_A.receiving ),
    .B(\deser_A.kept_shift_reg[1] ),
    .X(_0376_));
 sky130_fd_sc_hd__a221o_1 _1012_ (.A1(\deser_A.kept_shift_reg[0] ),
    .A2(_0419_),
    .B1(_0500_),
    .B2(net2),
    .C1(_0376_),
    .X(_0325_));
 sky130_fd_sc_hd__xor2_1 _1013_ (.A(\ser_C.bit_idx[0] ),
    .B(net7),
    .X(_0326_));
 sky130_fd_sc_hd__and3_1 _1014_ (.A(\ser_C.bit_idx[0] ),
    .B(\ser_C.bit_idx[1] ),
    .C(net7),
    .X(_0377_));
 sky130_fd_sc_hd__a21oi_1 _1015_ (.A1(\ser_C.bit_idx[0] ),
    .A2(net7),
    .B1(\ser_C.bit_idx[1] ),
    .Y(_0378_));
 sky130_fd_sc_hd__nor2_1 _1016_ (.A(_0377_),
    .B(_0378_),
    .Y(_0327_));
 sky130_fd_sc_hd__and4_1 _1017_ (.A(\ser_C.bit_idx[0] ),
    .B(\ser_C.bit_idx[1] ),
    .C(\ser_C.bit_idx[2] ),
    .D(net7),
    .X(_0379_));
 sky130_fd_sc_hd__nor2_1 _1018_ (.A(\ser_C.bit_idx[2] ),
    .B(_0377_),
    .Y(_0380_));
 sky130_fd_sc_hd__nor2_1 _1019_ (.A(_0379_),
    .B(_0380_),
    .Y(_0328_));
 sky130_fd_sc_hd__xor2_1 _1020_ (.A(\ser_C.bit_idx[3] ),
    .B(_0379_),
    .X(_0329_));
 sky130_fd_sc_hd__and3_1 _1021_ (.A(\ser_C.bit_idx[3] ),
    .B(\ser_C.bit_idx[4] ),
    .C(_0379_),
    .X(_0381_));
 sky130_fd_sc_hd__a21oi_1 _1022_ (.A1(\ser_C.bit_idx[3] ),
    .A2(_0379_),
    .B1(\ser_C.bit_idx[4] ),
    .Y(_0382_));
 sky130_fd_sc_hd__nor2_1 _1023_ (.A(_0381_),
    .B(_0382_),
    .Y(_0330_));
 sky130_fd_sc_hd__xor2_1 _1024_ (.A(\ser_C.bit_idx[5] ),
    .B(_0381_),
    .X(_0331_));
 sky130_fd_sc_hd__and3_1 _1025_ (.A(\ser_C.bit_idx[5] ),
    .B(\ser_C.bit_idx[6] ),
    .C(_0381_),
    .X(_0383_));
 sky130_fd_sc_hd__a21oi_1 _1026_ (.A1(\ser_C.bit_idx[5] ),
    .A2(_0381_),
    .B1(\ser_C.bit_idx[6] ),
    .Y(_0384_));
 sky130_fd_sc_hd__nor2_1 _1027_ (.A(_0383_),
    .B(_0384_),
    .Y(_0332_));
 sky130_fd_sc_hd__xor2_1 _1028_ (.A(\ser_C.bit_idx[7] ),
    .B(_0383_),
    .X(_0333_));
 sky130_fd_sc_hd__and3_1 _1029_ (.A(\ser_C.bit_idx[7] ),
    .B(\ser_C.bit_idx[8] ),
    .C(_0383_),
    .X(_0385_));
 sky130_fd_sc_hd__a21oi_1 _1030_ (.A1(\ser_C.bit_idx[7] ),
    .A2(_0383_),
    .B1(\ser_C.bit_idx[8] ),
    .Y(_0386_));
 sky130_fd_sc_hd__nor2_1 _1031_ (.A(_0385_),
    .B(_0386_),
    .Y(_0334_));
 sky130_fd_sc_hd__xor2_1 _1032_ (.A(\ser_C.bit_idx[9] ),
    .B(_0385_),
    .X(_0335_));
 sky130_fd_sc_hd__o21ai_1 _1033_ (.A1(_0404_),
    .A2(_0424_),
    .B1(_0348_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2_1 _1034_ (.A(\ser_C.kept_bit_idx[0] ),
    .B(net7),
    .Y(_0387_));
 sky130_fd_sc_hd__or2_1 _1035_ (.A(\ser_C.kept_bit_idx[0] ),
    .B(net7),
    .X(_0388_));
 sky130_fd_sc_hd__and2_1 _1036_ (.A(_0387_),
    .B(_0388_),
    .X(_0337_));
 sky130_fd_sc_hd__xnor2_1 _1037_ (.A(\ser_C.kept_bit_idx[1] ),
    .B(_0387_),
    .Y(_0338_));
 sky130_fd_sc_hd__and4_1 _1038_ (.A(\ser_C.kept_bit_idx[0] ),
    .B(net7),
    .C(\ser_C.kept_bit_idx[1] ),
    .D(\ser_C.kept_bit_idx[2] ),
    .X(_0389_));
 sky130_fd_sc_hd__a31o_1 _1039_ (.A1(\ser_C.kept_bit_idx[0] ),
    .A2(net7),
    .A3(\ser_C.kept_bit_idx[1] ),
    .B1(\ser_C.kept_bit_idx[2] ),
    .X(_0390_));
 sky130_fd_sc_hd__and2b_1 _1040_ (.A_N(_0389_),
    .B(_0390_),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_1 _1041_ (.A(\ser_C.kept_bit_idx[3] ),
    .B(_0389_),
    .Y(_0391_));
 sky130_fd_sc_hd__or2_1 _1042_ (.A(\ser_C.kept_bit_idx[3] ),
    .B(_0389_),
    .X(_0392_));
 sky130_fd_sc_hd__and2_1 _1043_ (.A(_0391_),
    .B(_0392_),
    .X(_0340_));
 sky130_fd_sc_hd__xnor2_1 _1044_ (.A(\ser_C.kept_bit_idx[4] ),
    .B(_0391_),
    .Y(_0341_));
 sky130_fd_sc_hd__and4_1 _1045_ (.A(\ser_C.kept_bit_idx[3] ),
    .B(\ser_C.kept_bit_idx[4] ),
    .C(\ser_C.kept_bit_idx[5] ),
    .D(_0389_),
    .X(_0393_));
 sky130_fd_sc_hd__a31o_1 _1046_ (.A1(\ser_C.kept_bit_idx[3] ),
    .A2(\ser_C.kept_bit_idx[4] ),
    .A3(_0389_),
    .B1(\ser_C.kept_bit_idx[5] ),
    .X(_0394_));
 sky130_fd_sc_hd__and2b_1 _1047_ (.A_N(_0393_),
    .B(_0394_),
    .X(_0342_));
 sky130_fd_sc_hd__xor2_1 _1048_ (.A(\ser_C.kept_bit_idx[6] ),
    .B(_0393_),
    .X(_0343_));
 sky130_fd_sc_hd__and3_1 _1049_ (.A(\ser_C.kept_bit_idx[6] ),
    .B(\ser_C.kept_bit_idx[7] ),
    .C(_0393_),
    .X(_0395_));
 sky130_fd_sc_hd__a21oi_1 _1050_ (.A1(\ser_C.kept_bit_idx[6] ),
    .A2(_0393_),
    .B1(\ser_C.kept_bit_idx[7] ),
    .Y(_0396_));
 sky130_fd_sc_hd__nor2_1 _1051_ (.A(_0395_),
    .B(_0396_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _1052_ (.A(\ser_C.kept_bit_idx[8] ),
    .B(_0395_),
    .Y(_0397_));
 sky130_fd_sc_hd__or2_1 _1053_ (.A(\ser_C.kept_bit_idx[8] ),
    .B(_0395_),
    .X(_0398_));
 sky130_fd_sc_hd__and2_1 _1054_ (.A(_0397_),
    .B(_0398_),
    .X(_0345_));
 sky130_fd_sc_hd__xnor2_1 _1055_ (.A(\ser_C.kept_bit_idx[9] ),
    .B(_0397_),
    .Y(_0346_));
 sky130_fd_sc_hd__dfrtp_1 _1056_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0005_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1057_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0006_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1058_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0007_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1059_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0008_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1060_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0009_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1061_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0010_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1062_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0011_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1063_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0012_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1064_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0013_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1065_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0014_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1066_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0015_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1067_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0016_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1068_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0017_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1069_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0018_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1070_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0019_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1071_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0020_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1072_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0021_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1073_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0022_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1074_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0023_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1075_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0024_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1076_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0025_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1077_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0026_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1078_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0027_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1079_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0028_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1080_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0029_),
    .RESET_B(net5),
    .Q(\systolic_inst.cycle_cnt[24] ));
 sky130_fd_sc_hd__dfrtp_1 _1081_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0030_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[25] ));
 sky130_fd_sc_hd__dfrtp_1 _1082_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0031_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[26] ));
 sky130_fd_sc_hd__dfrtp_1 _1083_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0032_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1084_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0033_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1085_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0034_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1086_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0035_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1087_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0036_),
    .RESET_B(net15),
    .Q(\systolic_inst.cycle_cnt[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1088_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0037_),
    .RESET_B(net14),
    .Q(\deser_A.bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1089_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0038_),
    .RESET_B(net14),
    .Q(\deser_A.bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1090_ (.CLK(clknet_4_8_0_A_in_serial_clk),
    .D(_0039_),
    .RESET_B(net14),
    .Q(\deser_A.bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1091_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0040_),
    .RESET_B(net14),
    .Q(\deser_A.bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1092_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0041_),
    .RESET_B(net14),
    .Q(\deser_A.bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1093_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0042_),
    .RESET_B(net14),
    .Q(\deser_A.bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1094_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0043_),
    .RESET_B(net14),
    .Q(\deser_A.bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1095_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0044_),
    .RESET_B(net14),
    .Q(\deser_A.bit_idx[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1096_ (.CLK(clknet_4_8_0_A_in_serial_clk),
    .D(_0045_),
    .RESET_B(net14),
    .Q(\deser_A.kept_bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0046_),
    .RESET_B(net14),
    .Q(\deser_A.kept_bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1098_ (.CLK(clknet_4_9_0_A_in_serial_clk),
    .D(_0047_),
    .RESET_B(net14),
    .Q(\deser_A.kept_bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1099_ (.CLK(clknet_4_9_0_A_in_serial_clk),
    .D(_0048_),
    .RESET_B(net14),
    .Q(\deser_A.kept_bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1100_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0049_),
    .RESET_B(net14),
    .Q(\deser_A.kept_bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1101_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0050_),
    .RESET_B(net14),
    .Q(\deser_A.kept_bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0051_),
    .RESET_B(net14),
    .Q(\deser_A.kept_bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0052_),
    .RESET_B(net14),
    .Q(\deser_A.kept_bit_idx[7] ));
 sky130_fd_sc_hd__dfrtp_4 _1104_ (.CLK(clknet_4_10_0_A_in_serial_clk),
    .D(_0000_),
    .RESET_B(net14),
    .Q(\deser_A.receiving ));
 sky130_fd_sc_hd__dfrtp_1 _1105_ (.CLK(clknet_4_8_0_A_in_serial_clk),
    .D(_0053_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1106_ (.CLK(clknet_4_8_0_A_in_serial_clk),
    .D(_0054_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1107_ (.CLK(clknet_4_8_0_A_in_serial_clk),
    .D(_0055_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1108_ (.CLK(clknet_4_8_0_A_in_serial_clk),
    .D(_0056_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1109_ (.CLK(clknet_4_9_0_A_in_serial_clk),
    .D(_0057_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1110_ (.CLK(clknet_4_9_0_A_in_serial_clk),
    .D(_0058_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1111_ (.CLK(clknet_4_9_0_A_in_serial_clk),
    .D(_0059_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_4_9_0_A_in_serial_clk),
    .D(_0060_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1113_ (.CLK(clknet_4_9_0_A_in_serial_clk),
    .D(_0061_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1114_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0062_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1115_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0063_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1116_ (.CLK(clknet_4_14_0_A_in_serial_clk),
    .D(_0064_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1117_ (.CLK(clknet_4_14_0_A_in_serial_clk),
    .D(_0065_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1118_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0066_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1119_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0067_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_4_14_0_A_in_serial_clk),
    .D(_0068_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1121_ (.CLK(clknet_4_14_0_A_in_serial_clk),
    .D(_0069_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1122_ (.CLK(clknet_4_14_0_A_in_serial_clk),
    .D(_0070_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1123_ (.CLK(clknet_4_14_0_A_in_serial_clk),
    .D(_0071_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1124_ (.CLK(clknet_4_12_0_A_in_serial_clk),
    .D(_0072_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_4_12_0_A_in_serial_clk),
    .D(_0073_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_4_12_0_A_in_serial_clk),
    .D(_0074_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_4_12_0_A_in_serial_clk),
    .D(_0075_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_4_12_0_A_in_serial_clk),
    .D(_0076_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[24] ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(clknet_4_12_0_A_in_serial_clk),
    .D(_0077_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[25] ));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(clknet_4_6_0_A_in_serial_clk),
    .D(_0078_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[26] ));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(clknet_4_6_0_A_in_serial_clk),
    .D(_0079_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1132_ (.CLK(clknet_4_3_0_A_in_serial_clk),
    .D(_0080_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1133_ (.CLK(clknet_4_3_0_A_in_serial_clk),
    .D(_0081_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(clknet_4_3_0_A_in_serial_clk),
    .D(_0082_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(clknet_4_3_0_A_in_serial_clk),
    .D(_0083_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0084_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[32] ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0085_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[33] ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0086_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[34] ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0087_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[35] ));
 sky130_fd_sc_hd__dfrtp_1 _1140_ (.CLK(clknet_4_3_0_A_in_serial_clk),
    .D(_0088_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[36] ));
 sky130_fd_sc_hd__dfrtp_1 _1141_ (.CLK(clknet_4_3_0_A_in_serial_clk),
    .D(_0089_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[37] ));
 sky130_fd_sc_hd__dfrtp_1 _1142_ (.CLK(clknet_4_3_0_A_in_serial_clk),
    .D(_0090_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[38] ));
 sky130_fd_sc_hd__dfrtp_1 _1143_ (.CLK(clknet_4_3_0_A_in_serial_clk),
    .D(_0091_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[39] ));
 sky130_fd_sc_hd__dfrtp_1 _1144_ (.CLK(clknet_4_6_0_A_in_serial_clk),
    .D(_0092_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[40] ));
 sky130_fd_sc_hd__dfrtp_1 _1145_ (.CLK(clknet_4_6_0_A_in_serial_clk),
    .D(_0093_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[41] ));
 sky130_fd_sc_hd__dfrtp_1 _1146_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0094_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[42] ));
 sky130_fd_sc_hd__dfrtp_1 _1147_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0095_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[43] ));
 sky130_fd_sc_hd__dfrtp_1 _1148_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0096_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[44] ));
 sky130_fd_sc_hd__dfrtp_1 _1149_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0097_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[45] ));
 sky130_fd_sc_hd__dfrtp_1 _1150_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0098_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[46] ));
 sky130_fd_sc_hd__dfrtp_1 _1151_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0099_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[47] ));
 sky130_fd_sc_hd__dfrtp_1 _1152_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0100_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[48] ));
 sky130_fd_sc_hd__dfrtp_1 _1153_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0101_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[49] ));
 sky130_fd_sc_hd__dfrtp_1 _1154_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0102_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[50] ));
 sky130_fd_sc_hd__dfrtp_1 _1155_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0103_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[51] ));
 sky130_fd_sc_hd__dfrtp_1 _1156_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0104_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[52] ));
 sky130_fd_sc_hd__dfrtp_1 _1157_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0105_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[53] ));
 sky130_fd_sc_hd__dfrtp_1 _1158_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0106_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[54] ));
 sky130_fd_sc_hd__dfrtp_1 _1159_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0107_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[55] ));
 sky130_fd_sc_hd__dfrtp_1 _1160_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0108_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[56] ));
 sky130_fd_sc_hd__dfrtp_1 _1161_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0109_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[57] ));
 sky130_fd_sc_hd__dfrtp_1 _1162_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0110_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[58] ));
 sky130_fd_sc_hd__dfrtp_1 _1163_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0111_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[59] ));
 sky130_fd_sc_hd__dfrtp_1 _1164_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0112_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[60] ));
 sky130_fd_sc_hd__dfrtp_1 _1165_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0113_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[61] ));
 sky130_fd_sc_hd__dfrtp_1 _1166_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0114_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[62] ));
 sky130_fd_sc_hd__dfrtp_1 _1167_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0115_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[63] ));
 sky130_fd_sc_hd__dfrtp_1 _1168_ (.CLK(clknet_4_14_0_A_in_serial_clk),
    .D(_0116_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[64] ));
 sky130_fd_sc_hd__dfrtp_1 _1169_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0117_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[65] ));
 sky130_fd_sc_hd__dfrtp_1 _1170_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0118_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[66] ));
 sky130_fd_sc_hd__dfrtp_1 _1171_ (.CLK(clknet_4_14_0_A_in_serial_clk),
    .D(_0119_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[67] ));
 sky130_fd_sc_hd__dfrtp_1 _1172_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0120_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[68] ));
 sky130_fd_sc_hd__dfrtp_1 _1173_ (.CLK(clknet_4_15_0_A_in_serial_clk),
    .D(_0121_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[69] ));
 sky130_fd_sc_hd__dfrtp_1 _1174_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0122_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[70] ));
 sky130_fd_sc_hd__dfrtp_1 _1175_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0123_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[71] ));
 sky130_fd_sc_hd__dfrtp_1 _1176_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0124_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[72] ));
 sky130_fd_sc_hd__dfrtp_1 _1177_ (.CLK(clknet_4_13_0_A_in_serial_clk),
    .D(_0125_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[73] ));
 sky130_fd_sc_hd__dfrtp_1 _1178_ (.CLK(clknet_4_12_0_A_in_serial_clk),
    .D(_0126_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[74] ));
 sky130_fd_sc_hd__dfrtp_1 _1179_ (.CLK(clknet_4_6_0_A_in_serial_clk),
    .D(_0127_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[75] ));
 sky130_fd_sc_hd__dfrtp_1 _1180_ (.CLK(clknet_4_7_0_A_in_serial_clk),
    .D(_0128_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[76] ));
 sky130_fd_sc_hd__dfrtp_1 _1181_ (.CLK(clknet_4_6_0_A_in_serial_clk),
    .D(_0129_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[77] ));
 sky130_fd_sc_hd__dfrtp_1 _1182_ (.CLK(clknet_4_6_0_A_in_serial_clk),
    .D(_0130_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[78] ));
 sky130_fd_sc_hd__dfrtp_1 _1183_ (.CLK(clknet_4_6_0_A_in_serial_clk),
    .D(_0131_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[79] ));
 sky130_fd_sc_hd__dfrtp_1 _1184_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0132_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[80] ));
 sky130_fd_sc_hd__dfrtp_1 _1185_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0133_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[81] ));
 sky130_fd_sc_hd__dfrtp_1 _1186_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0134_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[82] ));
 sky130_fd_sc_hd__dfrtp_1 _1187_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0135_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[83] ));
 sky130_fd_sc_hd__dfrtp_1 _1188_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0136_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[84] ));
 sky130_fd_sc_hd__dfrtp_1 _1189_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0137_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[85] ));
 sky130_fd_sc_hd__dfrtp_1 _1190_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0138_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[86] ));
 sky130_fd_sc_hd__dfrtp_1 _1191_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0139_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[87] ));
 sky130_fd_sc_hd__dfrtp_1 _1192_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0140_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[88] ));
 sky130_fd_sc_hd__dfrtp_1 _1193_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0141_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[89] ));
 sky130_fd_sc_hd__dfrtp_1 _1194_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0142_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[90] ));
 sky130_fd_sc_hd__dfrtp_1 _1195_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0143_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[91] ));
 sky130_fd_sc_hd__dfrtp_1 _1196_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0144_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[92] ));
 sky130_fd_sc_hd__dfrtp_1 _1197_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0145_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[93] ));
 sky130_fd_sc_hd__dfrtp_1 _1198_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0146_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[94] ));
 sky130_fd_sc_hd__dfrtp_1 _1199_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0147_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[95] ));
 sky130_fd_sc_hd__dfrtp_1 _1200_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0148_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[96] ));
 sky130_fd_sc_hd__dfrtp_1 _1201_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0149_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[97] ));
 sky130_fd_sc_hd__dfrtp_1 _1202_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0150_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[98] ));
 sky130_fd_sc_hd__dfrtp_1 _1203_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0151_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[99] ));
 sky130_fd_sc_hd__dfrtp_1 _1204_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0152_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[100] ));
 sky130_fd_sc_hd__dfrtp_1 _1205_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0153_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[101] ));
 sky130_fd_sc_hd__dfrtp_1 _1206_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0154_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[102] ));
 sky130_fd_sc_hd__dfrtp_1 _1207_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0155_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[103] ));
 sky130_fd_sc_hd__dfrtp_1 _1208_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0156_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[104] ));
 sky130_fd_sc_hd__dfrtp_1 _1209_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0157_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[105] ));
 sky130_fd_sc_hd__dfrtp_1 _1210_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0158_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[106] ));
 sky130_fd_sc_hd__dfrtp_1 _1211_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0159_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[107] ));
 sky130_fd_sc_hd__dfrtp_1 _1212_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0160_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[108] ));
 sky130_fd_sc_hd__dfrtp_1 _1213_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0161_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[109] ));
 sky130_fd_sc_hd__dfrtp_1 _1214_ (.CLK(clknet_4_5_0_A_in_serial_clk),
    .D(_0162_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[110] ));
 sky130_fd_sc_hd__dfrtp_1 _1215_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0163_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[111] ));
 sky130_fd_sc_hd__dfrtp_1 _1216_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0164_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[112] ));
 sky130_fd_sc_hd__dfrtp_1 _1217_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0165_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[113] ));
 sky130_fd_sc_hd__dfrtp_1 _1218_ (.CLK(clknet_4_4_0_A_in_serial_clk),
    .D(_0166_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[114] ));
 sky130_fd_sc_hd__dfrtp_1 _1219_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0167_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[115] ));
 sky130_fd_sc_hd__dfrtp_1 _1220_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0168_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[116] ));
 sky130_fd_sc_hd__dfrtp_1 _1221_ (.CLK(clknet_4_1_0_A_in_serial_clk),
    .D(_0169_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[117] ));
 sky130_fd_sc_hd__dfrtp_1 _1222_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0170_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[118] ));
 sky130_fd_sc_hd__dfrtp_1 _1223_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0171_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[119] ));
 sky130_fd_sc_hd__dfrtp_1 _1224_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0172_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[120] ));
 sky130_fd_sc_hd__dfrtp_1 _1225_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0173_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[121] ));
 sky130_fd_sc_hd__dfrtp_1 _1226_ (.CLK(clknet_4_0_0_A_in_serial_clk),
    .D(_0174_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[122] ));
 sky130_fd_sc_hd__dfrtp_1 _1227_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0175_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[123] ));
 sky130_fd_sc_hd__dfrtp_1 _1228_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0176_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[124] ));
 sky130_fd_sc_hd__dfrtp_1 _1229_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0177_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[125] ));
 sky130_fd_sc_hd__dfrtp_1 _1230_ (.CLK(clknet_4_8_0_A_in_serial_clk),
    .D(_0178_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[126] ));
 sky130_fd_sc_hd__dfrtp_1 _1231_ (.CLK(clknet_4_2_0_A_in_serial_clk),
    .D(_0179_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[127] ));
 sky130_fd_sc_hd__dfrtp_1 _1232_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0180_),
    .RESET_B(net15),
    .Q(\deser_B.bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1233_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0181_),
    .RESET_B(net15),
    .Q(\deser_B.bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1234_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0182_),
    .RESET_B(net15),
    .Q(\deser_B.bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1235_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0183_),
    .RESET_B(net15),
    .Q(\deser_B.bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1236_ (.CLK(clknet_4_12_0_B_in_serial_clk),
    .D(_0184_),
    .RESET_B(net15),
    .Q(\deser_B.bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1237_ (.CLK(clknet_4_15_0_B_in_serial_clk),
    .D(_0185_),
    .RESET_B(net15),
    .Q(\deser_B.bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1238_ (.CLK(clknet_4_15_0_B_in_serial_clk),
    .D(_0186_),
    .RESET_B(net15),
    .Q(\deser_B.bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1239_ (.CLK(clknet_4_14_0_B_in_serial_clk),
    .D(_0187_),
    .RESET_B(net15),
    .Q(\deser_B.bit_idx[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1240_ (.CLK(clknet_4_15_0_B_in_serial_clk),
    .D(_0188_),
    .RESET_B(net15),
    .Q(\deser_B.kept_bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1241_ (.CLK(clknet_4_15_0_B_in_serial_clk),
    .D(_0189_),
    .RESET_B(net15),
    .Q(\deser_B.kept_bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1242_ (.CLK(clknet_4_15_0_B_in_serial_clk),
    .D(_0190_),
    .RESET_B(net15),
    .Q(\deser_B.kept_bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1243_ (.CLK(clknet_4_15_0_B_in_serial_clk),
    .D(_0191_),
    .RESET_B(net15),
    .Q(\deser_B.kept_bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1244_ (.CLK(clknet_4_15_0_B_in_serial_clk),
    .D(_0192_),
    .RESET_B(net15),
    .Q(\deser_B.kept_bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1245_ (.CLK(clknet_4_15_0_B_in_serial_clk),
    .D(_0193_),
    .RESET_B(net15),
    .Q(\deser_B.kept_bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1246_ (.CLK(clknet_4_14_0_B_in_serial_clk),
    .D(_0194_),
    .RESET_B(net15),
    .Q(\deser_B.kept_bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1247_ (.CLK(clknet_4_14_0_B_in_serial_clk),
    .D(_0195_),
    .RESET_B(net15),
    .Q(\deser_B.kept_bit_idx[7] ));
 sky130_fd_sc_hd__dfrtp_4 _1248_ (.CLK(clknet_4_14_0_B_in_serial_clk),
    .D(_0001_),
    .RESET_B(net15),
    .Q(\deser_B.receiving ));
 sky130_fd_sc_hd__dfrtp_1 _1249_ (.CLK(clknet_4_11_0_A_in_serial_clk),
    .D(_0196_),
    .RESET_B(net14),
    .Q(\deser_A.kept_receiving ));
 sky130_fd_sc_hd__dfrtp_1 _1250_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0197_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1251_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0198_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1252_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0199_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1253_ (.CLK(clknet_4_12_0_B_in_serial_clk),
    .D(_0200_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1254_ (.CLK(clknet_4_12_0_B_in_serial_clk),
    .D(_0201_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1255_ (.CLK(clknet_4_12_0_B_in_serial_clk),
    .D(_0202_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1256_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0203_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1257_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0204_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1258_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0205_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1259_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0206_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1260_ (.CLK(clknet_4_14_0_B_in_serial_clk),
    .D(_0207_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1261_ (.CLK(clknet_4_14_0_B_in_serial_clk),
    .D(_0208_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1262_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0209_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1263_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0210_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1264_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0211_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1265_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0212_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1266_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0213_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1267_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0214_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1268_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0215_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1269_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0216_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1270_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0217_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1271_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0218_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1272_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0219_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1273_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0220_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[24] ));
 sky130_fd_sc_hd__dfrtp_1 _1274_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0221_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[25] ));
 sky130_fd_sc_hd__dfrtp_1 _1275_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0222_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[26] ));
 sky130_fd_sc_hd__dfrtp_1 _1276_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0223_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1277_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0224_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1278_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0225_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1279_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0226_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1280_ (.CLK(clknet_4_3_0_B_in_serial_clk),
    .D(_0227_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1281_ (.CLK(clknet_4_3_0_B_in_serial_clk),
    .D(_0228_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[32] ));
 sky130_fd_sc_hd__dfrtp_1 _1282_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0229_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[33] ));
 sky130_fd_sc_hd__dfrtp_1 _1283_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0230_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[34] ));
 sky130_fd_sc_hd__dfrtp_1 _1284_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0231_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[35] ));
 sky130_fd_sc_hd__dfrtp_1 _1285_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0232_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[36] ));
 sky130_fd_sc_hd__dfrtp_1 _1286_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0233_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[37] ));
 sky130_fd_sc_hd__dfrtp_1 _1287_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0234_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[38] ));
 sky130_fd_sc_hd__dfrtp_1 _1288_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0235_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[39] ));
 sky130_fd_sc_hd__dfrtp_1 _1289_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0236_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[40] ));
 sky130_fd_sc_hd__dfrtp_1 _1290_ (.CLK(clknet_4_11_0_B_in_serial_clk),
    .D(_0237_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[41] ));
 sky130_fd_sc_hd__dfrtp_1 _1291_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0238_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[42] ));
 sky130_fd_sc_hd__dfrtp_1 _1292_ (.CLK(clknet_4_10_0_B_in_serial_clk),
    .D(_0239_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[43] ));
 sky130_fd_sc_hd__dfrtp_1 _1293_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0240_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[44] ));
 sky130_fd_sc_hd__dfrtp_1 _1294_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0241_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[45] ));
 sky130_fd_sc_hd__dfrtp_1 _1295_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0242_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[46] ));
 sky130_fd_sc_hd__dfrtp_1 _1296_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0243_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[47] ));
 sky130_fd_sc_hd__dfrtp_1 _1297_ (.CLK(clknet_4_8_0_B_in_serial_clk),
    .D(_0244_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[48] ));
 sky130_fd_sc_hd__dfrtp_1 _1298_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0245_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[49] ));
 sky130_fd_sc_hd__dfrtp_1 _1299_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0246_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[50] ));
 sky130_fd_sc_hd__dfrtp_1 _1300_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0247_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[51] ));
 sky130_fd_sc_hd__dfrtp_1 _1301_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0248_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[52] ));
 sky130_fd_sc_hd__dfrtp_1 _1302_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0249_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[53] ));
 sky130_fd_sc_hd__dfrtp_1 _1303_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0250_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[54] ));
 sky130_fd_sc_hd__dfrtp_1 _1304_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0251_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[55] ));
 sky130_fd_sc_hd__dfrtp_1 _1305_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0252_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[56] ));
 sky130_fd_sc_hd__dfrtp_1 _1306_ (.CLK(clknet_4_1_0_B_in_serial_clk),
    .D(_0253_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[57] ));
 sky130_fd_sc_hd__dfrtp_1 _1307_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0254_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[58] ));
 sky130_fd_sc_hd__dfrtp_1 _1308_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0255_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[59] ));
 sky130_fd_sc_hd__dfrtp_1 _1309_ (.CLK(clknet_4_2_0_B_in_serial_clk),
    .D(_0256_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[60] ));
 sky130_fd_sc_hd__dfrtp_1 _1310_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0257_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[61] ));
 sky130_fd_sc_hd__dfrtp_1 _1311_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0258_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[62] ));
 sky130_fd_sc_hd__dfrtp_1 _1312_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0259_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[63] ));
 sky130_fd_sc_hd__dfrtp_1 _1313_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0260_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[64] ));
 sky130_fd_sc_hd__dfrtp_1 _1314_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0261_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[65] ));
 sky130_fd_sc_hd__dfrtp_1 _1315_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0262_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[66] ));
 sky130_fd_sc_hd__dfrtp_1 _1316_ (.CLK(clknet_4_0_0_B_in_serial_clk),
    .D(_0263_),
    .RESET_B(net14),
    .Q(\deser_B.kept_shift_reg[67] ));
 sky130_fd_sc_hd__dfrtp_1 _1317_ (.CLK(clknet_4_1_0_B_in_serial_clk),
    .D(_0264_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[68] ));
 sky130_fd_sc_hd__dfrtp_1 _1318_ (.CLK(clknet_4_1_0_B_in_serial_clk),
    .D(_0265_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[69] ));
 sky130_fd_sc_hd__dfrtp_1 _1319_ (.CLK(clknet_4_1_0_B_in_serial_clk),
    .D(_0266_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[70] ));
 sky130_fd_sc_hd__dfrtp_1 _1320_ (.CLK(clknet_4_1_0_B_in_serial_clk),
    .D(_0267_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[71] ));
 sky130_fd_sc_hd__dfrtp_1 _1321_ (.CLK(clknet_4_1_0_B_in_serial_clk),
    .D(_0268_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[72] ));
 sky130_fd_sc_hd__dfrtp_1 _1322_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0269_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[73] ));
 sky130_fd_sc_hd__dfrtp_1 _1323_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0270_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[74] ));
 sky130_fd_sc_hd__dfrtp_1 _1324_ (.CLK(clknet_4_1_0_B_in_serial_clk),
    .D(_0271_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[75] ));
 sky130_fd_sc_hd__dfrtp_1 _1325_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0272_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[76] ));
 sky130_fd_sc_hd__dfrtp_1 _1326_ (.CLK(clknet_4_1_0_B_in_serial_clk),
    .D(_0273_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[77] ));
 sky130_fd_sc_hd__dfrtp_1 _1327_ (.CLK(clknet_4_3_0_B_in_serial_clk),
    .D(_0274_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[78] ));
 sky130_fd_sc_hd__dfrtp_1 _1328_ (.CLK(clknet_4_3_0_B_in_serial_clk),
    .D(_0275_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[79] ));
 sky130_fd_sc_hd__dfrtp_1 _1329_ (.CLK(clknet_4_3_0_B_in_serial_clk),
    .D(_0276_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[80] ));
 sky130_fd_sc_hd__dfrtp_1 _1330_ (.CLK(clknet_4_3_0_B_in_serial_clk),
    .D(_0277_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[81] ));
 sky130_fd_sc_hd__dfrtp_1 _1331_ (.CLK(clknet_4_3_0_B_in_serial_clk),
    .D(_0278_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[82] ));
 sky130_fd_sc_hd__dfrtp_1 _1332_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0279_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[83] ));
 sky130_fd_sc_hd__dfrtp_1 _1333_ (.CLK(clknet_4_12_0_B_in_serial_clk),
    .D(_0280_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[84] ));
 sky130_fd_sc_hd__dfrtp_1 _1334_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0281_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[85] ));
 sky130_fd_sc_hd__dfrtp_1 _1335_ (.CLK(clknet_4_9_0_B_in_serial_clk),
    .D(_0282_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[86] ));
 sky130_fd_sc_hd__dfrtp_1 _1336_ (.CLK(clknet_4_12_0_B_in_serial_clk),
    .D(_0283_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[87] ));
 sky130_fd_sc_hd__dfrtp_1 _1337_ (.CLK(clknet_4_12_0_B_in_serial_clk),
    .D(_0284_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[88] ));
 sky130_fd_sc_hd__dfrtp_1 _1338_ (.CLK(clknet_4_6_0_B_in_serial_clk),
    .D(_0285_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[89] ));
 sky130_fd_sc_hd__dfrtp_1 _1339_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0286_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[90] ));
 sky130_fd_sc_hd__dfrtp_1 _1340_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0287_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[91] ));
 sky130_fd_sc_hd__dfrtp_1 _1341_ (.CLK(clknet_4_6_0_B_in_serial_clk),
    .D(_0288_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[92] ));
 sky130_fd_sc_hd__dfrtp_1 _1342_ (.CLK(clknet_4_6_0_B_in_serial_clk),
    .D(_0289_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[93] ));
 sky130_fd_sc_hd__dfrtp_1 _1343_ (.CLK(clknet_4_6_0_B_in_serial_clk),
    .D(_0290_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[94] ));
 sky130_fd_sc_hd__dfrtp_1 _1344_ (.CLK(clknet_4_6_0_B_in_serial_clk),
    .D(_0291_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[95] ));
 sky130_fd_sc_hd__dfrtp_1 _1345_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0292_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[96] ));
 sky130_fd_sc_hd__dfrtp_1 _1346_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0293_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[97] ));
 sky130_fd_sc_hd__dfrtp_1 _1347_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0294_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[98] ));
 sky130_fd_sc_hd__dfrtp_1 _1348_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0295_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[99] ));
 sky130_fd_sc_hd__dfrtp_1 _1349_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0296_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[100] ));
 sky130_fd_sc_hd__dfrtp_1 _1350_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0297_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[101] ));
 sky130_fd_sc_hd__dfrtp_1 _1351_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0298_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[102] ));
 sky130_fd_sc_hd__dfrtp_1 _1352_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0299_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[103] ));
 sky130_fd_sc_hd__dfrtp_1 _1353_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0300_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[104] ));
 sky130_fd_sc_hd__dfrtp_1 _1354_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0301_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[105] ));
 sky130_fd_sc_hd__dfrtp_1 _1355_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0302_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[106] ));
 sky130_fd_sc_hd__dfrtp_1 _1356_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0303_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[107] ));
 sky130_fd_sc_hd__dfrtp_1 _1357_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0304_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[108] ));
 sky130_fd_sc_hd__dfrtp_1 _1358_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0305_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[109] ));
 sky130_fd_sc_hd__dfrtp_1 _1359_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0306_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[110] ));
 sky130_fd_sc_hd__dfrtp_1 _1360_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0307_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[111] ));
 sky130_fd_sc_hd__dfrtp_1 _1361_ (.CLK(clknet_4_4_0_B_in_serial_clk),
    .D(_0308_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[112] ));
 sky130_fd_sc_hd__dfrtp_1 _1362_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0309_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[113] ));
 sky130_fd_sc_hd__dfrtp_1 _1363_ (.CLK(clknet_4_6_0_B_in_serial_clk),
    .D(_0310_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[114] ));
 sky130_fd_sc_hd__dfrtp_1 _1364_ (.CLK(clknet_4_6_0_B_in_serial_clk),
    .D(_0311_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[115] ));
 sky130_fd_sc_hd__dfrtp_1 _1365_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0312_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[116] ));
 sky130_fd_sc_hd__dfrtp_1 _1366_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0313_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[117] ));
 sky130_fd_sc_hd__dfrtp_1 _1367_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0314_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[118] ));
 sky130_fd_sc_hd__dfrtp_1 _1368_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0315_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[119] ));
 sky130_fd_sc_hd__dfrtp_1 _1369_ (.CLK(clknet_4_5_0_B_in_serial_clk),
    .D(_0316_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[120] ));
 sky130_fd_sc_hd__dfrtp_1 _1370_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0317_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[121] ));
 sky130_fd_sc_hd__dfrtp_1 _1371_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0318_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[122] ));
 sky130_fd_sc_hd__dfrtp_1 _1372_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0319_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[123] ));
 sky130_fd_sc_hd__dfrtp_1 _1373_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0320_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[124] ));
 sky130_fd_sc_hd__dfrtp_1 _1374_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0321_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[125] ));
 sky130_fd_sc_hd__dfrtp_1 _1375_ (.CLK(clknet_4_7_0_B_in_serial_clk),
    .D(_0322_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[126] ));
 sky130_fd_sc_hd__dfrtp_1 _1376_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0323_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[127] ));
 sky130_fd_sc_hd__dfrtp_1 _1377_ (.CLK(clknet_4_13_0_B_in_serial_clk),
    .D(_0324_),
    .RESET_B(net15),
    .Q(\deser_B.kept_shift_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1378_ (.CLK(clknet_4_8_0_A_in_serial_clk),
    .D(_0325_),
    .RESET_B(net14),
    .Q(\deser_A.kept_shift_reg[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1379_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0004_),
    .RESET_B(net5),
    .Q(\systolic_inst.ce_local ));
 sky130_fd_sc_hd__dfrtp_1 _1380_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0003_),
    .RESET_B(net5),
    .Q(net9));
 sky130_fd_sc_hd__dfrtp_1 _1381_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0326_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1382_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0327_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1383_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0328_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1384_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0329_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1385_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0330_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1386_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0331_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1387_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0332_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1388_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0333_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1389_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0334_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1390_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0335_),
    .RESET_B(net5),
    .Q(\ser_C.bit_idx[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1391_ (.CLK(clknet_4_14_0_B_in_serial_clk),
    .D(_0336_),
    .RESET_B(net15),
    .Q(\deser_B.kept_receiving ));
 sky130_fd_sc_hd__dfrtp_4 _1392_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0002_),
    .RESET_B(net5),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _1393_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0337_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1394_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0338_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1395_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0339_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1396_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0340_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1397_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0341_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1398_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0342_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1399_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0343_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1400_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0344_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1401_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0345_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1402_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0346_),
    .RESET_B(net5),
    .Q(\ser_C.kept_bit_idx[9] ));
 sky130_fd_sc_hd__clkinv_4 clkload29 (.A(clknet_4_15_0_B_in_serial_clk));
 sky130_fd_sc_hd__inv_6 clkload28 (.A(clknet_4_14_0_B_in_serial_clk));
 sky130_fd_sc_hd__bufinv_16 clkload27 (.A(clknet_4_13_0_B_in_serial_clk));
 sky130_fd_sc_hd__inv_6 clkload26 (.A(clknet_4_12_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkinv_2 clkload25 (.A(clknet_4_11_0_B_in_serial_clk));
 sky130_fd_sc_hd__bufinv_16 clkload24 (.A(clknet_4_10_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload23 (.A(clknet_4_9_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload22 (.A(clknet_4_8_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload21 (.A(clknet_4_7_0_B_in_serial_clk));
 sky130_fd_sc_hd__inv_6 clkload20 (.A(clknet_4_6_0_B_in_serial_clk));
 sky130_fd_sc_hd__bufinv_16 clkload19 (.A(clknet_4_4_0_B_in_serial_clk));
 sky130_fd_sc_hd__inv_6 clkload18 (.A(clknet_4_3_0_B_in_serial_clk));
 sky130_fd_sc_hd__bufinv_16 clkload17 (.A(clknet_4_2_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkinv_4 clkload16 (.A(clknet_4_1_0_B_in_serial_clk));
 sky130_fd_sc_hd__bufinv_16 clkload15 (.A(clknet_4_0_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_15_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_14_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_13_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_12_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_11_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_10_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_9_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_8_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_7_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_6_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_5_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_4_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_3_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_2_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_1_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_B_in_serial_clk (.A(clknet_0_B_in_serial_clk),
    .X(clknet_4_0_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_B_in_serial_clk (.A(B_in_serial_clk),
    .X(clknet_0_B_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload14 (.A(clknet_4_15_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_4_14_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload12 (.A(clknet_4_13_0_A_in_serial_clk));
 sky130_fd_sc_hd__bufinv_16 clkload11 (.A(clknet_4_12_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_4_11_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload9 (.A(clknet_4_10_0_A_in_serial_clk));
 sky130_fd_sc_hd__bufinv_16 clkload8 (.A(clknet_4_9_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_4_8_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkinv_2 clkload6 (.A(clknet_4_6_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload5 (.A(clknet_4_4_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_4_3_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_4_1_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_15_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_14_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_13_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_12_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_11_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_10_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_9_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_8_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_7_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_6_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_5_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_4_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_3_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_2_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_1_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_A_in_serial_clk (.A(clknet_0_A_in_serial_clk),
    .X(clknet_4_0_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_A_in_serial_clk (.A(A_in_serial_clk),
    .X(clknet_0_A_in_serial_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__inv_4 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_2 _1917_ (.A(clknet_2_0__leaf_clk),
    .X(net8));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_573 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(A_in_frame_sync),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(A_in_serial_data),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(B_in_frame_sync),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(B_in_serial_data),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(rst_n),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(start),
    .X(net6));
 sky130_fd_sc_hd__buf_1 output7 (.A(net7),
    .X(C_out_frame_sync));
 sky130_fd_sc_hd__buf_1 output8 (.A(net8),
    .X(C_out_serial_clk));
 sky130_fd_sc_hd__buf_1 output9 (.A(net9),
    .X(done));
 sky130_fd_sc_hd__buf_12 max_cap10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__buf_12 max_cap11 (.A(\deser_B.receiving ),
    .X(net11));
 sky130_fd_sc_hd__buf_12 max_cap12 (.A(\deser_A.receiving ),
    .X(net12));
 sky130_fd_sc_hd__buf_12 max_cap13 (.A(\deser_A.receiving ),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_16 load_slew14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_16 load_slew15 (.A(net5),
    .X(net15));
 sky130_fd_sc_hd__conb_1 Systolic4x4_serial_io_16 (.LO(net16));
 assign C_out_serial_data = net16;
endmodule
