magic
tech sky130A
magscale 1 2
timestamp 1757868665
<< checkpaint >>
rect -3932 -3932 42140 44284
<< viali >>
rect 32137 37893 32171 37927
rect 32353 37893 32387 37927
rect 13553 37825 13587 37859
rect 16037 37825 16071 37859
rect 16129 37825 16163 37859
rect 18613 37825 18647 37859
rect 23581 37825 23615 37859
rect 25237 37825 25271 37859
rect 27445 37825 27479 37859
rect 29745 37825 29779 37859
rect 30757 37825 30791 37859
rect 31769 37825 31803 37859
rect 13645 37757 13679 37791
rect 13737 37757 13771 37791
rect 16313 37757 16347 37791
rect 18705 37757 18739 37791
rect 18889 37757 18923 37791
rect 23673 37757 23707 37791
rect 23765 37757 23799 37791
rect 27537 37757 27571 37791
rect 29193 37757 29227 37791
rect 30021 37757 30055 37791
rect 30941 37757 30975 37791
rect 31493 37757 31527 37791
rect 31677 37689 31711 37723
rect 13185 37621 13219 37655
rect 15669 37621 15703 37655
rect 18245 37621 18279 37655
rect 23213 37621 23247 37655
rect 25421 37621 25455 37655
rect 27261 37621 27295 37655
rect 28733 37621 28767 37655
rect 31585 37621 31619 37655
rect 32321 37621 32355 37655
rect 32505 37621 32539 37655
rect 14749 37417 14783 37451
rect 18981 37417 19015 37451
rect 24409 37417 24443 37451
rect 28089 37417 28123 37451
rect 31585 37417 31619 37451
rect 23857 37349 23891 37383
rect 13461 37281 13495 37315
rect 16221 37281 16255 37315
rect 17509 37281 17543 37315
rect 19441 37281 19475 37315
rect 22385 37281 22419 37315
rect 30113 37281 30147 37315
rect 1409 37213 1443 37247
rect 13737 37213 13771 37247
rect 16497 37213 16531 37247
rect 17233 37213 17267 37247
rect 21833 37213 21867 37247
rect 22109 37213 22143 37247
rect 26157 37213 26191 37247
rect 26249 37213 26283 37247
rect 28273 37213 28307 37247
rect 28549 37213 28583 37247
rect 28733 37213 28767 37247
rect 29837 37213 29871 37247
rect 31677 37213 31711 37247
rect 2605 37145 2639 37179
rect 19533 37145 19567 37179
rect 21557 37145 21591 37179
rect 25881 37145 25915 37179
rect 26525 37145 26559 37179
rect 29285 37145 29319 37179
rect 31953 37145 31987 37179
rect 11989 37077 12023 37111
rect 19625 37077 19659 37111
rect 19993 37077 20027 37111
rect 20085 37077 20119 37111
rect 27997 37077 28031 37111
rect 28457 37077 28491 37111
rect 33425 37077 33459 37111
rect 12541 36873 12575 36907
rect 16497 36873 16531 36907
rect 17049 36873 17083 36907
rect 18429 36873 18463 36907
rect 18797 36873 18831 36907
rect 24777 36873 24811 36907
rect 25605 36873 25639 36907
rect 26065 36873 26099 36907
rect 26801 36873 26835 36907
rect 29285 36873 29319 36907
rect 32965 36873 32999 36907
rect 34989 36873 35023 36907
rect 26433 36805 26467 36839
rect 27721 36805 27755 36839
rect 32137 36805 32171 36839
rect 32353 36805 32387 36839
rect 32597 36805 32631 36839
rect 12449 36737 12483 36771
rect 14657 36737 14691 36771
rect 14749 36737 14783 36771
rect 18337 36737 18371 36771
rect 21097 36737 21131 36771
rect 23581 36737 23615 36771
rect 24041 36737 24075 36771
rect 24869 36737 24903 36771
rect 25697 36737 25731 36771
rect 26157 36737 26191 36771
rect 26250 36737 26284 36771
rect 26525 36737 26559 36771
rect 26622 36737 26656 36771
rect 27077 36737 27111 36771
rect 27261 36737 27295 36771
rect 29469 36737 29503 36771
rect 29745 36737 29779 36771
rect 30389 36737 30423 36771
rect 31033 36737 31067 36771
rect 31953 36737 31987 36771
rect 32781 36737 32815 36771
rect 32873 36737 32907 36771
rect 33241 36737 33275 36771
rect 12725 36669 12759 36703
rect 14381 36669 14415 36703
rect 15025 36669 15059 36703
rect 17141 36669 17175 36703
rect 17325 36669 17359 36703
rect 18613 36669 18647 36703
rect 20269 36669 20303 36703
rect 20545 36669 20579 36703
rect 20821 36669 20855 36703
rect 21005 36669 21039 36703
rect 23305 36669 23339 36703
rect 24133 36669 24167 36703
rect 24317 36669 24351 36703
rect 24593 36669 24627 36703
rect 25513 36669 25547 36703
rect 27445 36669 27479 36703
rect 29561 36669 29595 36703
rect 33517 36669 33551 36703
rect 16681 36601 16715 36635
rect 21465 36601 21499 36635
rect 23673 36601 23707 36635
rect 27261 36601 27295 36635
rect 12081 36533 12115 36567
rect 12909 36533 12943 36567
rect 17969 36533 18003 36567
rect 21833 36533 21867 36567
rect 25237 36533 25271 36567
rect 29193 36533 29227 36567
rect 31493 36533 31527 36567
rect 32321 36533 32355 36567
rect 32505 36533 32539 36567
rect 33149 36533 33183 36567
rect 13185 36329 13219 36363
rect 14197 36329 14231 36363
rect 18981 36329 19015 36363
rect 21741 36329 21775 36363
rect 22293 36329 22327 36363
rect 26157 36329 26191 36363
rect 28549 36329 28583 36363
rect 33517 36329 33551 36363
rect 25053 36261 25087 36295
rect 34713 36261 34747 36295
rect 11713 36193 11747 36227
rect 14841 36193 14875 36227
rect 17233 36193 17267 36227
rect 17509 36193 17543 36227
rect 20269 36193 20303 36227
rect 26801 36193 26835 36227
rect 27077 36193 27111 36227
rect 28917 36193 28951 36227
rect 30113 36193 30147 36227
rect 30297 36193 30331 36227
rect 31033 36193 31067 36227
rect 32597 36193 32631 36227
rect 11437 36125 11471 36159
rect 14565 36125 14599 36159
rect 14657 36125 14691 36159
rect 19993 36125 20027 36159
rect 25329 36125 25363 36159
rect 25881 36125 25915 36159
rect 25973 36125 26007 36159
rect 29285 36125 29319 36159
rect 30757 36125 30791 36159
rect 30941 36125 30975 36159
rect 31585 36125 31619 36159
rect 32045 36125 32079 36159
rect 32229 36125 32263 36159
rect 33241 36125 33275 36159
rect 33333 36125 33367 36159
rect 33517 36125 33551 36159
rect 33609 36125 33643 36159
rect 33885 36125 33919 36159
rect 34897 36125 34931 36159
rect 34989 36125 35023 36159
rect 23581 36057 23615 36091
rect 25605 36057 25639 36091
rect 31401 36057 31435 36091
rect 31953 36057 31987 36091
rect 34713 36057 34747 36091
rect 25513 35989 25547 36023
rect 29653 35989 29687 36023
rect 32229 35989 32263 36023
rect 32781 35989 32815 36023
rect 13001 35785 13035 35819
rect 18705 35785 18739 35819
rect 20913 35785 20947 35819
rect 21281 35785 21315 35819
rect 21373 35785 21407 35819
rect 23673 35785 23707 35819
rect 26341 35785 26375 35819
rect 27245 35785 27279 35819
rect 32137 35785 32171 35819
rect 16129 35717 16163 35751
rect 21833 35717 21867 35751
rect 25145 35717 25179 35751
rect 27445 35717 27479 35751
rect 27537 35717 27571 35751
rect 29653 35717 29687 35751
rect 30113 35717 30147 35751
rect 13093 35649 13127 35683
rect 18613 35649 18647 35683
rect 23581 35649 23615 35683
rect 27997 35649 28031 35683
rect 28181 35649 28215 35683
rect 28917 35649 28951 35683
rect 29561 35649 29595 35683
rect 29745 35649 29779 35683
rect 29837 35649 29871 35683
rect 31677 35649 31711 35683
rect 31861 35649 31895 35683
rect 31953 35649 31987 35683
rect 33333 35649 33367 35683
rect 33425 35649 33459 35683
rect 33609 35649 33643 35683
rect 33701 35649 33735 35683
rect 12909 35581 12943 35615
rect 16221 35581 16255 35615
rect 16405 35581 16439 35615
rect 18889 35581 18923 35615
rect 21465 35581 21499 35615
rect 25421 35581 25455 35615
rect 26801 35581 26835 35615
rect 28273 35581 28307 35615
rect 28641 35581 28675 35615
rect 32597 35581 32631 35615
rect 33241 35581 33275 35615
rect 33977 35581 34011 35615
rect 27077 35513 27111 35547
rect 31677 35513 31711 35547
rect 32229 35513 32263 35547
rect 32781 35513 32815 35547
rect 33609 35513 33643 35547
rect 13461 35445 13495 35479
rect 15761 35445 15795 35479
rect 18245 35445 18279 35479
rect 27261 35445 27295 35479
rect 31585 35445 31619 35479
rect 35449 35445 35483 35479
rect 11897 35241 11931 35275
rect 16957 35241 16991 35275
rect 19073 35241 19107 35275
rect 26157 35241 26191 35275
rect 26249 35241 26283 35275
rect 31493 35241 31527 35275
rect 35817 35241 35851 35275
rect 31309 35173 31343 35207
rect 34345 35173 34379 35207
rect 13645 35105 13679 35139
rect 15209 35105 15243 35139
rect 17325 35105 17359 35139
rect 17601 35105 17635 35139
rect 19717 35105 19751 35139
rect 19809 35105 19843 35139
rect 27997 35105 28031 35139
rect 29561 35105 29595 35139
rect 31769 35105 31803 35139
rect 31953 35105 31987 35139
rect 32505 35105 32539 35139
rect 32597 35105 32631 35139
rect 33517 35105 33551 35139
rect 33885 35105 33919 35139
rect 24409 35037 24443 35071
rect 28089 35037 28123 35071
rect 28549 35037 28583 35071
rect 28733 35037 28767 35071
rect 28825 35037 28859 35071
rect 29929 35037 29963 35071
rect 30205 35037 30239 35071
rect 30849 35037 30883 35071
rect 31677 35037 31711 35071
rect 31861 35037 31895 35071
rect 32229 35037 32263 35071
rect 33149 35037 33183 35071
rect 33333 35037 33367 35071
rect 33609 35037 33643 35071
rect 33701 35037 33735 35071
rect 34805 35037 34839 35071
rect 35541 35037 35575 35071
rect 35633 35037 35667 35071
rect 36093 35037 36127 35071
rect 13369 34969 13403 35003
rect 15485 34969 15519 35003
rect 24685 34969 24719 35003
rect 27721 34969 27755 35003
rect 29837 34969 29871 35003
rect 35173 34969 35207 35003
rect 35817 34969 35851 35003
rect 19257 34901 19291 34935
rect 19625 34901 19659 34935
rect 29745 34901 29779 34935
rect 30113 34901 30147 34935
rect 30665 34901 30699 34935
rect 35909 34901 35943 34935
rect 12357 34697 12391 34731
rect 15945 34697 15979 34731
rect 20545 34697 20579 34731
rect 25421 34697 25455 34731
rect 27905 34697 27939 34731
rect 28457 34697 28491 34731
rect 28549 34697 28583 34731
rect 32413 34697 32447 34731
rect 32597 34697 32631 34731
rect 33333 34697 33367 34731
rect 33609 34697 33643 34731
rect 12265 34629 12299 34663
rect 13185 34629 13219 34663
rect 27537 34629 27571 34663
rect 27753 34629 27787 34663
rect 33057 34629 33091 34663
rect 13093 34561 13127 34595
rect 14197 34561 14231 34595
rect 17141 34561 17175 34595
rect 17325 34561 17359 34595
rect 17417 34561 17451 34595
rect 18797 34561 18831 34595
rect 20637 34561 20671 34595
rect 22477 34561 22511 34595
rect 25513 34561 25547 34595
rect 27997 34561 28031 34595
rect 29377 34561 29411 34595
rect 29561 34561 29595 34595
rect 30481 34561 30515 34595
rect 30941 34561 30975 34595
rect 31585 34561 31619 34595
rect 31953 34561 31987 34595
rect 32321 34561 32355 34595
rect 32689 34561 32723 34595
rect 33241 34561 33275 34595
rect 33425 34561 33459 34595
rect 33701 34561 33735 34595
rect 33977 34561 34011 34595
rect 12541 34493 12575 34527
rect 13369 34493 13403 34527
rect 16681 34493 16715 34527
rect 19073 34493 19107 34527
rect 22569 34493 22603 34527
rect 22753 34493 22787 34527
rect 25697 34493 25731 34527
rect 28181 34493 28215 34527
rect 28273 34493 28307 34527
rect 28641 34493 28675 34527
rect 29101 34493 29135 34527
rect 29837 34493 29871 34527
rect 32781 34493 32815 34527
rect 33793 34493 33827 34527
rect 34253 34493 34287 34527
rect 35725 34493 35759 34527
rect 11897 34357 11931 34391
rect 12725 34357 12759 34391
rect 14460 34357 14494 34391
rect 22109 34357 22143 34391
rect 25053 34357 25087 34391
rect 27721 34357 27755 34391
rect 30573 34357 30607 34391
rect 32965 34357 32999 34391
rect 13553 34153 13587 34187
rect 17601 34153 17635 34187
rect 23305 34153 23339 34187
rect 28457 34153 28491 34187
rect 29101 34153 29135 34187
rect 33241 34153 33275 34187
rect 11805 34017 11839 34051
rect 12081 34017 12115 34051
rect 14749 34017 14783 34051
rect 19349 34017 19383 34051
rect 24685 34017 24719 34051
rect 26709 34017 26743 34051
rect 26985 34017 27019 34051
rect 29837 34017 29871 34051
rect 31493 34017 31527 34051
rect 35265 34017 35299 34051
rect 15669 33949 15703 33983
rect 18153 33949 18187 33983
rect 21557 33949 21591 33983
rect 24409 33949 24443 33983
rect 29285 33949 29319 33983
rect 29377 33949 29411 33983
rect 29561 33949 29595 33983
rect 31125 33949 31159 33983
rect 33517 33949 33551 33983
rect 34345 33949 34379 33983
rect 35633 33949 35667 33983
rect 35725 33949 35759 33983
rect 35909 33949 35943 33983
rect 15577 33881 15611 33915
rect 15945 33881 15979 33915
rect 17877 33881 17911 33915
rect 19625 33881 19659 33915
rect 21833 33881 21867 33915
rect 30573 33881 30607 33915
rect 31776 33881 31810 33915
rect 35817 33881 35851 33915
rect 17417 33813 17451 33847
rect 18061 33813 18095 33847
rect 21097 33813 21131 33847
rect 26157 33813 26191 33847
rect 34805 33813 34839 33847
rect 35449 33813 35483 33847
rect 13277 33609 13311 33643
rect 15761 33609 15795 33643
rect 16681 33609 16715 33643
rect 17049 33609 17083 33643
rect 19717 33609 19751 33643
rect 20177 33609 20211 33643
rect 22201 33609 22235 33643
rect 26341 33609 26375 33643
rect 33793 33609 33827 33643
rect 34437 33609 34471 33643
rect 11805 33541 11839 33575
rect 14289 33541 14323 33575
rect 20545 33541 20579 33575
rect 21373 33541 21407 33575
rect 32137 33541 32171 33575
rect 32873 33541 32907 33575
rect 34589 33541 34623 33575
rect 34805 33541 34839 33575
rect 11529 33473 11563 33507
rect 17141 33473 17175 33507
rect 17877 33473 17911 33507
rect 20085 33473 20119 33507
rect 22661 33473 22695 33507
rect 24593 33473 24627 33507
rect 27905 33473 27939 33507
rect 28181 33473 28215 33507
rect 28273 33473 28307 33507
rect 28733 33473 28767 33507
rect 28917 33473 28951 33507
rect 29377 33473 29411 33507
rect 29653 33473 29687 33507
rect 29837 33473 29871 33507
rect 31677 33473 31711 33507
rect 33241 33473 33275 33507
rect 34253 33473 34287 33507
rect 35081 33473 35115 33507
rect 14013 33405 14047 33439
rect 17325 33405 17359 33439
rect 17693 33405 17727 33439
rect 17785 33405 17819 33439
rect 20269 33405 20303 33439
rect 22293 33405 22327 33439
rect 22385 33405 22419 33439
rect 22937 33405 22971 33439
rect 24869 33405 24903 33439
rect 27077 33405 27111 33439
rect 29009 33405 29043 33439
rect 30113 33405 30147 33439
rect 31585 33405 31619 33439
rect 33977 33405 34011 33439
rect 34069 33405 34103 33439
rect 34161 33405 34195 33439
rect 35265 33405 35299 33439
rect 29469 33337 29503 33371
rect 34897 33337 34931 33371
rect 18245 33269 18279 33303
rect 21833 33269 21867 33303
rect 24409 33269 24443 33303
rect 28089 33269 28123 33303
rect 31861 33269 31895 33303
rect 34621 33269 34655 33303
rect 17049 33065 17083 33099
rect 22569 33065 22603 33099
rect 23121 33065 23155 33099
rect 25237 33065 25271 33099
rect 28549 33065 28583 33099
rect 28733 33065 28767 33099
rect 30113 33065 30147 33099
rect 30297 33065 30331 33099
rect 34345 33065 34379 33099
rect 13185 32929 13219 32963
rect 13369 32929 13403 32963
rect 18521 32929 18555 32963
rect 19717 32929 19751 32963
rect 19809 32929 19843 32963
rect 21097 32929 21131 32963
rect 23765 32929 23799 32963
rect 25789 32929 25823 32963
rect 29009 32929 29043 32963
rect 30573 32929 30607 32963
rect 30665 32929 30699 32963
rect 30757 32929 30791 32963
rect 14841 32861 14875 32895
rect 18797 32861 18831 32895
rect 20177 32861 20211 32895
rect 20821 32861 20855 32895
rect 23489 32861 23523 32895
rect 26065 32861 26099 32895
rect 29193 32861 29227 32895
rect 29377 32861 29411 32895
rect 30205 32861 30239 32895
rect 30481 32861 30515 32895
rect 31125 32861 31159 32895
rect 32413 32861 32447 32895
rect 33885 32861 33919 32895
rect 34161 32861 34195 32895
rect 19625 32793 19659 32827
rect 25605 32793 25639 32827
rect 28717 32793 28751 32827
rect 28917 32793 28951 32827
rect 31401 32793 31435 32827
rect 32137 32793 32171 32827
rect 33333 32793 33367 32827
rect 12725 32725 12759 32759
rect 13093 32725 13127 32759
rect 19257 32725 19291 32759
rect 23581 32725 23615 32759
rect 25697 32725 25731 32759
rect 31033 32725 31067 32759
rect 33977 32725 34011 32759
rect 18061 32521 18095 32555
rect 22201 32521 22235 32555
rect 28917 32521 28951 32555
rect 35265 32521 35299 32555
rect 14841 32453 14875 32487
rect 19533 32453 19567 32487
rect 20361 32453 20395 32487
rect 25881 32453 25915 32487
rect 30173 32453 30207 32487
rect 30389 32453 30423 32487
rect 31125 32453 31159 32487
rect 17049 32385 17083 32419
rect 25789 32385 25823 32419
rect 26617 32385 26651 32419
rect 27169 32385 27203 32419
rect 29745 32385 29779 32419
rect 29929 32385 29963 32419
rect 30757 32385 30791 32419
rect 31861 32385 31895 32419
rect 32597 32385 32631 32419
rect 32965 32385 32999 32419
rect 34989 32385 35023 32419
rect 35173 32385 35207 32419
rect 35449 32385 35483 32419
rect 12909 32317 12943 32351
rect 13185 32317 13219 32351
rect 15577 32317 15611 32351
rect 17141 32317 17175 32351
rect 17325 32317 17359 32351
rect 19809 32317 19843 32351
rect 21097 32317 21131 32351
rect 22293 32317 22327 32351
rect 22477 32317 22511 32351
rect 27445 32317 27479 32351
rect 30481 32317 30515 32351
rect 33149 32317 33183 32351
rect 33425 32317 33459 32351
rect 30665 32249 30699 32283
rect 31309 32249 31343 32283
rect 35081 32249 35115 32283
rect 14657 32181 14691 32215
rect 16681 32181 16715 32215
rect 21833 32181 21867 32215
rect 29929 32181 29963 32215
rect 30021 32181 30055 32215
rect 30205 32181 30239 32215
rect 30573 32181 30607 32215
rect 34897 32181 34931 32215
rect 13553 31977 13587 32011
rect 17049 31977 17083 32011
rect 22477 31977 22511 32011
rect 27445 31909 27479 31943
rect 34345 31909 34379 31943
rect 12081 31841 12115 31875
rect 14933 31841 14967 31875
rect 15025 31841 15059 31875
rect 15577 31841 15611 31875
rect 20729 31841 20763 31875
rect 21005 31841 21039 31875
rect 23581 31841 23615 31875
rect 23765 31841 23799 31875
rect 24961 31841 24995 31875
rect 25605 31841 25639 31875
rect 27077 31841 27111 31875
rect 27353 31841 27387 31875
rect 27997 31841 28031 31875
rect 30757 31841 30791 31875
rect 32597 31841 32631 31875
rect 35449 31841 35483 31875
rect 11805 31773 11839 31807
rect 15301 31773 15335 31807
rect 28917 31773 28951 31807
rect 29193 31773 29227 31807
rect 29377 31773 29411 31807
rect 29929 31773 29963 31807
rect 30113 31773 30147 31807
rect 30481 31773 30515 31807
rect 32505 31773 32539 31807
rect 34713 31773 34747 31807
rect 23489 31705 23523 31739
rect 24777 31705 24811 31739
rect 27813 31705 27847 31739
rect 32873 31705 32907 31739
rect 14473 31637 14507 31671
rect 14841 31637 14875 31671
rect 23121 31637 23155 31671
rect 24409 31637 24443 31671
rect 24869 31637 24903 31671
rect 27905 31637 27939 31671
rect 29837 31637 29871 31671
rect 13369 31433 13403 31467
rect 13829 31433 13863 31467
rect 15945 31433 15979 31467
rect 17233 31433 17267 31467
rect 21649 31433 21683 31467
rect 23949 31433 23983 31467
rect 25789 31433 25823 31467
rect 26341 31433 26375 31467
rect 28825 31433 28859 31467
rect 31861 31433 31895 31467
rect 13737 31365 13771 31399
rect 14473 31365 14507 31399
rect 22477 31365 22511 31399
rect 24317 31365 24351 31399
rect 30297 31365 30331 31399
rect 33885 31365 33919 31399
rect 9965 31297 9999 31331
rect 14197 31297 14231 31331
rect 17141 31297 17175 31331
rect 18061 31297 18095 31331
rect 26249 31297 26283 31331
rect 30573 31297 30607 31331
rect 31953 31297 31987 31331
rect 32413 31297 32447 31331
rect 34345 31297 34379 31331
rect 34529 31297 34563 31331
rect 34621 31297 34655 31331
rect 8125 31229 8159 31263
rect 8401 31229 8435 31263
rect 13921 31229 13955 31263
rect 17417 31229 17451 31263
rect 18337 31229 18371 31263
rect 19901 31229 19935 31263
rect 20177 31229 20211 31263
rect 22201 31229 22235 31263
rect 24041 31229 24075 31263
rect 26525 31229 26559 31263
rect 26985 31229 27019 31263
rect 27261 31229 27295 31263
rect 33149 31229 33183 31263
rect 9873 31093 9907 31127
rect 10057 31093 10091 31127
rect 16773 31093 16807 31127
rect 19809 31093 19843 31127
rect 25881 31093 25915 31127
rect 28733 31093 28767 31127
rect 8953 30889 8987 30923
rect 19257 30889 19291 30923
rect 20361 30889 20395 30923
rect 26157 30889 26191 30923
rect 26985 30889 27019 30923
rect 29824 30889 29858 30923
rect 31309 30889 31343 30923
rect 6653 30753 6687 30787
rect 6745 30753 6779 30787
rect 9505 30753 9539 30787
rect 13461 30753 13495 30787
rect 15485 30753 15519 30787
rect 17325 30753 17359 30787
rect 19073 30753 19107 30787
rect 19717 30753 19751 30787
rect 19901 30753 19935 30787
rect 20913 30753 20947 30787
rect 24685 30753 24719 30787
rect 27537 30753 27571 30787
rect 29561 30753 29595 30787
rect 32045 30753 32079 30787
rect 34989 30753 35023 30787
rect 3893 30685 3927 30719
rect 4077 30685 4111 30719
rect 9781 30685 9815 30719
rect 9965 30685 9999 30719
rect 19625 30685 19659 30719
rect 20821 30685 20855 30719
rect 24409 30685 24443 30719
rect 27353 30685 27387 30719
rect 31861 30685 31895 30719
rect 32597 30685 32631 30719
rect 33609 30685 33643 30719
rect 35081 30685 35115 30719
rect 35265 30685 35299 30719
rect 6377 30617 6411 30651
rect 7021 30617 7055 30651
rect 9321 30617 9355 30651
rect 9873 30617 9907 30651
rect 15761 30617 15795 30651
rect 17601 30617 17635 30651
rect 20729 30617 20763 30651
rect 31769 30617 31803 30651
rect 35725 30617 35759 30651
rect 3985 30549 4019 30583
rect 4905 30549 4939 30583
rect 8493 30549 8527 30583
rect 9413 30549 9447 30583
rect 12817 30549 12851 30583
rect 13185 30549 13219 30583
rect 13277 30549 13311 30583
rect 17233 30549 17267 30583
rect 27445 30549 27479 30583
rect 31401 30549 31435 30583
rect 6377 30345 6411 30379
rect 8585 30345 8619 30379
rect 9229 30345 9263 30379
rect 17877 30345 17911 30379
rect 18245 30345 18279 30379
rect 18337 30345 18371 30379
rect 26341 30345 26375 30379
rect 32413 30345 32447 30379
rect 8309 30277 8343 30311
rect 8753 30277 8787 30311
rect 8953 30277 8987 30311
rect 9321 30277 9355 30311
rect 25789 30277 25823 30311
rect 33885 30277 33919 30311
rect 1777 30209 1811 30243
rect 3341 30209 3375 30243
rect 5641 30209 5675 30243
rect 5825 30209 5859 30243
rect 6745 30209 6779 30243
rect 8033 30209 8067 30243
rect 8125 30209 8159 30243
rect 9413 30209 9447 30243
rect 10425 30209 10459 30243
rect 11621 30209 11655 30243
rect 15485 30209 15519 30243
rect 23949 30209 23983 30243
rect 26249 30209 26283 30243
rect 30205 30209 30239 30243
rect 34161 30209 34195 30243
rect 3433 30141 3467 30175
rect 3709 30141 3743 30175
rect 5733 30141 5767 30175
rect 6837 30141 6871 30175
rect 6929 30141 6963 30175
rect 10517 30141 10551 30175
rect 10609 30141 10643 30175
rect 11897 30141 11931 30175
rect 15209 30141 15243 30175
rect 18429 30141 18463 30175
rect 23673 30141 23707 30175
rect 26525 30141 26559 30175
rect 30481 30141 30515 30175
rect 8309 30073 8343 30107
rect 9045 30073 9079 30107
rect 9597 30073 9631 30107
rect 24501 30073 24535 30107
rect 5181 30005 5215 30039
rect 8769 30005 8803 30039
rect 10057 30005 10091 30039
rect 13369 30005 13403 30039
rect 13737 30005 13771 30039
rect 22201 30005 22235 30039
rect 25881 30005 25915 30039
rect 31953 30005 31987 30039
rect 3801 29801 3835 29835
rect 7849 29801 7883 29835
rect 8125 29801 8159 29835
rect 15301 29801 15335 29835
rect 27629 29801 27663 29835
rect 4629 29733 4663 29767
rect 27721 29733 27755 29767
rect 2145 29665 2179 29699
rect 4445 29665 4479 29699
rect 5181 29665 5215 29699
rect 9689 29665 9723 29699
rect 9965 29665 9999 29699
rect 14657 29665 14691 29699
rect 17509 29665 17543 29699
rect 25053 29665 25087 29699
rect 25145 29665 25179 29699
rect 25881 29665 25915 29699
rect 26157 29665 26191 29699
rect 28365 29665 28399 29699
rect 30205 29665 30239 29699
rect 31033 29665 31067 29699
rect 33425 29665 33459 29699
rect 1869 29597 1903 29631
rect 4169 29597 4203 29631
rect 4813 29597 4847 29631
rect 4905 29597 4939 29631
rect 7757 29597 7791 29631
rect 7941 29597 7975 29631
rect 8033 29597 8067 29631
rect 8217 29597 8251 29631
rect 8309 29597 8343 29631
rect 8493 29597 8527 29631
rect 8677 29597 8711 29631
rect 11529 29597 11563 29631
rect 14933 29597 14967 29631
rect 19257 29597 19291 29631
rect 21189 29597 21223 29631
rect 21373 29597 21407 29631
rect 23581 29597 23615 29631
rect 28089 29597 28123 29631
rect 32229 29597 32263 29631
rect 33241 29597 33275 29631
rect 5457 29529 5491 29563
rect 11805 29529 11839 29563
rect 17233 29529 17267 29563
rect 19533 29529 19567 29563
rect 23305 29529 23339 29563
rect 3617 29461 3651 29495
rect 4261 29461 4295 29495
rect 6929 29461 6963 29495
rect 9321 29461 9355 29495
rect 9505 29461 9539 29495
rect 11437 29461 11471 29495
rect 13277 29461 13311 29495
rect 14841 29461 14875 29495
rect 15761 29461 15795 29495
rect 21005 29461 21039 29495
rect 21833 29461 21867 29495
rect 24593 29461 24627 29495
rect 24961 29461 24995 29495
rect 28181 29461 28215 29495
rect 29561 29461 29595 29495
rect 29929 29461 29963 29495
rect 30021 29461 30055 29495
rect 32873 29461 32907 29495
rect 33333 29461 33367 29495
rect 3157 29257 3191 29291
rect 4261 29257 4295 29291
rect 5457 29257 5491 29291
rect 5549 29257 5583 29291
rect 7113 29257 7147 29291
rect 7297 29257 7331 29291
rect 10517 29257 10551 29291
rect 12541 29257 12575 29291
rect 12909 29257 12943 29291
rect 15669 29257 15703 29291
rect 17417 29257 17451 29291
rect 19717 29257 19751 29291
rect 20085 29257 20119 29291
rect 23305 29257 23339 29291
rect 23673 29257 23707 29291
rect 28825 29257 28859 29291
rect 33977 29257 34011 29291
rect 3893 29189 3927 29223
rect 4093 29189 4127 29223
rect 5089 29189 5123 29223
rect 5305 29189 5339 29223
rect 9597 29189 9631 29223
rect 10793 29189 10827 29223
rect 13001 29189 13035 29223
rect 23581 29189 23615 29223
rect 25145 29189 25179 29223
rect 32505 29189 32539 29223
rect 5733 29121 5767 29155
rect 6009 29121 6043 29155
rect 9873 29121 9907 29155
rect 10609 29121 10643 29155
rect 10701 29121 10735 29155
rect 10885 29121 10919 29155
rect 17049 29121 17083 29155
rect 18889 29121 18923 29155
rect 18981 29121 19015 29155
rect 20177 29121 20211 29155
rect 21281 29121 21315 29155
rect 21373 29121 21407 29155
rect 25421 29121 25455 29155
rect 26985 29121 27019 29155
rect 31309 29121 31343 29155
rect 31493 29121 31527 29155
rect 1409 29053 1443 29087
rect 1685 29053 1719 29087
rect 7481 29053 7515 29087
rect 7757 29053 7791 29087
rect 9689 29053 9723 29087
rect 13185 29053 13219 29087
rect 13921 29053 13955 29087
rect 14197 29053 14231 29087
rect 16773 29053 16807 29087
rect 16957 29053 16991 29087
rect 19165 29053 19199 29087
rect 20269 29053 20303 29087
rect 21465 29053 21499 29087
rect 27261 29053 27295 29087
rect 30481 29053 30515 29087
rect 30757 29053 30791 29087
rect 30849 29053 30883 29087
rect 31585 29053 31619 29087
rect 32229 29053 32263 29087
rect 9229 28985 9263 29019
rect 10057 28985 10091 29019
rect 4077 28917 4111 28951
rect 5273 28917 5307 28951
rect 5917 28917 5951 28951
rect 9597 28917 9631 28951
rect 18521 28917 18555 28951
rect 20913 28917 20947 28951
rect 28733 28917 28767 28951
rect 29009 28917 29043 28951
rect 2053 28713 2087 28747
rect 4629 28713 4663 28747
rect 6009 28713 6043 28747
rect 7941 28713 7975 28747
rect 8309 28713 8343 28747
rect 14841 28713 14875 28747
rect 17325 28713 17359 28747
rect 22201 28713 22235 28747
rect 23029 28713 23063 28747
rect 23857 28713 23891 28747
rect 27261 28713 27295 28747
rect 29377 28713 29411 28747
rect 4353 28645 4387 28679
rect 30113 28645 30147 28679
rect 2697 28577 2731 28611
rect 3893 28577 3927 28611
rect 3985 28577 4019 28611
rect 13185 28577 13219 28611
rect 15485 28577 15519 28611
rect 18797 28577 18831 28611
rect 19073 28577 19107 28611
rect 20085 28577 20119 28611
rect 20729 28577 20763 28611
rect 22385 28577 22419 28611
rect 22569 28577 22603 28611
rect 23305 28577 23339 28611
rect 25881 28577 25915 28611
rect 26157 28577 26191 28611
rect 27905 28577 27939 28611
rect 28825 28577 28859 28611
rect 28917 28577 28951 28611
rect 31585 28577 31619 28611
rect 33425 28577 33459 28611
rect 2421 28509 2455 28543
rect 2881 28509 2915 28543
rect 3065 28509 3099 28543
rect 4077 28509 4111 28543
rect 4169 28509 4203 28543
rect 8125 28509 8159 28543
rect 8401 28509 8435 28543
rect 13093 28509 13127 28543
rect 15209 28509 15243 28543
rect 20453 28509 20487 28543
rect 22661 28509 22695 28543
rect 23397 28509 23431 28543
rect 27629 28509 27663 28543
rect 27721 28509 27755 28543
rect 29009 28509 29043 28543
rect 31861 28509 31895 28543
rect 33149 28509 33183 28543
rect 33333 28509 33367 28543
rect 4445 28441 4479 28475
rect 5977 28441 6011 28475
rect 6193 28441 6227 28475
rect 15301 28441 15335 28475
rect 19901 28441 19935 28475
rect 19993 28441 20027 28475
rect 32689 28441 32723 28475
rect 2513 28373 2547 28407
rect 2973 28373 3007 28407
rect 4645 28373 4679 28407
rect 4813 28373 4847 28407
rect 5825 28373 5859 28407
rect 12633 28373 12667 28407
rect 13001 28373 13035 28407
rect 19533 28373 19567 28407
rect 23489 28373 23523 28407
rect 24409 28373 24443 28407
rect 3065 28169 3099 28203
rect 5641 28169 5675 28203
rect 16497 28169 16531 28203
rect 28181 28169 28215 28203
rect 33885 28169 33919 28203
rect 3217 28101 3251 28135
rect 3433 28101 3467 28135
rect 5273 28101 5307 28135
rect 5473 28101 5507 28135
rect 5733 28101 5767 28135
rect 11989 28101 12023 28135
rect 29653 28101 29687 28135
rect 32413 28101 32447 28135
rect 2237 28033 2271 28067
rect 2697 28033 2731 28067
rect 2881 28033 2915 28067
rect 2973 28033 3007 28067
rect 3893 28033 3927 28067
rect 3985 28033 4019 28067
rect 4169 28033 4203 28067
rect 6009 28033 6043 28067
rect 6561 28033 6595 28067
rect 6745 28033 6779 28067
rect 10793 28033 10827 28067
rect 11713 28033 11747 28067
rect 21373 28033 21407 28067
rect 26065 28033 26099 28067
rect 30481 28033 30515 28067
rect 30941 28033 30975 28067
rect 2421 27965 2455 27999
rect 2513 27965 2547 27999
rect 5917 27965 5951 27999
rect 6653 27965 6687 27999
rect 6837 27965 6871 27999
rect 8769 27965 8803 27999
rect 9045 27965 9079 27999
rect 10977 27965 11011 27999
rect 14749 27965 14783 27999
rect 15025 27965 15059 27999
rect 18153 27965 18187 27999
rect 18429 27965 18463 27999
rect 19625 27965 19659 27999
rect 26157 27965 26191 27999
rect 26249 27965 26283 27999
rect 29929 27965 29963 27999
rect 30297 27965 30331 27999
rect 30389 27965 30423 27999
rect 31677 27965 31711 27999
rect 32137 27965 32171 27999
rect 4353 27897 4387 27931
rect 6377 27897 6411 27931
rect 10609 27897 10643 27931
rect 2053 27829 2087 27863
rect 3249 27829 3283 27863
rect 5457 27829 5491 27863
rect 5917 27829 5951 27863
rect 6193 27829 6227 27863
rect 10517 27829 10551 27863
rect 13461 27829 13495 27863
rect 16681 27829 16715 27863
rect 25697 27829 25731 27863
rect 30849 27829 30883 27863
rect 2132 27625 2166 27659
rect 3617 27625 3651 27659
rect 4169 27625 4203 27659
rect 6377 27625 6411 27659
rect 9505 27625 9539 27659
rect 18245 27625 18279 27659
rect 19520 27625 19554 27659
rect 31051 27625 31085 27659
rect 32492 27625 32526 27659
rect 33977 27625 34011 27659
rect 5273 27557 5307 27591
rect 12081 27557 12115 27591
rect 16313 27557 16347 27591
rect 21005 27557 21039 27591
rect 3801 27489 3835 27523
rect 7849 27489 7883 27523
rect 8125 27489 8159 27523
rect 12173 27489 12207 27523
rect 16773 27489 16807 27523
rect 16865 27489 16899 27523
rect 17693 27489 17727 27523
rect 19257 27489 19291 27523
rect 21189 27489 21223 27523
rect 22661 27489 22695 27523
rect 23581 27489 23615 27523
rect 23765 27489 23799 27523
rect 24869 27489 24903 27523
rect 27629 27489 27663 27523
rect 28917 27489 28951 27523
rect 1869 27421 1903 27455
rect 3985 27421 4019 27455
rect 5457 27421 5491 27455
rect 5641 27421 5675 27455
rect 6285 27421 6319 27455
rect 9229 27421 9263 27455
rect 9413 27421 9447 27455
rect 9689 27421 9723 27455
rect 9965 27421 9999 27455
rect 10149 27421 10183 27455
rect 10333 27421 10367 27455
rect 15853 27421 15887 27455
rect 17877 27421 17911 27455
rect 22017 27421 22051 27455
rect 27813 27421 27847 27455
rect 31309 27421 31343 27455
rect 32229 27421 32263 27455
rect 10609 27353 10643 27387
rect 12449 27353 12483 27387
rect 15577 27353 15611 27387
rect 16681 27353 16715 27387
rect 17785 27353 17819 27387
rect 22569 27353 22603 27387
rect 23857 27353 23891 27387
rect 25145 27353 25179 27387
rect 28641 27353 28675 27387
rect 5549 27285 5583 27319
rect 5825 27285 5859 27319
rect 6193 27285 6227 27319
rect 9413 27285 9447 27319
rect 13921 27285 13955 27319
rect 14105 27285 14139 27319
rect 22109 27285 22143 27319
rect 22477 27285 22511 27319
rect 24225 27285 24259 27319
rect 26617 27285 26651 27319
rect 27721 27285 27755 27319
rect 28181 27285 28215 27319
rect 28273 27285 28307 27319
rect 28733 27285 28767 27319
rect 29561 27285 29595 27319
rect 5565 27081 5599 27115
rect 6035 27081 6069 27115
rect 8585 27081 8619 27115
rect 10425 27081 10459 27115
rect 11069 27081 11103 27115
rect 13369 27081 13403 27115
rect 13829 27081 13863 27115
rect 18705 27081 18739 27115
rect 33241 27081 33275 27115
rect 33609 27081 33643 27115
rect 5365 27013 5399 27047
rect 5825 27013 5859 27047
rect 6745 27013 6779 27047
rect 6929 27013 6963 27047
rect 7145 27013 7179 27047
rect 7757 27013 7791 27047
rect 8769 27013 8803 27047
rect 9965 27013 9999 27047
rect 10165 27013 10199 27047
rect 10577 27013 10611 27047
rect 10793 27013 10827 27047
rect 14105 27013 14139 27047
rect 25329 27013 25363 27047
rect 26433 27013 26467 27047
rect 28457 27013 28491 27047
rect 30665 27013 30699 27047
rect 32137 27013 32171 27047
rect 6515 26979 6549 27013
rect 4905 26945 4939 26979
rect 7573 26945 7607 26979
rect 7665 26945 7699 26979
rect 8401 26945 8435 26979
rect 8493 26945 8527 26979
rect 10885 26945 10919 26979
rect 11161 26945 11195 26979
rect 13461 26945 13495 26979
rect 14841 26945 14875 26979
rect 15853 26945 15887 26979
rect 16405 26945 16439 26979
rect 17693 26945 17727 26979
rect 19257 26945 19291 26979
rect 19901 26945 19935 26979
rect 25605 26945 25639 26979
rect 25697 26945 25731 26979
rect 31033 26945 31067 26979
rect 32597 26945 32631 26979
rect 32781 26945 32815 26979
rect 32873 26945 32907 26979
rect 1409 26877 1443 26911
rect 1685 26877 1719 26911
rect 5181 26877 5215 26911
rect 13277 26877 13311 26911
rect 15025 26877 15059 26911
rect 17785 26877 17819 26911
rect 17877 26877 17911 26911
rect 18797 26877 18831 26911
rect 18889 26877 18923 26911
rect 20177 26877 20211 26911
rect 23489 26877 23523 26911
rect 23765 26877 23799 26911
rect 26985 26877 27019 26911
rect 28733 26877 28767 26911
rect 29193 26877 29227 26911
rect 30941 26877 30975 26911
rect 33701 26877 33735 26911
rect 33885 26877 33919 26911
rect 5089 26809 5123 26843
rect 6377 26809 6411 26843
rect 7297 26809 7331 26843
rect 7389 26809 7423 26843
rect 8217 26809 8251 26843
rect 10333 26809 10367 26843
rect 10885 26809 10919 26843
rect 3157 26741 3191 26775
rect 4721 26741 4755 26775
rect 5549 26741 5583 26775
rect 5733 26741 5767 26775
rect 6009 26741 6043 26775
rect 6193 26741 6227 26775
rect 6561 26741 6595 26775
rect 7113 26741 7147 26775
rect 7941 26741 7975 26775
rect 10149 26741 10183 26775
rect 10609 26741 10643 26775
rect 17325 26741 17359 26775
rect 18337 26741 18371 26775
rect 21649 26741 21683 26775
rect 22017 26741 22051 26775
rect 23857 26741 23891 26775
rect 1961 26537 1995 26571
rect 4432 26537 4466 26571
rect 5917 26537 5951 26571
rect 6377 26537 6411 26571
rect 8309 26537 8343 26571
rect 9505 26537 9539 26571
rect 10057 26537 10091 26571
rect 13001 26537 13035 26571
rect 18889 26537 18923 26571
rect 22845 26537 22879 26571
rect 24409 26537 24443 26571
rect 26985 26537 27019 26571
rect 31493 26537 31527 26571
rect 9229 26469 9263 26503
rect 21833 26469 21867 26503
rect 2605 26401 2639 26435
rect 4169 26401 4203 26435
rect 6469 26401 6503 26435
rect 9321 26401 9355 26435
rect 13461 26401 13495 26435
rect 13645 26401 13679 26435
rect 14565 26401 14599 26435
rect 14749 26401 14783 26435
rect 17141 26401 17175 26435
rect 19993 26401 20027 26435
rect 20269 26401 20303 26435
rect 21741 26401 21775 26435
rect 22293 26401 22327 26435
rect 22477 26401 22511 26435
rect 23305 26401 23339 26435
rect 23397 26401 23431 26435
rect 25881 26401 25915 26435
rect 26157 26401 26191 26435
rect 28457 26401 28491 26435
rect 28733 26401 28767 26435
rect 29745 26401 29779 26435
rect 33609 26401 33643 26435
rect 6653 26333 6687 26367
rect 8953 26333 8987 26367
rect 9045 26333 9079 26367
rect 9597 26333 9631 26367
rect 9965 26333 9999 26367
rect 10149 26333 10183 26367
rect 10333 26333 10367 26367
rect 13369 26333 13403 26367
rect 14933 26333 14967 26367
rect 22201 26333 22235 26367
rect 23213 26333 23247 26367
rect 31585 26333 31619 26367
rect 33333 26333 33367 26367
rect 2329 26265 2363 26299
rect 6377 26265 6411 26299
rect 7021 26265 7055 26299
rect 9229 26265 9263 26299
rect 9321 26265 9355 26299
rect 10609 26265 10643 26299
rect 17417 26265 17451 26299
rect 26709 26265 26743 26299
rect 30021 26265 30055 26299
rect 32321 26265 32355 26299
rect 2421 26197 2455 26231
rect 6837 26197 6871 26231
rect 12081 26197 12115 26231
rect 14105 26197 14139 26231
rect 14473 26197 14507 26231
rect 32965 26197 32999 26231
rect 33425 26197 33459 26231
rect 3709 25993 3743 26027
rect 4721 25993 4755 26027
rect 9689 25993 9723 26027
rect 10977 25993 11011 26027
rect 14565 25993 14599 26027
rect 17049 25993 17083 26027
rect 17417 25993 17451 26027
rect 33885 25993 33919 26027
rect 3525 25925 3559 25959
rect 6193 25925 6227 25959
rect 10885 25925 10919 25959
rect 17969 25925 18003 25959
rect 24409 25925 24443 25959
rect 25789 25925 25823 25959
rect 30113 25925 30147 25959
rect 32413 25925 32447 25959
rect 3341 25857 3375 25891
rect 4261 25857 4295 25891
rect 6561 25857 6595 25891
rect 7297 25857 7331 25891
rect 7941 25857 7975 25891
rect 10149 25857 10183 25891
rect 10609 25857 10643 25891
rect 11161 25857 11195 25891
rect 12817 25857 12851 25891
rect 21465 25857 21499 25891
rect 25329 25857 25363 25891
rect 25421 25857 25455 25891
rect 28089 25857 28123 25891
rect 28273 25857 28307 25891
rect 29377 25857 29411 25891
rect 29469 25857 29503 25891
rect 29653 25857 29687 25891
rect 6653 25789 6687 25823
rect 6745 25789 6779 25823
rect 6837 25789 6871 25823
rect 8217 25789 8251 25823
rect 9965 25789 9999 25823
rect 10057 25789 10091 25823
rect 10241 25789 10275 25823
rect 10793 25789 10827 25823
rect 11345 25789 11379 25823
rect 13093 25789 13127 25823
rect 16865 25789 16899 25823
rect 16957 25789 16991 25823
rect 17693 25789 17727 25823
rect 25513 25789 25547 25823
rect 26525 25789 26559 25823
rect 27629 25789 27663 25823
rect 28365 25789 28399 25823
rect 30205 25789 30239 25823
rect 30481 25789 30515 25823
rect 32137 25789 32171 25823
rect 9781 25721 9815 25755
rect 24961 25721 24995 25755
rect 6377 25653 6411 25687
rect 10425 25653 10459 25687
rect 10885 25653 10919 25687
rect 19441 25653 19475 25687
rect 31953 25653 31987 25687
rect 3249 25449 3283 25483
rect 5917 25449 5951 25483
rect 6101 25449 6135 25483
rect 7021 25449 7055 25483
rect 10149 25449 10183 25483
rect 10609 25449 10643 25483
rect 10793 25449 10827 25483
rect 12068 25449 12102 25483
rect 14105 25449 14139 25483
rect 16681 25449 16715 25483
rect 18705 25449 18739 25483
rect 1409 25381 1443 25415
rect 3065 25381 3099 25415
rect 6561 25381 6595 25415
rect 9873 25381 9907 25415
rect 2237 25313 2271 25347
rect 2789 25313 2823 25347
rect 3801 25313 3835 25347
rect 5549 25313 5583 25347
rect 6469 25313 6503 25347
rect 10241 25313 10275 25347
rect 14565 25313 14599 25347
rect 14749 25313 14783 25347
rect 16957 25313 16991 25347
rect 17233 25313 17267 25347
rect 21925 25313 21959 25347
rect 24961 25313 24995 25347
rect 28917 25313 28951 25347
rect 34069 25313 34103 25347
rect 1593 25245 1627 25279
rect 1869 25245 1903 25279
rect 2053 25245 2087 25279
rect 2145 25245 2179 25279
rect 2329 25245 2363 25279
rect 5733 25245 5767 25279
rect 5917 25245 5951 25279
rect 6377 25245 6411 25279
rect 6653 25245 6687 25279
rect 10057 25245 10091 25279
rect 11805 25245 11839 25279
rect 14933 25245 14967 25279
rect 20545 25245 20579 25279
rect 21649 25245 21683 25279
rect 21833 25245 21867 25279
rect 22753 25245 22787 25279
rect 22937 25245 22971 25279
rect 23029 25245 23063 25279
rect 30021 25245 30055 25279
rect 31125 25245 31159 25279
rect 33793 25245 33827 25279
rect 33977 25245 34011 25279
rect 4077 25177 4111 25211
rect 6989 25177 7023 25211
rect 7205 25177 7239 25211
rect 10333 25177 10367 25211
rect 10425 25177 10459 25211
rect 10625 25177 10659 25211
rect 15209 25177 15243 25211
rect 19717 25177 19751 25211
rect 21189 25177 21223 25211
rect 22293 25177 22327 25211
rect 25237 25177 25271 25211
rect 27169 25177 27203 25211
rect 30665 25177 30699 25211
rect 33333 25177 33367 25211
rect 1961 25109 1995 25143
rect 6193 25109 6227 25143
rect 6837 25109 6871 25143
rect 13553 25109 13587 25143
rect 14473 25109 14507 25143
rect 26709 25109 26743 25143
rect 1409 24905 1443 24939
rect 4353 24905 4387 24939
rect 5917 24905 5951 24939
rect 6009 24905 6043 24939
rect 14013 24905 14047 24939
rect 15669 24905 15703 24939
rect 16037 24905 16071 24939
rect 28917 24905 28951 24939
rect 34437 24905 34471 24939
rect 4721 24837 4755 24871
rect 5825 24837 5859 24871
rect 22109 24837 22143 24871
rect 3157 24769 3191 24803
rect 3249 24769 3283 24803
rect 4169 24769 4203 24803
rect 4813 24769 4847 24803
rect 5181 24769 5215 24803
rect 5365 24769 5399 24803
rect 6193 24769 6227 24803
rect 6837 24769 6871 24803
rect 11713 24769 11747 24803
rect 13921 24769 13955 24803
rect 18521 24769 18555 24803
rect 20821 24769 20855 24803
rect 21005 24769 21039 24803
rect 25881 24769 25915 24803
rect 29009 24769 29043 24803
rect 31217 24769 31251 24803
rect 2881 24701 2915 24735
rect 4905 24701 4939 24735
rect 5273 24701 5307 24735
rect 7113 24701 7147 24735
rect 13461 24701 13495 24735
rect 14197 24701 14231 24735
rect 16129 24701 16163 24735
rect 16313 24701 16347 24735
rect 18797 24701 18831 24735
rect 20361 24701 20395 24735
rect 21097 24701 21131 24735
rect 21833 24701 21867 24735
rect 23581 24701 23615 24735
rect 23673 24701 23707 24735
rect 23949 24701 23983 24735
rect 25973 24701 26007 24735
rect 26065 24701 26099 24735
rect 27169 24701 27203 24735
rect 27445 24701 27479 24735
rect 29285 24701 29319 24735
rect 31309 24701 31343 24735
rect 31493 24701 31527 24735
rect 32689 24701 32723 24735
rect 32965 24701 32999 24735
rect 20269 24633 20303 24667
rect 25513 24633 25547 24667
rect 3709 24565 3743 24599
rect 5641 24565 5675 24599
rect 8585 24565 8619 24599
rect 13553 24565 13587 24599
rect 25421 24565 25455 24599
rect 30757 24565 30791 24599
rect 30849 24565 30883 24599
rect 7389 24361 7423 24395
rect 13921 24361 13955 24395
rect 16221 24361 16255 24395
rect 22293 24361 22327 24395
rect 26157 24361 26191 24395
rect 27997 24361 28031 24395
rect 31309 24361 31343 24395
rect 34529 24361 34563 24395
rect 7481 24293 7515 24327
rect 31401 24293 31435 24327
rect 1593 24225 1627 24259
rect 3617 24225 3651 24259
rect 12173 24225 12207 24259
rect 12449 24225 12483 24259
rect 18153 24225 18187 24259
rect 20545 24225 20579 24259
rect 20821 24225 20855 24259
rect 24409 24225 24443 24259
rect 24685 24225 24719 24259
rect 28641 24225 28675 24259
rect 29377 24225 29411 24259
rect 29837 24225 29871 24259
rect 31861 24225 31895 24259
rect 32045 24225 32079 24259
rect 32781 24225 32815 24259
rect 7113 24157 7147 24191
rect 7389 24157 7423 24191
rect 7757 24157 7791 24191
rect 14473 24157 14507 24191
rect 19717 24157 19751 24191
rect 19901 24157 19935 24191
rect 19993 24157 20027 24191
rect 26249 24157 26283 24191
rect 28733 24157 28767 24191
rect 28917 24157 28951 24191
rect 29561 24157 29595 24191
rect 31769 24157 31803 24191
rect 1869 24089 1903 24123
rect 7205 24089 7239 24123
rect 7481 24089 7515 24123
rect 14749 24089 14783 24123
rect 17877 24089 17911 24123
rect 19257 24089 19291 24123
rect 24133 24089 24167 24123
rect 26525 24089 26559 24123
rect 33057 24089 33091 24123
rect 7665 24021 7699 24055
rect 16405 24021 16439 24055
rect 22845 24021 22879 24055
rect 9505 23817 9539 23851
rect 10149 23817 10183 23851
rect 13553 23817 13587 23851
rect 15485 23817 15519 23851
rect 15853 23817 15887 23851
rect 17785 23817 17819 23851
rect 18521 23817 18555 23851
rect 25329 23817 25363 23851
rect 25789 23817 25823 23851
rect 26985 23817 27019 23851
rect 27353 23817 27387 23851
rect 34345 23817 34379 23851
rect 34713 23817 34747 23851
rect 4997 23749 5031 23783
rect 5197 23749 5231 23783
rect 9137 23749 9171 23783
rect 9337 23749 9371 23783
rect 10241 23749 10275 23783
rect 15945 23749 15979 23783
rect 17417 23749 17451 23783
rect 19993 23749 20027 23783
rect 23949 23749 23983 23783
rect 25697 23749 25731 23783
rect 27445 23749 27479 23783
rect 10471 23715 10505 23749
rect 1409 23681 1443 23715
rect 1685 23681 1719 23715
rect 6561 23681 6595 23715
rect 6745 23681 6779 23715
rect 8217 23681 8251 23715
rect 8401 23681 8435 23715
rect 8677 23681 8711 23715
rect 8769 23681 8803 23715
rect 9689 23681 9723 23715
rect 9965 23681 9999 23715
rect 13461 23681 13495 23715
rect 20269 23681 20303 23715
rect 23213 23681 23247 23715
rect 23305 23681 23339 23715
rect 23489 23681 23523 23715
rect 25053 23681 25087 23715
rect 30573 23681 30607 23715
rect 30757 23681 30791 23715
rect 32597 23681 32631 23715
rect 32781 23681 32815 23715
rect 32873 23681 32907 23715
rect 33701 23681 33735 23715
rect 33885 23681 33919 23715
rect 9873 23613 9907 23647
rect 13737 23613 13771 23647
rect 16129 23613 16163 23647
rect 17141 23613 17175 23647
rect 17325 23613 17359 23647
rect 24225 23613 24259 23647
rect 25973 23613 26007 23647
rect 27537 23613 27571 23647
rect 30113 23613 30147 23647
rect 30849 23613 30883 23647
rect 32137 23613 32171 23647
rect 33241 23613 33275 23647
rect 33977 23613 34011 23647
rect 34805 23613 34839 23647
rect 34897 23613 34931 23647
rect 5181 23477 5215 23511
rect 5365 23477 5399 23511
rect 6377 23477 6411 23511
rect 8217 23477 8251 23511
rect 9321 23477 9355 23511
rect 9689 23477 9723 23511
rect 10425 23477 10459 23511
rect 10609 23477 10643 23511
rect 13093 23477 13127 23511
rect 4813 23273 4847 23307
rect 6745 23273 6779 23307
rect 8769 23273 8803 23307
rect 9137 23273 9171 23307
rect 9321 23273 9355 23307
rect 10149 23273 10183 23307
rect 13921 23273 13955 23307
rect 31677 23273 31711 23307
rect 34437 23273 34471 23307
rect 4997 23137 5031 23171
rect 5273 23137 5307 23171
rect 7021 23137 7055 23171
rect 10333 23137 10367 23171
rect 12173 23137 12207 23171
rect 12449 23137 12483 23171
rect 14565 23137 14599 23171
rect 14657 23137 14691 23171
rect 20729 23137 20763 23171
rect 22937 23137 22971 23171
rect 25237 23137 25271 23171
rect 28733 23137 28767 23171
rect 30205 23137 30239 23171
rect 32689 23137 32723 23171
rect 2789 23069 2823 23103
rect 2973 23069 3007 23103
rect 3801 23069 3835 23103
rect 3985 23069 4019 23103
rect 4721 23069 4755 23103
rect 9689 23069 9723 23103
rect 9781 23069 9815 23103
rect 9873 23069 9907 23103
rect 9965 23069 9999 23103
rect 15301 23069 15335 23103
rect 18521 23069 18555 23103
rect 18705 23069 18739 23103
rect 18797 23069 18831 23103
rect 20453 23069 20487 23103
rect 20637 23069 20671 23103
rect 21649 23069 21683 23103
rect 21833 23069 21867 23103
rect 21925 23069 21959 23103
rect 22845 23069 22879 23103
rect 27537 23069 27571 23103
rect 27721 23069 27755 23103
rect 27813 23069 27847 23103
rect 28641 23069 28675 23103
rect 29929 23069 29963 23103
rect 7297 23001 7331 23035
rect 9505 23001 9539 23035
rect 10609 23001 10643 23035
rect 15577 23001 15611 23035
rect 18061 23001 18095 23035
rect 19993 23001 20027 23035
rect 21189 23001 21223 23035
rect 22753 23001 22787 23035
rect 25513 23001 25547 23035
rect 27077 23001 27111 23035
rect 32965 23001 32999 23035
rect 2789 22933 2823 22967
rect 3893 22933 3927 22967
rect 9305 22933 9339 22967
rect 12081 22933 12115 22967
rect 14105 22933 14139 22967
rect 14473 22933 14507 22967
rect 17049 22933 17083 22967
rect 22385 22933 22419 22967
rect 26985 22933 27019 22967
rect 28181 22933 28215 22967
rect 28549 22933 28583 22967
rect 8217 22729 8251 22763
rect 8585 22729 8619 22763
rect 8677 22729 8711 22763
rect 9413 22729 9447 22763
rect 10057 22729 10091 22763
rect 10149 22729 10183 22763
rect 10517 22729 10551 22763
rect 17233 22729 17267 22763
rect 23673 22729 23707 22763
rect 28733 22729 28767 22763
rect 30757 22729 30791 22763
rect 33885 22729 33919 22763
rect 2697 22661 2731 22695
rect 3433 22661 3467 22695
rect 5181 22661 5215 22695
rect 5549 22661 5583 22695
rect 5825 22661 5859 22695
rect 6041 22661 6075 22695
rect 6377 22661 6411 22695
rect 9045 22661 9079 22695
rect 9245 22661 9279 22695
rect 18061 22661 18095 22695
rect 19901 22661 19935 22695
rect 22201 22661 22235 22695
rect 27261 22661 27295 22695
rect 32413 22661 32447 22695
rect 2053 22593 2087 22627
rect 3157 22593 3191 22627
rect 5365 22593 5399 22627
rect 5457 22593 5491 22627
rect 9505 22593 9539 22627
rect 9689 22593 9723 22627
rect 10241 22593 10275 22627
rect 10333 22593 10367 22627
rect 10517 22593 10551 22627
rect 10609 22593 10643 22627
rect 10701 22593 10735 22627
rect 10885 22593 10919 22627
rect 12265 22593 12299 22627
rect 14105 22593 14139 22627
rect 17325 22593 17359 22627
rect 19625 22593 19659 22627
rect 21925 22593 21959 22627
rect 23765 22593 23799 22627
rect 25973 22593 26007 22627
rect 29009 22593 29043 22627
rect 32137 22593 32171 22627
rect 2789 22525 2823 22559
rect 2973 22525 3007 22559
rect 8861 22525 8895 22559
rect 9597 22525 9631 22559
rect 9781 22525 9815 22559
rect 10793 22525 10827 22559
rect 12541 22525 12575 22559
rect 14381 22525 14415 22559
rect 17417 22525 17451 22559
rect 17785 22525 17819 22559
rect 19533 22525 19567 22559
rect 24041 22525 24075 22559
rect 26065 22525 26099 22559
rect 26157 22525 26191 22559
rect 26985 22525 27019 22559
rect 29285 22525 29319 22559
rect 2329 22457 2363 22491
rect 5733 22457 5767 22491
rect 21373 22457 21407 22491
rect 25605 22457 25639 22491
rect 1961 22389 1995 22423
rect 4905 22389 4939 22423
rect 6009 22389 6043 22423
rect 6193 22389 6227 22423
rect 7665 22389 7699 22423
rect 9229 22389 9263 22423
rect 14013 22389 14047 22423
rect 15853 22389 15887 22423
rect 16865 22389 16899 22423
rect 25513 22389 25547 22423
rect 1672 22185 1706 22219
rect 3801 22185 3835 22219
rect 5641 22185 5675 22219
rect 6285 22185 6319 22219
rect 6561 22185 6595 22219
rect 6745 22185 6779 22219
rect 10774 22185 10808 22219
rect 14565 22185 14599 22219
rect 15577 22185 15611 22219
rect 16668 22185 16702 22219
rect 20992 22185 21026 22219
rect 22477 22185 22511 22219
rect 24672 22185 24706 22219
rect 26157 22185 26191 22219
rect 26249 22185 26283 22219
rect 27892 22185 27926 22219
rect 29377 22185 29411 22219
rect 3157 22117 3191 22151
rect 7481 22049 7515 22083
rect 12265 22049 12299 22083
rect 15025 22049 15059 22083
rect 15117 22049 15151 22083
rect 16037 22049 16071 22083
rect 16129 22049 16163 22083
rect 18153 22049 18187 22083
rect 20729 22049 20763 22083
rect 24409 22049 24443 22083
rect 26709 22049 26743 22083
rect 26801 22049 26835 22083
rect 27629 22049 27663 22083
rect 29561 22049 29595 22083
rect 30297 22049 30331 22083
rect 1409 21981 1443 22015
rect 3801 21981 3835 22015
rect 3985 21981 4019 22015
rect 4077 21981 4111 22015
rect 4174 21981 4208 22015
rect 4629 21981 4663 22015
rect 5549 21981 5583 22015
rect 5641 21981 5675 22015
rect 5917 21981 5951 22015
rect 7297 21981 7331 22015
rect 10517 21981 10551 22015
rect 14933 21981 14967 22015
rect 16405 21981 16439 22015
rect 23489 21981 23523 22015
rect 23581 21981 23615 22015
rect 23765 21981 23799 22015
rect 24225 21981 24259 22015
rect 26617 21981 26651 22015
rect 30021 21981 30055 22015
rect 30205 21981 30239 22015
rect 4353 21913 4387 21947
rect 5365 21913 5399 21947
rect 6713 21913 6747 21947
rect 6929 21913 6963 21947
rect 15945 21913 15979 21947
rect 4451 21845 4485 21879
rect 4537 21845 4571 21879
rect 5825 21845 5859 21879
rect 6285 21845 6319 21879
rect 6469 21845 6503 21879
rect 7113 21845 7147 21879
rect 6745 21641 6779 21675
rect 9965 21641 9999 21675
rect 10517 21641 10551 21675
rect 9137 21573 9171 21607
rect 9229 21573 9263 21607
rect 9505 21573 9539 21607
rect 6561 21505 6595 21539
rect 6837 21505 6871 21539
rect 9045 21505 9079 21539
rect 9689 21505 9723 21539
rect 9781 21505 9815 21539
rect 28549 21505 28583 21539
rect 28641 21505 28675 21539
rect 30665 21505 30699 21539
rect 31493 21505 31527 21539
rect 32689 21505 32723 21539
rect 3157 21437 3191 21471
rect 3433 21437 3467 21471
rect 9413 21437 9447 21471
rect 10609 21437 10643 21471
rect 10793 21437 10827 21471
rect 28733 21437 28767 21471
rect 30757 21437 30791 21471
rect 30849 21437 30883 21471
rect 31585 21437 31619 21471
rect 31677 21437 31711 21471
rect 32781 21437 32815 21471
rect 32873 21437 32907 21471
rect 8861 21369 8895 21403
rect 4905 21301 4939 21335
rect 6377 21301 6411 21335
rect 9505 21301 9539 21335
rect 10149 21301 10183 21335
rect 28181 21301 28215 21335
rect 30297 21301 30331 21335
rect 31125 21301 31159 21335
rect 32321 21301 32355 21335
rect 4077 21097 4111 21131
rect 4629 21097 4663 21131
rect 9965 21097 9999 21131
rect 11805 21097 11839 21131
rect 29561 21097 29595 21131
rect 31493 21097 31527 21131
rect 7297 21029 7331 21063
rect 1409 20961 1443 20995
rect 6101 20961 6135 20995
rect 6929 20961 6963 20995
rect 7021 20961 7055 20995
rect 7849 20961 7883 20995
rect 9045 20961 9079 20995
rect 9321 20961 9355 20995
rect 10057 20961 10091 20995
rect 10333 20961 10367 20995
rect 21373 20961 21407 20995
rect 25145 20961 25179 20995
rect 27629 20961 27663 20995
rect 31033 20961 31067 20995
rect 31309 20961 31343 20995
rect 33241 20961 33275 20995
rect 3801 20893 3835 20927
rect 3893 20893 3927 20927
rect 4077 20893 4111 20927
rect 6377 20893 6411 20927
rect 6837 20893 6871 20927
rect 7297 20893 7331 20927
rect 7481 20893 7515 20927
rect 7665 20893 7699 20927
rect 8033 20893 8067 20927
rect 8309 20893 8343 20927
rect 8401 20893 8435 20927
rect 8585 20893 8619 20927
rect 8953 20893 8987 20927
rect 9413 20893 9447 20927
rect 9781 20893 9815 20927
rect 9965 20893 9999 20927
rect 16773 20893 16807 20927
rect 16865 20893 16899 20927
rect 22569 20893 22603 20927
rect 22753 20893 22787 20927
rect 22845 20893 22879 20927
rect 24869 20893 24903 20927
rect 25053 20893 25087 20927
rect 27353 20893 27387 20927
rect 33793 20893 33827 20927
rect 33977 20893 34011 20927
rect 34069 20893 34103 20927
rect 34713 20893 34747 20927
rect 1685 20825 1719 20859
rect 16497 20825 16531 20859
rect 17141 20825 17175 20859
rect 22109 20825 22143 20859
rect 24409 20825 24443 20859
rect 32965 20825 32999 20859
rect 33333 20825 33367 20859
rect 34989 20825 35023 20859
rect 3157 20757 3191 20791
rect 6469 20757 6503 20791
rect 7757 20757 7791 20791
rect 7941 20757 7975 20791
rect 8769 20757 8803 20791
rect 9137 20757 9171 20791
rect 9597 20757 9631 20791
rect 15025 20757 15059 20791
rect 18613 20757 18647 20791
rect 20729 20757 20763 20791
rect 21097 20757 21131 20791
rect 21189 20757 21223 20791
rect 29101 20757 29135 20791
rect 36461 20757 36495 20791
rect 8125 20553 8159 20587
rect 8677 20553 8711 20587
rect 9597 20553 9631 20587
rect 16129 20553 16163 20587
rect 23581 20553 23615 20587
rect 23673 20553 23707 20587
rect 29745 20553 29779 20587
rect 32321 20553 32355 20587
rect 6653 20485 6687 20519
rect 17509 20485 17543 20519
rect 22109 20485 22143 20519
rect 25145 20485 25179 20519
rect 26249 20485 26283 20519
rect 31217 20485 31251 20519
rect 33793 20485 33827 20519
rect 35173 20485 35207 20519
rect 2237 20417 2271 20451
rect 8585 20417 8619 20451
rect 9229 20417 9263 20451
rect 11345 20417 11379 20451
rect 16037 20417 16071 20451
rect 17969 20417 18003 20451
rect 18153 20417 18187 20451
rect 26157 20417 26191 20451
rect 28733 20417 28767 20451
rect 34069 20417 34103 20451
rect 34437 20417 34471 20451
rect 34529 20417 34563 20451
rect 34713 20417 34747 20451
rect 1869 20349 1903 20383
rect 2329 20349 2363 20383
rect 6377 20349 6411 20383
rect 8769 20349 8803 20383
rect 9045 20349 9079 20383
rect 11069 20349 11103 20383
rect 13829 20349 13863 20383
rect 14105 20349 14139 20383
rect 16313 20349 16347 20383
rect 18245 20349 18279 20383
rect 19809 20349 19843 20383
rect 20085 20349 20119 20383
rect 21557 20349 21591 20383
rect 21833 20349 21867 20383
rect 25421 20349 25455 20383
rect 26341 20349 26375 20383
rect 28457 20349 28491 20383
rect 31493 20349 31527 20383
rect 8217 20281 8251 20315
rect 9413 20281 9447 20315
rect 15669 20281 15703 20315
rect 15577 20213 15611 20247
rect 25789 20213 25823 20247
rect 26985 20213 27019 20247
rect 2973 20009 3007 20043
rect 7941 20009 7975 20043
rect 8125 20009 8159 20043
rect 10149 20009 10183 20043
rect 18429 20009 18463 20043
rect 24041 20009 24075 20043
rect 26525 20009 26559 20043
rect 9781 19873 9815 19907
rect 19257 19873 19291 19907
rect 24777 19873 24811 19907
rect 27721 19873 27755 19907
rect 28457 19873 28491 19907
rect 35449 19873 35483 19907
rect 2421 19805 2455 19839
rect 2605 19805 2639 19839
rect 9965 19805 9999 19839
rect 16681 19805 16715 19839
rect 22293 19805 22327 19839
rect 27077 19805 27111 19839
rect 27261 19805 27295 19839
rect 27353 19805 27387 19839
rect 28181 19805 28215 19839
rect 28365 19805 28399 19839
rect 30021 19805 30055 19839
rect 30205 19805 30239 19839
rect 30297 19805 30331 19839
rect 31125 19805 31159 19839
rect 31309 19805 31343 19839
rect 31401 19805 31435 19839
rect 35173 19805 35207 19839
rect 35357 19805 35391 19839
rect 3157 19737 3191 19771
rect 7757 19737 7791 19771
rect 7957 19737 7991 19771
rect 16957 19737 16991 19771
rect 19533 19737 19567 19771
rect 22569 19737 22603 19771
rect 25053 19737 25087 19771
rect 26617 19737 26651 19771
rect 29561 19737 29595 19771
rect 30665 19737 30699 19771
rect 34713 19737 34747 19771
rect 2513 19669 2547 19703
rect 2789 19669 2823 19703
rect 2957 19669 2991 19703
rect 21005 19669 21039 19703
rect 1862 19465 1896 19499
rect 8217 19465 8251 19499
rect 23305 19465 23339 19499
rect 23673 19465 23707 19499
rect 31217 19465 31251 19499
rect 35817 19465 35851 19499
rect 1777 19397 1811 19431
rect 1961 19397 1995 19431
rect 16681 19397 16715 19431
rect 18153 19397 18187 19431
rect 18337 19397 18371 19431
rect 20177 19397 20211 19431
rect 26525 19397 26559 19431
rect 1685 19329 1719 19363
rect 4169 19329 4203 19363
rect 4353 19329 4387 19363
rect 6193 19329 6227 19363
rect 9965 19329 9999 19363
rect 14105 19329 14139 19363
rect 17141 19329 17175 19363
rect 17325 19329 17359 19363
rect 17417 19329 17451 19363
rect 20637 19329 20671 19363
rect 20821 19329 20855 19363
rect 20913 19329 20947 19363
rect 29653 19329 29687 19363
rect 29745 19329 29779 19363
rect 30941 19329 30975 19363
rect 31585 19329 31619 19363
rect 34069 19329 34103 19363
rect 2053 19261 2087 19295
rect 2329 19261 2363 19295
rect 4261 19261 4295 19295
rect 5917 19261 5951 19295
rect 9689 19261 9723 19295
rect 14381 19261 14415 19295
rect 18429 19261 18463 19295
rect 23765 19261 23799 19295
rect 23857 19261 23891 19295
rect 25053 19261 25087 19295
rect 26801 19261 26835 19295
rect 31677 19261 31711 19295
rect 31861 19261 31895 19295
rect 34345 19261 34379 19295
rect 17877 19193 17911 19227
rect 3801 19125 3835 19159
rect 4445 19125 4479 19159
rect 15853 19125 15887 19159
rect 28365 19125 28399 19159
rect 8769 18921 8803 18955
rect 18705 18921 18739 18955
rect 29285 18921 29319 18955
rect 31309 18921 31343 18955
rect 21465 18853 21499 18887
rect 35357 18853 35391 18887
rect 1409 18785 1443 18819
rect 4077 18785 4111 18819
rect 4629 18785 4663 18819
rect 5089 18785 5123 18819
rect 6653 18785 6687 18819
rect 7297 18785 7331 18819
rect 15025 18785 15059 18819
rect 15761 18785 15795 18819
rect 16589 18785 16623 18819
rect 16681 18785 16715 18819
rect 19533 18785 19567 18819
rect 21925 18785 21959 18819
rect 29561 18785 29595 18819
rect 29837 18785 29871 18819
rect 32045 18785 32079 18819
rect 32321 18785 32355 18819
rect 3801 18717 3835 18751
rect 4169 18717 4203 18751
rect 4721 18717 4755 18751
rect 6929 18717 6963 18751
rect 7021 18717 7055 18751
rect 15485 18717 15519 18751
rect 15669 18717 15703 18751
rect 16957 18717 16991 18751
rect 24685 18717 24719 18751
rect 24803 18717 24837 18751
rect 24961 18717 24995 18751
rect 26157 18717 26191 18751
rect 26249 18717 26283 18751
rect 27537 18717 27571 18751
rect 35081 18717 35115 18751
rect 1685 18649 1719 18683
rect 4286 18649 4320 18683
rect 17233 18649 17267 18683
rect 19809 18649 19843 18683
rect 22017 18649 22051 18683
rect 25421 18649 25455 18683
rect 25513 18649 25547 18683
rect 26019 18649 26053 18683
rect 27813 18649 27847 18683
rect 34805 18649 34839 18683
rect 3157 18581 3191 18615
rect 4445 18581 4479 18615
rect 5181 18581 5215 18615
rect 16129 18581 16163 18615
rect 16497 18581 16531 18615
rect 21281 18581 21315 18615
rect 21925 18581 21959 18615
rect 33793 18581 33827 18615
rect 34897 18581 34931 18615
rect 3985 18377 4019 18411
rect 4153 18377 4187 18411
rect 16405 18377 16439 18411
rect 18043 18377 18077 18411
rect 28733 18377 28767 18411
rect 4353 18309 4387 18343
rect 6193 18309 6227 18343
rect 7757 18309 7791 18343
rect 9505 18309 9539 18343
rect 14933 18309 14967 18343
rect 18337 18309 18371 18343
rect 18521 18309 18555 18343
rect 20269 18309 20303 18343
rect 25605 18309 25639 18343
rect 32873 18309 32907 18343
rect 1593 18241 1627 18275
rect 2237 18241 2271 18275
rect 9597 18241 9631 18275
rect 14657 18241 14691 18275
rect 20729 18241 20763 18275
rect 20913 18241 20947 18275
rect 22293 18241 22327 18275
rect 25881 18241 25915 18275
rect 30573 18241 30607 18275
rect 31309 18241 31343 18275
rect 31493 18241 31527 18275
rect 1869 18173 1903 18207
rect 2329 18173 2363 18207
rect 9873 18173 9907 18207
rect 18613 18173 18647 18207
rect 21005 18173 21039 18207
rect 22569 18173 22603 18207
rect 24041 18173 24075 18207
rect 24133 18173 24167 18207
rect 26985 18173 27019 18207
rect 27261 18173 27295 18207
rect 31217 18173 31251 18207
rect 31953 18173 31987 18207
rect 32597 18173 32631 18207
rect 34345 18173 34379 18207
rect 1409 18037 1443 18071
rect 4169 18037 4203 18071
rect 4721 18037 4755 18071
rect 11345 18037 11379 18071
rect 29101 18037 29135 18071
rect 1869 17833 1903 17867
rect 5089 17833 5123 17867
rect 10241 17833 10275 17867
rect 10701 17833 10735 17867
rect 19073 17833 19107 17867
rect 22385 17833 22419 17867
rect 23397 17833 23431 17867
rect 24777 17833 24811 17867
rect 28365 17833 28399 17867
rect 31861 17833 31895 17867
rect 33333 17833 33367 17867
rect 4261 17765 4295 17799
rect 11253 17765 11287 17799
rect 6285 17697 6319 17731
rect 17325 17697 17359 17731
rect 20637 17697 20671 17731
rect 23949 17697 23983 17731
rect 26525 17697 26559 17731
rect 28825 17697 28859 17731
rect 30113 17697 30147 17731
rect 33793 17697 33827 17731
rect 33885 17697 33919 17731
rect 2053 17629 2087 17663
rect 3985 17629 4019 17663
rect 4353 17629 4387 17663
rect 4537 17629 4571 17663
rect 4629 17629 4663 17663
rect 5089 17629 5123 17663
rect 5365 17629 5399 17663
rect 10057 17629 10091 17663
rect 10241 17629 10275 17663
rect 10977 17629 11011 17663
rect 11253 17629 11287 17663
rect 15761 17629 15795 17663
rect 15945 17629 15979 17663
rect 16037 17629 16071 17663
rect 23765 17629 23799 17663
rect 23857 17629 23891 17663
rect 26801 17629 26835 17663
rect 27353 17629 27387 17663
rect 32413 17629 32447 17663
rect 4261 17561 4295 17595
rect 6561 17561 6595 17595
rect 10685 17561 10719 17595
rect 10885 17561 10919 17595
rect 15301 17561 15335 17595
rect 17601 17561 17635 17595
rect 20913 17561 20947 17595
rect 26249 17561 26283 17595
rect 28181 17561 28215 17595
rect 28917 17561 28951 17595
rect 30389 17561 30423 17595
rect 4077 17493 4111 17527
rect 4445 17493 4479 17527
rect 5273 17493 5307 17527
rect 8033 17493 8067 17527
rect 10517 17493 10551 17527
rect 11069 17493 11103 17527
rect 28825 17493 28859 17527
rect 33793 17493 33827 17527
rect 5825 17289 5859 17323
rect 7113 17289 7147 17323
rect 18705 17289 18739 17323
rect 19073 17289 19107 17323
rect 23397 17289 23431 17323
rect 26801 17289 26835 17323
rect 35725 17289 35759 17323
rect 3617 17221 3651 17255
rect 3817 17221 3851 17255
rect 4353 17221 4387 17255
rect 14565 17221 14599 17255
rect 20637 17221 20671 17255
rect 22569 17221 22603 17255
rect 29745 17221 29779 17255
rect 31677 17221 31711 17255
rect 1685 17153 1719 17187
rect 4077 17153 4111 17187
rect 7481 17153 7515 17187
rect 7757 17153 7791 17187
rect 9781 17153 9815 17187
rect 9965 17153 9999 17187
rect 10425 17153 10459 17187
rect 14289 17153 14323 17187
rect 20729 17153 20763 17187
rect 21833 17153 21867 17187
rect 25053 17153 25087 17187
rect 29009 17153 29043 17187
rect 29561 17153 29595 17187
rect 31953 17153 31987 17187
rect 1961 17085 1995 17119
rect 7573 17085 7607 17119
rect 8033 17085 8067 17119
rect 10517 17085 10551 17119
rect 16865 17085 16899 17119
rect 17141 17085 17175 17119
rect 18613 17085 18647 17119
rect 19165 17085 19199 17119
rect 19349 17085 19383 17119
rect 20821 17085 20855 17119
rect 23305 17085 23339 17119
rect 23489 17085 23523 17119
rect 25329 17085 25363 17119
rect 29837 17085 29871 17119
rect 32137 17085 32171 17119
rect 32413 17085 32447 17119
rect 33977 17085 34011 17119
rect 34253 17085 34287 17119
rect 3433 16949 3467 16983
rect 3801 16949 3835 16983
rect 3985 16949 4019 16983
rect 9505 16949 9539 16983
rect 9597 16949 9631 16983
rect 10793 16949 10827 16983
rect 16037 16949 16071 16983
rect 20269 16949 20303 16983
rect 22937 16949 22971 16983
rect 29285 16949 29319 16983
rect 30205 16949 30239 16983
rect 33885 16949 33919 16983
rect 1777 16745 1811 16779
rect 8309 16745 8343 16779
rect 12357 16745 12391 16779
rect 20453 16745 20487 16779
rect 25132 16745 25166 16779
rect 26801 16745 26835 16779
rect 29285 16745 29319 16779
rect 30849 16677 30883 16711
rect 2237 16609 2271 16643
rect 4537 16609 4571 16643
rect 5181 16609 5215 16643
rect 10609 16609 10643 16643
rect 10885 16609 10919 16643
rect 14105 16609 14139 16643
rect 14381 16609 14415 16643
rect 16589 16609 16623 16643
rect 21925 16609 21959 16643
rect 22201 16609 22235 16643
rect 22385 16609 22419 16643
rect 24869 16609 24903 16643
rect 27537 16609 27571 16643
rect 27813 16609 27847 16643
rect 31677 16609 31711 16643
rect 32413 16609 32447 16643
rect 32689 16609 32723 16643
rect 34253 16609 34287 16643
rect 36461 16609 36495 16643
rect 2145 16541 2179 16575
rect 3801 16541 3835 16575
rect 4077 16541 4111 16575
rect 4169 16541 4203 16575
rect 4445 16541 4479 16575
rect 4721 16541 4755 16575
rect 4813 16541 4847 16575
rect 8493 16541 8527 16575
rect 8585 16541 8619 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 17785 16541 17819 16575
rect 18245 16541 18279 16575
rect 18429 16541 18463 16575
rect 18521 16541 18555 16575
rect 27077 16541 27111 16575
rect 31769 16541 31803 16575
rect 31953 16541 31987 16575
rect 3893 16473 3927 16507
rect 4905 16473 4939 16507
rect 5457 16473 5491 16507
rect 7205 16473 7239 16507
rect 9045 16473 9079 16507
rect 17325 16473 17359 16507
rect 22661 16473 22695 16507
rect 27353 16473 27387 16507
rect 29561 16473 29595 16507
rect 33425 16473 33459 16507
rect 33517 16473 33551 16507
rect 36645 16473 36679 16507
rect 4353 16405 4387 16439
rect 15853 16405 15887 16439
rect 24133 16405 24167 16439
rect 26617 16405 26651 16439
rect 27261 16405 27295 16439
rect 3893 16201 3927 16235
rect 4077 16201 4111 16235
rect 20821 16201 20855 16235
rect 30389 16201 30423 16235
rect 32689 16201 32723 16235
rect 33517 16201 33551 16235
rect 33977 16201 34011 16235
rect 10517 16133 10551 16167
rect 19349 16133 19383 16167
rect 22661 16133 22695 16167
rect 25973 16133 26007 16167
rect 26157 16133 26191 16167
rect 26985 16133 27019 16167
rect 27721 16133 27755 16167
rect 33609 16133 33643 16167
rect 2243 16065 2277 16099
rect 2421 16065 2455 16099
rect 3709 16065 3743 16099
rect 3801 16065 3835 16099
rect 14657 16065 14691 16099
rect 15209 16065 15243 16099
rect 15393 16065 15427 16099
rect 18429 16065 18463 16099
rect 19073 16065 19107 16099
rect 21649 16065 21683 16099
rect 23121 16065 23155 16099
rect 23305 16065 23339 16099
rect 28641 16065 28675 16099
rect 30481 16065 30515 16099
rect 31769 16065 31803 16099
rect 7481 15997 7515 16031
rect 14749 15997 14783 16031
rect 15485 15997 15519 16031
rect 18153 15997 18187 16031
rect 23397 15997 23431 16031
rect 23765 15997 23799 16031
rect 24041 15997 24075 16031
rect 25513 15997 25547 16031
rect 26249 15997 26283 16031
rect 28917 15997 28951 16031
rect 30849 15997 30883 16031
rect 32597 15997 32631 16031
rect 32781 15997 32815 16031
rect 33333 15997 33367 16031
rect 3525 15929 3559 15963
rect 7113 15929 7147 15963
rect 10793 15929 10827 15963
rect 25697 15929 25731 15963
rect 2421 15861 2455 15895
rect 7021 15861 7055 15895
rect 10977 15861 11011 15895
rect 16681 15861 16715 15895
rect 32229 15861 32263 15895
rect 3433 15657 3467 15691
rect 4353 15657 4387 15691
rect 10517 15657 10551 15691
rect 15853 15657 15887 15691
rect 15945 15657 15979 15691
rect 23581 15657 23615 15691
rect 28733 15657 28767 15691
rect 31309 15589 31343 15623
rect 32597 15589 32631 15623
rect 1685 15521 1719 15555
rect 3157 15521 3191 15555
rect 7205 15521 7239 15555
rect 10609 15521 10643 15555
rect 10885 15521 10919 15555
rect 14381 15521 14415 15555
rect 16405 15521 16439 15555
rect 16497 15521 16531 15555
rect 16865 15521 16899 15555
rect 18061 15521 18095 15555
rect 18797 15521 18831 15555
rect 20177 15521 20211 15555
rect 24409 15521 24443 15555
rect 25145 15521 25179 15555
rect 28181 15521 28215 15555
rect 29561 15521 29595 15555
rect 29837 15521 29871 15555
rect 33057 15521 33091 15555
rect 1409 15453 1443 15487
rect 3249 15453 3283 15487
rect 3433 15453 3467 15487
rect 4077 15453 4111 15487
rect 6929 15453 6963 15487
rect 9321 15453 9355 15487
rect 9597 15453 9631 15487
rect 9781 15453 9815 15487
rect 10333 15453 10367 15487
rect 14105 15453 14139 15487
rect 16313 15453 16347 15487
rect 18153 15453 18187 15487
rect 18337 15453 18371 15487
rect 20637 15453 20671 15487
rect 21189 15453 21223 15487
rect 21373 15453 21407 15487
rect 21465 15453 21499 15487
rect 21833 15453 21867 15487
rect 24869 15453 24903 15487
rect 25053 15453 25087 15487
rect 27997 15453 28031 15487
rect 31861 15453 31895 15487
rect 32045 15453 32079 15487
rect 32137 15453 32171 15487
rect 33149 15453 33183 15487
rect 3801 15385 3835 15419
rect 9505 15385 9539 15419
rect 9965 15385 9999 15419
rect 10241 15385 10275 15419
rect 17693 15385 17727 15419
rect 20729 15385 20763 15419
rect 22109 15385 22143 15419
rect 29009 15385 29043 15419
rect 29285 15385 29319 15419
rect 31401 15385 31435 15419
rect 33057 15385 33091 15419
rect 3985 15317 4019 15351
rect 4169 15317 4203 15351
rect 8677 15317 8711 15351
rect 9137 15317 9171 15351
rect 9689 15317 9723 15351
rect 10149 15317 10183 15351
rect 12357 15317 12391 15351
rect 27629 15317 27663 15351
rect 28089 15317 28123 15351
rect 29193 15317 29227 15351
rect 3525 15113 3559 15147
rect 7297 15113 7331 15147
rect 7665 15113 7699 15147
rect 7757 15113 7791 15147
rect 11069 15113 11103 15147
rect 22937 15113 22971 15147
rect 23305 15113 23339 15147
rect 28825 15113 28859 15147
rect 30205 15113 30239 15147
rect 3157 15045 3191 15079
rect 3357 15045 3391 15079
rect 5733 15045 5767 15079
rect 7389 15045 7423 15079
rect 20453 15045 20487 15079
rect 22753 15045 22787 15079
rect 25973 15045 26007 15079
rect 27353 15045 27387 15079
rect 5273 14977 5307 15011
rect 5549 14977 5583 15011
rect 5917 14977 5951 15011
rect 6009 14967 6043 15001
rect 6193 14977 6227 15011
rect 7481 14977 7515 15011
rect 8217 14977 8251 15011
rect 10609 14977 10643 15011
rect 10885 14977 10919 15011
rect 15485 14977 15519 15011
rect 15669 14977 15703 15011
rect 20729 14977 20763 15011
rect 21925 14977 21959 15011
rect 26065 14977 26099 15011
rect 31493 14977 31527 15011
rect 5457 14909 5491 14943
rect 7941 14909 7975 14943
rect 8033 14909 8067 14943
rect 8125 14909 8159 14943
rect 8585 14909 8619 14943
rect 8861 14909 8895 14943
rect 10333 14909 10367 14943
rect 10701 14909 10735 14943
rect 10793 14909 10827 14943
rect 15025 14909 15059 14943
rect 15761 14909 15795 14943
rect 16681 14909 16715 14943
rect 16957 14909 16991 14943
rect 18981 14909 19015 14943
rect 23397 14909 23431 14943
rect 23581 14909 23615 14943
rect 25973 14909 26007 14943
rect 27077 14909 27111 14943
rect 32597 14909 32631 14943
rect 32873 14909 32907 14943
rect 34437 14909 34471 14943
rect 34713 14909 34747 14943
rect 7113 14841 7147 14875
rect 3341 14773 3375 14807
rect 5089 14773 5123 14807
rect 6101 14773 6135 14807
rect 18429 14773 18463 14807
rect 25513 14773 25547 14807
rect 34345 14773 34379 14807
rect 36185 14773 36219 14807
rect 6745 14569 6779 14603
rect 11621 14569 11655 14603
rect 14105 14569 14139 14603
rect 23949 14569 23983 14603
rect 27997 14569 28031 14603
rect 29929 14569 29963 14603
rect 33517 14569 33551 14603
rect 3433 14501 3467 14535
rect 1685 14433 1719 14467
rect 1961 14433 1995 14467
rect 4997 14433 5031 14467
rect 5273 14433 5307 14467
rect 9505 14433 9539 14467
rect 9873 14433 9907 14467
rect 15853 14433 15887 14467
rect 18613 14433 18647 14467
rect 22201 14433 22235 14467
rect 24409 14433 24443 14467
rect 31401 14433 31435 14467
rect 31677 14433 31711 14467
rect 31769 14433 31803 14467
rect 32045 14433 32079 14467
rect 34713 14433 34747 14467
rect 35449 14433 35483 14467
rect 1593 14365 1627 14399
rect 3157 14365 3191 14399
rect 3801 14365 3835 14399
rect 3985 14365 4019 14399
rect 9413 14365 9447 14399
rect 26249 14365 26283 14399
rect 35173 14365 35207 14399
rect 35357 14365 35391 14399
rect 3433 14297 3467 14331
rect 10149 14297 10183 14331
rect 15577 14297 15611 14331
rect 18337 14297 18371 14331
rect 20361 14297 20395 14331
rect 22477 14297 22511 14331
rect 24685 14297 24719 14331
rect 26525 14297 26559 14331
rect 3249 14229 3283 14263
rect 3893 14229 3927 14263
rect 9781 14229 9815 14263
rect 16865 14229 16899 14263
rect 21833 14229 21867 14263
rect 26157 14229 26191 14263
rect 1409 14025 1443 14059
rect 2973 14025 3007 14059
rect 17601 14025 17635 14059
rect 17969 14025 18003 14059
rect 18061 14025 18095 14059
rect 19625 14025 19659 14059
rect 26985 14025 27019 14059
rect 27353 14025 27387 14059
rect 4445 13957 4479 13991
rect 9045 13957 9079 13991
rect 18429 13957 18463 13991
rect 22937 13957 22971 13991
rect 25237 13957 25271 13991
rect 32321 13957 32355 13991
rect 33057 13957 33091 13991
rect 1593 13889 1627 13923
rect 4721 13889 4755 13923
rect 5733 13889 5767 13923
rect 6377 13889 6411 13923
rect 9229 13889 9263 13923
rect 9413 13889 9447 13923
rect 18889 13889 18923 13923
rect 19073 13889 19107 13923
rect 19165 13889 19199 13923
rect 21373 13889 21407 13923
rect 22293 13889 22327 13923
rect 22477 13889 22511 13923
rect 23397 13889 23431 13923
rect 23581 13889 23615 13923
rect 23673 13889 23707 13923
rect 24961 13889 24995 13923
rect 29653 13889 29687 13923
rect 29837 13889 29871 13923
rect 32229 13889 32263 13923
rect 33517 13889 33551 13923
rect 33701 13889 33735 13923
rect 33793 13889 33827 13923
rect 5641 13821 5675 13855
rect 8125 13821 8159 13855
rect 14289 13821 14323 13855
rect 14565 13821 14599 13855
rect 18153 13821 18187 13855
rect 21097 13821 21131 13855
rect 21833 13821 21867 13855
rect 22569 13821 22603 13855
rect 26709 13821 26743 13855
rect 27445 13821 27479 13855
rect 27629 13821 27663 13855
rect 28917 13821 28951 13855
rect 29193 13821 29227 13855
rect 29561 13821 29595 13855
rect 30297 13821 30331 13855
rect 32413 13821 32447 13855
rect 6009 13685 6043 13719
rect 6634 13685 6668 13719
rect 16037 13685 16071 13719
rect 32781 13685 32815 13719
rect 3341 13481 3375 13515
rect 22569 13481 22603 13515
rect 32413 13481 32447 13515
rect 28089 13413 28123 13447
rect 1593 13345 1627 13379
rect 1869 13345 1903 13379
rect 15117 13345 15151 13379
rect 15853 13345 15887 13379
rect 16773 13345 16807 13379
rect 20821 13345 20855 13379
rect 24409 13345 24443 13379
rect 25145 13345 25179 13379
rect 28641 13345 28675 13379
rect 32321 13345 32355 13379
rect 34161 13345 34195 13379
rect 35265 13345 35299 13379
rect 15577 13277 15611 13311
rect 15761 13277 15795 13311
rect 24869 13277 24903 13311
rect 25053 13277 25087 13311
rect 17049 13209 17083 13243
rect 21097 13209 21131 13243
rect 28365 13209 28399 13243
rect 28549 13209 28583 13243
rect 32045 13209 32079 13243
rect 33885 13209 33919 13243
rect 35357 13209 35391 13243
rect 18521 13141 18555 13175
rect 30573 13141 30607 13175
rect 34787 13141 34821 13175
rect 35265 13141 35299 13175
rect 24961 12937 24995 12971
rect 25421 12937 25455 12971
rect 28549 12937 28583 12971
rect 30021 12869 30055 12903
rect 32137 12869 32171 12903
rect 33701 12869 33735 12903
rect 14381 12801 14415 12835
rect 18889 12801 18923 12835
rect 21833 12801 21867 12835
rect 22293 12801 22327 12835
rect 22477 12801 22511 12835
rect 22569 12801 22603 12835
rect 23213 12801 23247 12835
rect 27353 12801 27387 12835
rect 30665 12801 30699 12835
rect 30757 12801 30791 12835
rect 30941 12801 30975 12835
rect 32597 12801 32631 12835
rect 32781 12801 32815 12835
rect 14657 12733 14691 12767
rect 18429 12733 18463 12767
rect 18981 12733 19015 12767
rect 19257 12733 19291 12767
rect 20729 12733 20763 12767
rect 23489 12733 23523 12767
rect 25513 12733 25547 12767
rect 25697 12733 25731 12767
rect 27445 12733 27479 12767
rect 27537 12733 27571 12767
rect 30297 12733 30331 12767
rect 31401 12733 31435 12767
rect 32873 12733 32907 12767
rect 33425 12733 33459 12767
rect 25053 12665 25087 12699
rect 16129 12597 16163 12631
rect 26985 12597 27019 12631
rect 35173 12597 35207 12631
rect 20992 12393 21026 12427
rect 22569 12393 22603 12427
rect 29561 12393 29595 12427
rect 32781 12393 32815 12427
rect 23029 12257 23063 12291
rect 23213 12257 23247 12291
rect 24133 12257 24167 12291
rect 28365 12257 28399 12291
rect 31309 12257 31343 12291
rect 35449 12257 35483 12291
rect 15117 12189 15151 12223
rect 15577 12189 15611 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 18245 12189 18279 12223
rect 19625 12189 19659 12223
rect 20085 12189 20119 12223
rect 20269 12189 20303 12223
rect 20361 12189 20395 12223
rect 20729 12189 20763 12223
rect 25053 12189 25087 12223
rect 28641 12189 28675 12223
rect 34529 12189 34563 12223
rect 35173 12189 35207 12223
rect 35357 12189 35391 12223
rect 17969 12121 18003 12155
rect 26617 12121 26651 12155
rect 31033 12121 31067 12155
rect 34253 12121 34287 12155
rect 34713 12121 34747 12155
rect 16497 12053 16531 12087
rect 22477 12053 22511 12087
rect 22937 12053 22971 12087
rect 23489 12053 23523 12087
rect 23857 12053 23891 12087
rect 23949 12053 23983 12087
rect 26893 12053 26927 12087
rect 15669 11849 15703 11883
rect 16129 11849 16163 11883
rect 16221 11849 16255 11883
rect 24317 11849 24351 11883
rect 27261 11849 27295 11883
rect 17509 11781 17543 11815
rect 22845 11781 22879 11815
rect 17969 11713 18003 11747
rect 18153 11713 18187 11747
rect 18245 11713 18279 11747
rect 29009 11713 29043 11747
rect 30665 11713 30699 11747
rect 31217 11713 31251 11747
rect 31585 11713 31619 11747
rect 13921 11645 13955 11679
rect 14197 11645 14231 11679
rect 16313 11645 16347 11679
rect 18613 11645 18647 11679
rect 18889 11645 18923 11679
rect 22569 11645 22603 11679
rect 24409 11645 24443 11679
rect 24685 11645 24719 11679
rect 28733 11645 28767 11679
rect 31309 11645 31343 11679
rect 31493 11645 31527 11679
rect 31677 11645 31711 11679
rect 31769 11645 31803 11679
rect 15761 11577 15795 11611
rect 20361 11509 20395 11543
rect 26157 11509 26191 11543
rect 30849 11509 30883 11543
rect 31125 11509 31159 11543
rect 24685 11305 24719 11339
rect 26249 11305 26283 11339
rect 28469 11305 28503 11339
rect 31658 11305 31692 11339
rect 33149 11305 33183 11339
rect 16313 11237 16347 11271
rect 26985 11237 27019 11271
rect 18061 11169 18095 11203
rect 18797 11169 18831 11203
rect 21005 11169 21039 11203
rect 21281 11169 21315 11203
rect 23765 11169 23799 11203
rect 23857 11169 23891 11203
rect 25329 11169 25363 11203
rect 26709 11169 26743 11203
rect 28733 11169 28767 11203
rect 29561 11169 29595 11203
rect 29837 11169 29871 11203
rect 31401 11169 31435 11203
rect 19257 11101 19291 11135
rect 22017 11101 22051 11135
rect 22477 11101 22511 11135
rect 22569 11101 22603 11135
rect 22753 11101 22787 11135
rect 23673 11101 23707 11135
rect 25053 11101 25087 11135
rect 26801 11101 26835 11135
rect 33701 11101 33735 11135
rect 33885 11101 33919 11135
rect 33977 11101 34011 11135
rect 34345 11101 34379 11135
rect 17785 11033 17819 11067
rect 18521 11033 18555 11067
rect 19533 11033 19567 11067
rect 23213 11033 23247 11067
rect 26709 11033 26743 11067
rect 33241 11033 33275 11067
rect 18153 10965 18187 10999
rect 18613 10965 18647 10999
rect 23305 10965 23339 10999
rect 25145 10965 25179 10999
rect 31309 10965 31343 10999
rect 34437 10965 34471 10999
rect 15485 10761 15519 10795
rect 15945 10761 15979 10795
rect 16037 10761 16071 10795
rect 26341 10761 26375 10795
rect 30395 10761 30429 10795
rect 18245 10693 18279 10727
rect 21097 10693 21131 10727
rect 26433 10693 26467 10727
rect 30481 10693 30515 10727
rect 31677 10693 31711 10727
rect 31861 10693 31895 10727
rect 32965 10693 32999 10727
rect 13737 10625 13771 10659
rect 17601 10625 17635 10659
rect 17785 10625 17819 10659
rect 18889 10625 18923 10659
rect 22017 10625 22051 10659
rect 22845 10625 22879 10659
rect 23305 10625 23339 10659
rect 25145 10625 25179 10659
rect 25237 10625 25271 10659
rect 27445 10625 27479 10659
rect 30297 10625 30331 10659
rect 30573 10625 30607 10659
rect 31493 10625 31527 10659
rect 31953 10625 31987 10659
rect 32689 10625 32723 10659
rect 14013 10557 14047 10591
rect 16221 10557 16255 10591
rect 17509 10557 17543 10591
rect 21189 10557 21223 10591
rect 21373 10557 21407 10591
rect 23397 10557 23431 10591
rect 23489 10557 23523 10591
rect 25421 10557 25455 10591
rect 26249 10557 26283 10591
rect 28181 10557 28215 10591
rect 28457 10557 28491 10591
rect 28733 10557 28767 10591
rect 31217 10557 31251 10591
rect 34529 10557 34563 10591
rect 34805 10557 34839 10591
rect 15577 10489 15611 10523
rect 31677 10489 31711 10523
rect 20177 10421 20211 10455
rect 20729 10421 20763 10455
rect 22937 10421 22971 10455
rect 24777 10421 24811 10455
rect 26801 10421 26835 10455
rect 30205 10421 30239 10455
rect 34437 10421 34471 10455
rect 36277 10421 36311 10455
rect 17877 10217 17911 10251
rect 20900 10217 20934 10251
rect 22385 10217 22419 10251
rect 26157 10217 26191 10251
rect 30297 10217 30331 10251
rect 31769 10217 31803 10251
rect 34989 10217 35023 10251
rect 35449 10217 35483 10251
rect 29929 10149 29963 10183
rect 16405 10081 16439 10115
rect 19073 10081 19107 10115
rect 20085 10081 20119 10115
rect 20637 10081 20671 10115
rect 23305 10081 23339 10115
rect 24409 10081 24443 10115
rect 24685 10081 24719 10115
rect 31401 10081 31435 10115
rect 33701 10081 33735 10115
rect 15209 10013 15243 10047
rect 15393 10013 15427 10047
rect 15485 10013 15519 10047
rect 16129 10013 16163 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 18613 10013 18647 10047
rect 19349 10013 19383 10047
rect 19809 10013 19843 10047
rect 19993 10013 20027 10047
rect 22569 10013 22603 10047
rect 27261 10013 27295 10047
rect 29653 10013 29687 10047
rect 29929 10013 29963 10047
rect 30205 10013 30239 10047
rect 30297 10013 30331 10047
rect 30481 10013 30515 10047
rect 30757 10013 30791 10047
rect 31677 10013 31711 10047
rect 31861 10013 31895 10047
rect 32045 10013 32079 10047
rect 32229 10013 32263 10047
rect 32505 10013 32539 10047
rect 32689 10013 32723 10047
rect 33977 10013 34011 10047
rect 34713 10013 34747 10047
rect 34805 10013 34839 10047
rect 35357 10013 35391 10047
rect 35541 10013 35575 10047
rect 14749 9945 14783 9979
rect 30113 9945 30147 9979
rect 33885 9945 33919 9979
rect 29837 9877 29871 9911
rect 31585 9877 31619 9911
rect 34069 9877 34103 9911
rect 34253 9877 34287 9911
rect 15393 9673 15427 9707
rect 18245 9673 18279 9707
rect 26157 9673 26191 9707
rect 28733 9673 28767 9707
rect 33793 9673 33827 9707
rect 13921 9605 13955 9639
rect 18153 9605 18187 9639
rect 19717 9605 19751 9639
rect 23305 9605 23339 9639
rect 26525 9605 26559 9639
rect 26709 9605 26743 9639
rect 27261 9605 27295 9639
rect 29285 9605 29319 9639
rect 31769 9605 31803 9639
rect 32321 9605 32355 9639
rect 33425 9605 33459 9639
rect 34405 9605 34439 9639
rect 34621 9605 34655 9639
rect 13645 9537 13679 9571
rect 16497 9537 16531 9571
rect 17417 9537 17451 9571
rect 17509 9537 17543 9571
rect 17693 9537 17727 9571
rect 21281 9537 21315 9571
rect 23581 9537 23615 9571
rect 23673 9537 23707 9571
rect 24409 9537 24443 9571
rect 29193 9537 29227 9571
rect 29837 9537 29871 9571
rect 30021 9537 30055 9571
rect 30297 9537 30331 9571
rect 30849 9537 30883 9571
rect 31125 9537 31159 9571
rect 32505 9537 32539 9571
rect 32689 9537 32723 9571
rect 33701 9537 33735 9571
rect 33977 9537 34011 9571
rect 34713 9537 34747 9571
rect 34989 9537 35023 9571
rect 15669 9469 15703 9503
rect 19993 9469 20027 9503
rect 20269 9469 20303 9503
rect 21833 9469 21867 9503
rect 24685 9469 24719 9503
rect 26985 9469 27019 9503
rect 29469 9469 29503 9503
rect 29653 9469 29687 9503
rect 30665 9469 30699 9503
rect 34161 9469 34195 9503
rect 28825 9333 28859 9367
rect 34253 9333 34287 9367
rect 34437 9333 34471 9367
rect 34805 9333 34839 9367
rect 23673 9129 23707 9163
rect 25513 9129 25547 9163
rect 28733 9129 28767 9163
rect 29193 9129 29227 9163
rect 29377 9129 29411 9163
rect 31217 9129 31251 9163
rect 31953 9129 31987 9163
rect 33535 9129 33569 9163
rect 16037 8993 16071 9027
rect 19717 8993 19751 9027
rect 21925 8993 21959 9027
rect 22201 8993 22235 9027
rect 26065 8993 26099 9027
rect 26985 8993 27019 9027
rect 27261 8993 27295 9027
rect 29745 8993 29779 9027
rect 31309 8993 31343 9027
rect 31677 8993 31711 9027
rect 31769 8993 31803 9027
rect 32045 8993 32079 9027
rect 33793 8993 33827 9027
rect 34713 8993 34747 9027
rect 15209 8925 15243 8959
rect 15393 8925 15427 8959
rect 15485 8925 15519 8959
rect 18337 8925 18371 8959
rect 18521 8925 18555 8959
rect 18613 8925 18647 8959
rect 21465 8925 21499 8959
rect 24869 8925 24903 8959
rect 25053 8925 25087 8959
rect 25145 8925 25179 8959
rect 25881 8925 25915 8959
rect 26893 8925 26927 8959
rect 30389 8925 30423 8959
rect 31033 8925 31067 8959
rect 31539 8925 31573 8959
rect 34253 8925 34287 8959
rect 34897 8925 34931 8959
rect 34989 8925 35023 8959
rect 14749 8857 14783 8891
rect 16313 8857 16347 8891
rect 17877 8857 17911 8891
rect 21189 8857 21223 8891
rect 24409 8857 24443 8891
rect 29009 8857 29043 8891
rect 30665 8857 30699 8891
rect 30941 8857 30975 8891
rect 31401 8857 31435 8891
rect 33885 8857 33919 8891
rect 34437 8857 34471 8891
rect 17785 8789 17819 8823
rect 25973 8789 26007 8823
rect 29219 8789 29253 8823
rect 30849 8789 30883 8823
rect 34713 8789 34747 8823
rect 15577 8585 15611 8619
rect 35633 8585 35667 8619
rect 14105 8517 14139 8551
rect 17601 8517 17635 8551
rect 23029 8517 23063 8551
rect 25605 8517 25639 8551
rect 27169 8517 27203 8551
rect 27629 8517 27663 8551
rect 28457 8517 28491 8551
rect 29009 8517 29043 8551
rect 29837 8517 29871 8551
rect 31553 8517 31587 8551
rect 31769 8517 31803 8551
rect 33057 8517 33091 8551
rect 33977 8517 34011 8551
rect 18521 8449 18555 8483
rect 18705 8449 18739 8483
rect 20453 8449 20487 8483
rect 20545 8449 20579 8483
rect 20729 8449 20763 8483
rect 21189 8449 21223 8483
rect 23765 8449 23799 8483
rect 23949 8449 23983 8483
rect 26801 8449 26835 8483
rect 26985 8449 27019 8483
rect 28917 8449 28951 8483
rect 33149 8449 33183 8483
rect 33333 8449 33367 8483
rect 33425 8449 33459 8483
rect 33701 8449 33735 8483
rect 35541 8449 35575 8483
rect 13829 8381 13863 8415
rect 16773 8381 16807 8415
rect 18420 8381 18454 8415
rect 19165 8381 19199 8415
rect 22201 8381 22235 8415
rect 23673 8381 23707 8415
rect 24409 8381 24443 8415
rect 29193 8381 29227 8415
rect 29561 8381 29595 8415
rect 32229 8381 32263 8415
rect 35449 8381 35483 8415
rect 31309 8313 31343 8347
rect 31401 8313 31435 8347
rect 33149 8313 33183 8347
rect 28549 8245 28583 8279
rect 31585 8245 31619 8279
rect 17325 8041 17359 8075
rect 26157 8041 26191 8075
rect 34989 8041 35023 8075
rect 23397 7973 23431 8007
rect 14289 7905 14323 7939
rect 18797 7905 18831 7939
rect 21465 7905 21499 7939
rect 21557 7905 21591 7939
rect 21833 7905 21867 7939
rect 23857 7905 23891 7939
rect 23949 7905 23983 7939
rect 28273 7905 28307 7939
rect 30205 7905 30239 7939
rect 30665 7905 30699 7939
rect 17233 7837 17267 7871
rect 19073 7837 19107 7871
rect 24409 7837 24443 7871
rect 29929 7837 29963 7871
rect 31769 7837 31803 7871
rect 32873 7837 32907 7871
rect 34069 7837 34103 7871
rect 34713 7837 34747 7871
rect 35357 7837 35391 7871
rect 35817 7837 35851 7871
rect 14565 7769 14599 7803
rect 21189 7769 21223 7803
rect 23765 7769 23799 7803
rect 24685 7769 24719 7803
rect 27997 7769 28031 7803
rect 32045 7769 32079 7803
rect 32965 7769 32999 7803
rect 36185 7769 36219 7803
rect 16037 7701 16071 7735
rect 19717 7701 19751 7735
rect 23305 7701 23339 7735
rect 26525 7701 26559 7735
rect 29561 7701 29595 7735
rect 30021 7701 30055 7735
rect 34253 7701 34287 7735
rect 22477 7497 22511 7531
rect 26065 7497 26099 7531
rect 27445 7497 27479 7531
rect 29929 7497 29963 7531
rect 15025 7429 15059 7463
rect 23949 7429 23983 7463
rect 24593 7429 24627 7463
rect 27353 7429 27387 7463
rect 28457 7429 28491 7463
rect 31677 7429 31711 7463
rect 31861 7429 31895 7463
rect 34161 7429 34195 7463
rect 34897 7429 34931 7463
rect 35265 7429 35299 7463
rect 15485 7361 15519 7395
rect 15669 7361 15703 7395
rect 15761 7361 15795 7395
rect 21189 7361 21223 7395
rect 28181 7361 28215 7395
rect 30297 7361 30331 7395
rect 31217 7361 31251 7395
rect 32137 7361 32171 7395
rect 34345 7361 34379 7395
rect 16681 7293 16715 7327
rect 16957 7293 16991 7327
rect 20913 7293 20947 7327
rect 24225 7293 24259 7327
rect 24317 7293 24351 7327
rect 27537 7293 27571 7327
rect 30021 7293 30055 7327
rect 32413 7293 32447 7327
rect 31401 7225 31435 7259
rect 35081 7225 35115 7259
rect 18429 7157 18463 7191
rect 19441 7157 19475 7191
rect 26985 7157 27019 7191
rect 22201 6953 22235 6987
rect 26328 6953 26362 6987
rect 27813 6953 27847 6987
rect 31125 6953 31159 6987
rect 34069 6953 34103 6987
rect 34345 6953 34379 6987
rect 30389 6885 30423 6919
rect 34161 6885 34195 6919
rect 16681 6817 16715 6851
rect 22845 6817 22879 6851
rect 24961 6817 24995 6851
rect 25697 6817 25731 6851
rect 30481 6817 30515 6851
rect 31493 6817 31527 6851
rect 32321 6817 32355 6851
rect 15393 6749 15427 6783
rect 15577 6749 15611 6783
rect 15669 6749 15703 6783
rect 19257 6749 19291 6783
rect 21005 6749 21039 6783
rect 21557 6749 21591 6783
rect 21741 6749 21775 6783
rect 21833 6749 21867 6783
rect 22661 6749 22695 6783
rect 25421 6749 25455 6783
rect 25605 6749 25639 6783
rect 26065 6749 26099 6783
rect 30941 6749 30975 6783
rect 31125 6749 31159 6783
rect 31401 6749 31435 6783
rect 31585 6749 31619 6783
rect 34713 6749 34747 6783
rect 34989 6749 35023 6783
rect 35357 6749 35391 6783
rect 14933 6681 14967 6715
rect 16957 6681 16991 6715
rect 21097 6681 21131 6715
rect 30021 6681 30055 6715
rect 32597 6681 32631 6715
rect 34529 6681 34563 6715
rect 18429 6613 18463 6647
rect 22569 6613 22603 6647
rect 34329 6613 34363 6647
rect 34805 6613 34839 6647
rect 35173 6613 35207 6647
rect 33885 6409 33919 6443
rect 17325 6341 17359 6375
rect 21189 6341 21223 6375
rect 27537 6341 27571 6375
rect 32781 6341 32815 6375
rect 33517 6341 33551 6375
rect 33733 6341 33767 6375
rect 34253 6341 34287 6375
rect 13829 6273 13863 6307
rect 17785 6273 17819 6307
rect 17969 6273 18003 6307
rect 18061 6273 18095 6307
rect 18521 6273 18555 6307
rect 18981 6273 19015 6307
rect 19165 6273 19199 6307
rect 19257 6273 19291 6307
rect 20453 6273 20487 6307
rect 20545 6273 20579 6307
rect 20729 6273 20763 6307
rect 22201 6273 22235 6307
rect 33149 6273 33183 6307
rect 33333 6273 33367 6307
rect 14105 6205 14139 6239
rect 22293 6205 22327 6239
rect 22477 6205 22511 6239
rect 23397 6205 23431 6239
rect 23673 6205 23707 6239
rect 27629 6205 27663 6239
rect 27813 6205 27847 6239
rect 28181 6205 28215 6239
rect 28457 6205 28491 6239
rect 30205 6205 30239 6239
rect 30481 6205 30515 6239
rect 31953 6205 31987 6239
rect 32689 6205 32723 6239
rect 33977 6205 34011 6239
rect 36737 6137 36771 6171
rect 15577 6069 15611 6103
rect 21833 6069 21867 6103
rect 25145 6069 25179 6103
rect 27169 6069 27203 6103
rect 29929 6069 29963 6103
rect 32229 6069 32263 6103
rect 33701 6069 33735 6103
rect 35725 6069 35759 6103
rect 21005 5865 21039 5899
rect 25960 5865 25994 5899
rect 27537 5865 27571 5899
rect 30205 5865 30239 5899
rect 33609 5865 33643 5899
rect 27445 5797 27479 5831
rect 15117 5729 15151 5763
rect 16589 5729 16623 5763
rect 19257 5729 19291 5763
rect 19533 5729 19567 5763
rect 21373 5729 21407 5763
rect 23949 5729 23983 5763
rect 24409 5729 24443 5763
rect 25145 5729 25179 5763
rect 27997 5729 28031 5763
rect 28181 5729 28215 5763
rect 30665 5729 30699 5763
rect 30849 5729 30883 5763
rect 31033 5729 31067 5763
rect 33149 5729 33183 5763
rect 33333 5729 33367 5763
rect 34713 5729 34747 5763
rect 14841 5661 14875 5695
rect 15025 5661 15059 5695
rect 15945 5661 15979 5695
rect 16129 5661 16163 5695
rect 16221 5661 16255 5695
rect 23121 5661 23155 5695
rect 23673 5661 23707 5695
rect 23857 5661 23891 5695
rect 24869 5661 24903 5695
rect 25053 5661 25087 5695
rect 25697 5661 25731 5695
rect 27905 5661 27939 5695
rect 28457 5661 28491 5695
rect 28549 5661 28583 5695
rect 31309 5661 31343 5695
rect 33241 5661 33275 5695
rect 33425 5661 33459 5695
rect 33701 5661 33735 5695
rect 33977 5661 34011 5695
rect 14381 5593 14415 5627
rect 15485 5593 15519 5627
rect 16865 5593 16899 5627
rect 22845 5593 22879 5627
rect 23213 5593 23247 5627
rect 34897 5593 34931 5627
rect 18337 5525 18371 5559
rect 28733 5525 28767 5559
rect 30573 5525 30607 5559
rect 15853 5321 15887 5355
rect 28733 5321 28767 5355
rect 30205 5321 30239 5355
rect 32305 5321 32339 5355
rect 14381 5253 14415 5287
rect 16957 5253 16991 5287
rect 23305 5253 23339 5287
rect 27261 5253 27295 5287
rect 29837 5253 29871 5287
rect 29929 5253 29963 5287
rect 30389 5253 30423 5287
rect 32505 5253 32539 5287
rect 34253 5253 34287 5287
rect 35081 5253 35115 5287
rect 14105 5185 14139 5219
rect 17417 5185 17451 5219
rect 17601 5185 17635 5219
rect 17693 5185 17727 5219
rect 18981 5185 19015 5219
rect 23581 5185 23615 5219
rect 25421 5185 25455 5219
rect 26985 5185 27019 5219
rect 29561 5185 29595 5219
rect 29654 5185 29688 5219
rect 30067 5185 30101 5219
rect 30297 5185 30331 5219
rect 30481 5185 30515 5219
rect 30849 5185 30883 5219
rect 31033 5185 31067 5219
rect 31125 5185 31159 5219
rect 31401 5185 31435 5219
rect 31493 5185 31527 5219
rect 32965 5185 32999 5219
rect 33149 5185 33183 5219
rect 33425 5185 33459 5219
rect 34161 5185 34195 5219
rect 34713 5185 34747 5219
rect 34897 5185 34931 5219
rect 35173 5185 35207 5219
rect 19257 5117 19291 5151
rect 21833 5117 21867 5151
rect 25145 5117 25179 5151
rect 30665 5117 30699 5151
rect 34069 5117 34103 5151
rect 34805 5117 34839 5151
rect 20729 5049 20763 5083
rect 32137 5049 32171 5083
rect 23673 4981 23707 5015
rect 31217 4981 31251 5015
rect 32321 4981 32355 5015
rect 35173 4981 35207 5015
rect 17049 4777 17083 4811
rect 35265 4777 35299 4811
rect 35541 4777 35575 4811
rect 34069 4709 34103 4743
rect 15301 4641 15335 4675
rect 15577 4641 15611 4675
rect 20821 4641 20855 4675
rect 24409 4641 24443 4675
rect 25145 4641 25179 4675
rect 31585 4641 31619 4675
rect 31861 4641 31895 4675
rect 32597 4641 32631 4675
rect 34989 4641 35023 4675
rect 35081 4641 35115 4675
rect 21281 4573 21315 4607
rect 21465 4573 21499 4607
rect 21557 4573 21591 4607
rect 24869 4573 24903 4607
rect 25053 4573 25087 4607
rect 30113 4573 30147 4607
rect 30297 4573 30331 4607
rect 30389 4573 30423 4607
rect 32137 4573 32171 4607
rect 32229 4573 32263 4607
rect 33241 4573 33275 4607
rect 33517 4573 33551 4607
rect 33609 4573 33643 4607
rect 34805 4573 34839 4607
rect 34897 4573 34931 4607
rect 29653 4505 29687 4539
rect 35525 4505 35559 4539
rect 35725 4505 35759 4539
rect 31953 4437 31987 4471
rect 32321 4437 32355 4471
rect 32505 4437 32539 4471
rect 35357 4437 35391 4471
rect 30389 4233 30423 4267
rect 31109 4233 31143 4267
rect 31861 4233 31895 4267
rect 32229 4233 32263 4267
rect 33333 4233 33367 4267
rect 33609 4233 33643 4267
rect 31309 4165 31343 4199
rect 33057 4165 33091 4199
rect 33149 4165 33183 4199
rect 35081 4165 35115 4199
rect 28457 4097 28491 4131
rect 32781 4097 32815 4131
rect 32965 4097 32999 4131
rect 28733 4029 28767 4063
rect 30205 4029 30239 4063
rect 30849 4029 30883 4063
rect 31401 4029 31435 4063
rect 32689 4029 32723 4063
rect 35357 4029 35391 4063
rect 30941 3893 30975 3927
rect 31125 3893 31159 3927
rect 32505 3689 32539 3723
rect 30297 3553 30331 3587
rect 31769 3553 31803 3587
rect 32689 3553 32723 3587
rect 33885 3553 33919 3587
rect 30021 3485 30055 3519
rect 32137 3485 32171 3519
rect 32413 3485 32447 3519
rect 32597 3485 32631 3519
rect 33149 3485 33183 3519
rect 33333 3485 33367 3519
rect 33425 3485 33459 3519
rect 33793 3485 33827 3519
rect 33977 3485 34011 3519
rect 32045 3349 32079 3383
rect 33885 3145 33919 3179
rect 30481 3077 30515 3111
rect 32413 3077 32447 3111
rect 30205 2941 30239 2975
rect 31953 2941 31987 2975
rect 32137 2941 32171 2975
rect 23489 2601 23523 2635
rect 23305 2397 23339 2431
<< metal1 >>
rect 1104 38106 37076 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 37076 38106
rect 1104 38032 37076 38054
rect 31938 37884 31944 37936
rect 31996 37924 32002 37936
rect 32125 37927 32183 37933
rect 32125 37924 32137 37927
rect 31996 37896 32137 37924
rect 31996 37884 32002 37896
rect 32125 37893 32137 37896
rect 32171 37893 32183 37927
rect 32125 37887 32183 37893
rect 32341 37927 32399 37933
rect 32341 37893 32353 37927
rect 32387 37924 32399 37927
rect 32950 37924 32956 37936
rect 32387 37896 32956 37924
rect 32387 37893 32399 37896
rect 32341 37887 32399 37893
rect 32950 37884 32956 37896
rect 33008 37884 33014 37936
rect 12526 37816 12532 37868
rect 12584 37856 12590 37868
rect 13541 37859 13599 37865
rect 13541 37856 13553 37859
rect 12584 37828 13553 37856
rect 12584 37816 12590 37828
rect 13541 37825 13553 37828
rect 13587 37825 13599 37859
rect 13541 37819 13599 37825
rect 16022 37816 16028 37868
rect 16080 37816 16086 37868
rect 16117 37859 16175 37865
rect 16117 37825 16129 37859
rect 16163 37856 16175 37859
rect 16390 37856 16396 37868
rect 16163 37828 16396 37856
rect 16163 37825 16175 37828
rect 16117 37819 16175 37825
rect 16390 37816 16396 37828
rect 16448 37816 16454 37868
rect 18598 37816 18604 37868
rect 18656 37816 18662 37868
rect 23569 37859 23627 37865
rect 23569 37825 23581 37859
rect 23615 37856 23627 37859
rect 23842 37856 23848 37868
rect 23615 37828 23848 37856
rect 23615 37825 23627 37828
rect 23569 37819 23627 37825
rect 23842 37816 23848 37828
rect 23900 37816 23906 37868
rect 25222 37816 25228 37868
rect 25280 37816 25286 37868
rect 27433 37859 27491 37865
rect 27433 37825 27445 37859
rect 27479 37856 27491 37859
rect 28074 37856 28080 37868
rect 27479 37828 28080 37856
rect 27479 37825 27491 37828
rect 27433 37819 27491 37825
rect 28074 37816 28080 37828
rect 28132 37816 28138 37868
rect 29730 37816 29736 37868
rect 29788 37816 29794 37868
rect 30745 37859 30803 37865
rect 30745 37825 30757 37859
rect 30791 37856 30803 37859
rect 31662 37856 31668 37868
rect 30791 37828 31668 37856
rect 30791 37825 30803 37828
rect 30745 37819 30803 37825
rect 31662 37816 31668 37828
rect 31720 37816 31726 37868
rect 31757 37859 31815 37865
rect 31757 37825 31769 37859
rect 31803 37856 31815 37859
rect 32858 37856 32864 37868
rect 31803 37828 32864 37856
rect 31803 37825 31815 37828
rect 31757 37819 31815 37825
rect 32858 37816 32864 37828
rect 32916 37816 32922 37868
rect 13078 37748 13084 37800
rect 13136 37788 13142 37800
rect 13633 37791 13691 37797
rect 13633 37788 13645 37791
rect 13136 37760 13645 37788
rect 13136 37748 13142 37760
rect 13633 37757 13645 37760
rect 13679 37757 13691 37791
rect 13633 37751 13691 37757
rect 13722 37748 13728 37800
rect 13780 37748 13786 37800
rect 16301 37791 16359 37797
rect 16301 37757 16313 37791
rect 16347 37757 16359 37791
rect 16301 37751 16359 37757
rect 16316 37720 16344 37751
rect 18690 37748 18696 37800
rect 18748 37748 18754 37800
rect 18874 37748 18880 37800
rect 18932 37748 18938 37800
rect 23658 37748 23664 37800
rect 23716 37748 23722 37800
rect 23753 37791 23811 37797
rect 23753 37757 23765 37791
rect 23799 37788 23811 37791
rect 24854 37788 24860 37800
rect 23799 37760 24860 37788
rect 23799 37757 23811 37760
rect 23753 37751 23811 37757
rect 24854 37748 24860 37760
rect 24912 37748 24918 37800
rect 27246 37748 27252 37800
rect 27304 37788 27310 37800
rect 27525 37791 27583 37797
rect 27525 37788 27537 37791
rect 27304 37760 27537 37788
rect 27304 37748 27310 37760
rect 27525 37757 27537 37760
rect 27571 37757 27583 37791
rect 27525 37751 27583 37757
rect 29178 37748 29184 37800
rect 29236 37748 29242 37800
rect 30009 37791 30067 37797
rect 30009 37757 30021 37791
rect 30055 37788 30067 37791
rect 30374 37788 30380 37800
rect 30055 37760 30380 37788
rect 30055 37757 30067 37760
rect 30009 37751 30067 37757
rect 30374 37748 30380 37760
rect 30432 37748 30438 37800
rect 30929 37791 30987 37797
rect 30929 37757 30941 37791
rect 30975 37788 30987 37791
rect 31481 37791 31539 37797
rect 31481 37788 31493 37791
rect 30975 37760 31493 37788
rect 30975 37757 30987 37760
rect 30929 37751 30987 37757
rect 31481 37757 31493 37760
rect 31527 37788 31539 37791
rect 31846 37788 31852 37800
rect 31527 37760 31852 37788
rect 31527 37757 31539 37760
rect 31481 37751 31539 37757
rect 31846 37748 31852 37760
rect 31904 37748 31910 37800
rect 18892 37720 18920 37748
rect 16316 37692 18920 37720
rect 31665 37723 31723 37729
rect 31665 37689 31677 37723
rect 31711 37720 31723 37723
rect 32214 37720 32220 37732
rect 31711 37692 32220 37720
rect 31711 37689 31723 37692
rect 31665 37683 31723 37689
rect 32214 37680 32220 37692
rect 32272 37680 32278 37732
rect 13173 37655 13231 37661
rect 13173 37621 13185 37655
rect 13219 37652 13231 37655
rect 13446 37652 13452 37664
rect 13219 37624 13452 37652
rect 13219 37621 13231 37624
rect 13173 37615 13231 37621
rect 13446 37612 13452 37624
rect 13504 37612 13510 37664
rect 15657 37655 15715 37661
rect 15657 37621 15669 37655
rect 15703 37652 15715 37655
rect 16206 37652 16212 37664
rect 15703 37624 16212 37652
rect 15703 37621 15715 37624
rect 15657 37615 15715 37621
rect 16206 37612 16212 37624
rect 16264 37612 16270 37664
rect 17494 37612 17500 37664
rect 17552 37652 17558 37664
rect 18233 37655 18291 37661
rect 18233 37652 18245 37655
rect 17552 37624 18245 37652
rect 17552 37612 17558 37624
rect 18233 37621 18245 37624
rect 18279 37621 18291 37655
rect 18233 37615 18291 37621
rect 22370 37612 22376 37664
rect 22428 37652 22434 37664
rect 23201 37655 23259 37661
rect 23201 37652 23213 37655
rect 22428 37624 23213 37652
rect 22428 37612 22434 37624
rect 23201 37621 23213 37624
rect 23247 37621 23259 37655
rect 23201 37615 23259 37621
rect 25406 37612 25412 37664
rect 25464 37612 25470 37664
rect 27249 37655 27307 37661
rect 27249 37621 27261 37655
rect 27295 37652 27307 37655
rect 27706 37652 27712 37664
rect 27295 37624 27712 37652
rect 27295 37621 27307 37624
rect 27249 37615 27307 37621
rect 27706 37612 27712 37624
rect 27764 37612 27770 37664
rect 27982 37612 27988 37664
rect 28040 37652 28046 37664
rect 28721 37655 28779 37661
rect 28721 37652 28733 37655
rect 28040 37624 28733 37652
rect 28040 37612 28046 37624
rect 28721 37621 28733 37624
rect 28767 37621 28779 37655
rect 28721 37615 28779 37621
rect 31570 37612 31576 37664
rect 31628 37612 31634 37664
rect 32306 37612 32312 37664
rect 32364 37612 32370 37664
rect 32490 37612 32496 37664
rect 32548 37612 32554 37664
rect 1104 37562 37076 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 37076 37562
rect 1104 37488 37076 37510
rect 14737 37451 14795 37457
rect 14737 37417 14749 37451
rect 14783 37448 14795 37451
rect 15470 37448 15476 37460
rect 14783 37420 15476 37448
rect 14783 37417 14795 37420
rect 14737 37411 14795 37417
rect 15470 37408 15476 37420
rect 15528 37448 15534 37460
rect 16022 37448 16028 37460
rect 15528 37420 16028 37448
rect 15528 37408 15534 37420
rect 16022 37408 16028 37420
rect 16080 37408 16086 37460
rect 18598 37408 18604 37460
rect 18656 37448 18662 37460
rect 18969 37451 19027 37457
rect 18969 37448 18981 37451
rect 18656 37420 18981 37448
rect 18656 37408 18662 37420
rect 18969 37417 18981 37420
rect 19015 37417 19027 37451
rect 18969 37411 19027 37417
rect 23658 37408 23664 37460
rect 23716 37448 23722 37460
rect 24394 37448 24400 37460
rect 23716 37420 24400 37448
rect 23716 37408 23722 37420
rect 24394 37408 24400 37420
rect 24452 37408 24458 37460
rect 28074 37408 28080 37460
rect 28132 37408 28138 37460
rect 31573 37451 31631 37457
rect 31573 37417 31585 37451
rect 31619 37448 31631 37451
rect 31938 37448 31944 37460
rect 31619 37420 31944 37448
rect 31619 37417 31631 37420
rect 31573 37411 31631 37417
rect 31938 37408 31944 37420
rect 31996 37408 32002 37460
rect 23842 37340 23848 37392
rect 23900 37340 23906 37392
rect 13446 37272 13452 37324
rect 13504 37272 13510 37324
rect 16206 37272 16212 37324
rect 16264 37272 16270 37324
rect 17494 37272 17500 37324
rect 17552 37272 17558 37324
rect 19429 37315 19487 37321
rect 19429 37281 19441 37315
rect 19475 37312 19487 37315
rect 21542 37312 21548 37324
rect 19475 37284 21548 37312
rect 19475 37281 19487 37284
rect 19429 37275 19487 37281
rect 21542 37272 21548 37284
rect 21600 37272 21606 37324
rect 22370 37272 22376 37324
rect 22428 37272 22434 37324
rect 30101 37315 30159 37321
rect 27540 37284 27752 37312
rect 27540 37256 27568 37284
rect 842 37204 848 37256
rect 900 37244 906 37256
rect 1397 37247 1455 37253
rect 1397 37244 1409 37247
rect 900 37216 1409 37244
rect 900 37204 906 37216
rect 1397 37213 1409 37216
rect 1443 37213 1455 37247
rect 1397 37207 1455 37213
rect 13725 37247 13783 37253
rect 13725 37213 13737 37247
rect 13771 37244 13783 37247
rect 14642 37244 14648 37256
rect 13771 37216 14648 37244
rect 13771 37213 13783 37216
rect 13725 37207 13783 37213
rect 14642 37204 14648 37216
rect 14700 37204 14706 37256
rect 16485 37247 16543 37253
rect 16485 37213 16497 37247
rect 16531 37244 16543 37247
rect 17221 37247 17279 37253
rect 17221 37244 17233 37247
rect 16531 37216 17233 37244
rect 16531 37213 16543 37216
rect 16485 37207 16543 37213
rect 17221 37213 17233 37216
rect 17267 37213 17279 37247
rect 17221 37207 17279 37213
rect 21821 37247 21879 37253
rect 21821 37213 21833 37247
rect 21867 37244 21879 37247
rect 22097 37247 22155 37253
rect 22097 37244 22109 37247
rect 21867 37216 22109 37244
rect 21867 37213 21879 37216
rect 21821 37207 21879 37213
rect 22097 37213 22109 37216
rect 22143 37213 22155 37247
rect 22097 37207 22155 37213
rect 2593 37179 2651 37185
rect 2593 37145 2605 37179
rect 2639 37176 2651 37179
rect 3326 37176 3332 37188
rect 2639 37148 3332 37176
rect 2639 37145 2651 37148
rect 2593 37139 2651 37145
rect 3326 37136 3332 37148
rect 3384 37136 3390 37188
rect 12986 37136 12992 37188
rect 13044 37136 13050 37188
rect 15562 37136 15568 37188
rect 15620 37136 15626 37188
rect 16500 37120 16528 37207
rect 19426 37176 19432 37188
rect 18722 37148 19432 37176
rect 19426 37136 19432 37148
rect 19484 37136 19490 37188
rect 19521 37179 19579 37185
rect 19521 37145 19533 37179
rect 19567 37176 19579 37179
rect 21266 37176 21272 37188
rect 19567 37148 20116 37176
rect 21114 37148 21272 37176
rect 19567 37145 19579 37148
rect 19521 37139 19579 37145
rect 20088 37120 20116 37148
rect 21266 37136 21272 37148
rect 21324 37136 21330 37188
rect 21450 37136 21456 37188
rect 21508 37176 21514 37188
rect 21545 37179 21603 37185
rect 21545 37176 21557 37179
rect 21508 37148 21557 37176
rect 21508 37136 21514 37148
rect 21545 37145 21557 37148
rect 21591 37145 21603 37179
rect 21545 37139 21603 37145
rect 11977 37111 12035 37117
rect 11977 37077 11989 37111
rect 12023 37108 12035 37111
rect 12526 37108 12532 37120
rect 12023 37080 12532 37108
rect 12023 37077 12035 37080
rect 11977 37071 12035 37077
rect 12526 37068 12532 37080
rect 12584 37068 12590 37120
rect 15194 37068 15200 37120
rect 15252 37108 15258 37120
rect 16482 37108 16488 37120
rect 15252 37080 16488 37108
rect 15252 37068 15258 37080
rect 16482 37068 16488 37080
rect 16540 37068 16546 37120
rect 18782 37068 18788 37120
rect 18840 37108 18846 37120
rect 19613 37111 19671 37117
rect 19613 37108 19625 37111
rect 18840 37080 19625 37108
rect 18840 37068 18846 37080
rect 19613 37077 19625 37080
rect 19659 37077 19671 37111
rect 19613 37071 19671 37077
rect 19886 37068 19892 37120
rect 19944 37108 19950 37120
rect 19981 37111 20039 37117
rect 19981 37108 19993 37111
rect 19944 37080 19993 37108
rect 19944 37068 19950 37080
rect 19981 37077 19993 37080
rect 20027 37077 20039 37111
rect 19981 37071 20039 37077
rect 20070 37068 20076 37120
rect 20128 37068 20134 37120
rect 20530 37068 20536 37120
rect 20588 37108 20594 37120
rect 21836 37108 21864 37207
rect 26142 37204 26148 37256
rect 26200 37244 26206 37256
rect 26237 37247 26295 37253
rect 26237 37244 26249 37247
rect 26200 37216 26249 37244
rect 26200 37204 26206 37216
rect 26237 37213 26249 37216
rect 26283 37213 26295 37247
rect 26237 37207 26295 37213
rect 27522 37204 27528 37256
rect 27580 37204 27586 37256
rect 27724 37244 27752 37284
rect 30101 37281 30113 37315
rect 30147 37312 30159 37315
rect 30466 37312 30472 37324
rect 30147 37284 30472 37312
rect 30147 37281 30159 37284
rect 30101 37275 30159 37281
rect 30466 37272 30472 37284
rect 30524 37272 30530 37324
rect 30558 37272 30564 37324
rect 30616 37312 30622 37324
rect 30616 37284 33088 37312
rect 30616 37272 30622 37284
rect 28261 37247 28319 37253
rect 28261 37244 28273 37247
rect 27724 37216 28273 37244
rect 28261 37213 28273 37216
rect 28307 37213 28319 37247
rect 28261 37207 28319 37213
rect 28534 37204 28540 37256
rect 28592 37204 28598 37256
rect 28718 37204 28724 37256
rect 28776 37204 28782 37256
rect 29822 37204 29828 37256
rect 29880 37204 29886 37256
rect 31665 37247 31723 37253
rect 31665 37244 31677 37247
rect 31496 37216 31677 37244
rect 22278 37136 22284 37188
rect 22336 37176 22342 37188
rect 22336 37148 22862 37176
rect 24412 37148 24702 37176
rect 22336 37136 22342 37148
rect 22002 37108 22008 37120
rect 20588 37080 22008 37108
rect 20588 37068 20594 37080
rect 22002 37068 22008 37080
rect 22060 37068 22066 37120
rect 22756 37108 22784 37148
rect 24412 37108 24440 37148
rect 25866 37136 25872 37188
rect 25924 37136 25930 37188
rect 26510 37136 26516 37188
rect 26568 37136 26574 37188
rect 28902 37176 28908 37188
rect 27738 37148 28908 37176
rect 28902 37136 28908 37148
rect 28960 37136 28966 37188
rect 29273 37179 29331 37185
rect 29273 37145 29285 37179
rect 29319 37176 29331 37179
rect 29730 37176 29736 37188
rect 29319 37148 29736 37176
rect 29319 37145 29331 37148
rect 29273 37139 29331 37145
rect 29730 37136 29736 37148
rect 29788 37136 29794 37188
rect 30558 37136 30564 37188
rect 30616 37136 30622 37188
rect 31496 37120 31524 37216
rect 31665 37213 31677 37216
rect 31711 37213 31723 37247
rect 33060 37244 33088 37284
rect 33962 37244 33968 37256
rect 33060 37230 33968 37244
rect 33074 37216 33968 37230
rect 31665 37207 31723 37213
rect 33962 37204 33968 37216
rect 34020 37204 34026 37256
rect 31570 37136 31576 37188
rect 31628 37176 31634 37188
rect 31941 37179 31999 37185
rect 31941 37176 31953 37179
rect 31628 37148 31953 37176
rect 31628 37136 31634 37148
rect 31941 37145 31953 37148
rect 31987 37145 31999 37179
rect 31941 37139 31999 37145
rect 22756 37080 24440 37108
rect 26602 37068 26608 37120
rect 26660 37108 26666 37120
rect 27985 37111 28043 37117
rect 27985 37108 27997 37111
rect 26660 37080 27997 37108
rect 26660 37068 26666 37080
rect 27985 37077 27997 37080
rect 28031 37077 28043 37111
rect 27985 37071 28043 37077
rect 28258 37068 28264 37120
rect 28316 37108 28322 37120
rect 28445 37111 28503 37117
rect 28445 37108 28457 37111
rect 28316 37080 28457 37108
rect 28316 37068 28322 37080
rect 28445 37077 28457 37080
rect 28491 37077 28503 37111
rect 28445 37071 28503 37077
rect 29822 37068 29828 37120
rect 29880 37108 29886 37120
rect 31478 37108 31484 37120
rect 29880 37080 31484 37108
rect 29880 37068 29886 37080
rect 31478 37068 31484 37080
rect 31536 37108 31542 37120
rect 33226 37108 33232 37120
rect 31536 37080 33232 37108
rect 31536 37068 31542 37080
rect 33226 37068 33232 37080
rect 33284 37068 33290 37120
rect 33410 37068 33416 37120
rect 33468 37068 33474 37120
rect 1104 37018 37076 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 37076 37018
rect 1104 36944 37076 36966
rect 12526 36864 12532 36916
rect 12584 36864 12590 36916
rect 16390 36864 16396 36916
rect 16448 36904 16454 36916
rect 16485 36907 16543 36913
rect 16485 36904 16497 36907
rect 16448 36876 16497 36904
rect 16448 36864 16454 36876
rect 16485 36873 16497 36876
rect 16531 36904 16543 36907
rect 17037 36907 17095 36913
rect 17037 36904 17049 36907
rect 16531 36876 17049 36904
rect 16531 36873 16543 36876
rect 16485 36867 16543 36873
rect 17037 36873 17049 36876
rect 17083 36873 17095 36907
rect 17037 36867 17095 36873
rect 18417 36907 18475 36913
rect 18417 36873 18429 36907
rect 18463 36904 18475 36907
rect 18598 36904 18604 36916
rect 18463 36876 18604 36904
rect 18463 36873 18475 36876
rect 18417 36867 18475 36873
rect 18598 36864 18604 36876
rect 18656 36864 18662 36916
rect 18690 36864 18696 36916
rect 18748 36904 18754 36916
rect 18785 36907 18843 36913
rect 18785 36904 18797 36907
rect 18748 36876 18797 36904
rect 18748 36864 18754 36876
rect 18785 36873 18797 36876
rect 18831 36873 18843 36907
rect 18785 36867 18843 36873
rect 18984 36876 20484 36904
rect 12342 36796 12348 36848
rect 12400 36836 12406 36848
rect 12986 36836 12992 36848
rect 12400 36808 12992 36836
rect 12400 36796 12406 36808
rect 12986 36796 12992 36808
rect 13044 36836 13050 36848
rect 13044 36808 13202 36836
rect 13044 36796 13050 36808
rect 15562 36796 15568 36848
rect 15620 36796 15626 36848
rect 12434 36728 12440 36780
rect 12492 36728 12498 36780
rect 14642 36728 14648 36780
rect 14700 36768 14706 36780
rect 14737 36771 14795 36777
rect 14737 36768 14749 36771
rect 14700 36740 14749 36768
rect 14700 36728 14706 36740
rect 14737 36737 14749 36740
rect 14783 36737 14795 36771
rect 14737 36731 14795 36737
rect 12713 36703 12771 36709
rect 12713 36669 12725 36703
rect 12759 36700 12771 36703
rect 13722 36700 13728 36712
rect 12759 36672 13728 36700
rect 12759 36669 12771 36672
rect 12713 36663 12771 36669
rect 13722 36660 13728 36672
rect 13780 36660 13786 36712
rect 14366 36660 14372 36712
rect 14424 36660 14430 36712
rect 11698 36524 11704 36576
rect 11756 36564 11762 36576
rect 12069 36567 12127 36573
rect 12069 36564 12081 36567
rect 11756 36536 12081 36564
rect 11756 36524 11762 36536
rect 12069 36533 12081 36536
rect 12115 36533 12127 36567
rect 12069 36527 12127 36533
rect 12897 36567 12955 36573
rect 12897 36533 12909 36567
rect 12943 36564 12955 36567
rect 13078 36564 13084 36576
rect 12943 36536 13084 36564
rect 12943 36533 12955 36536
rect 12897 36527 12955 36533
rect 13078 36524 13084 36536
rect 13136 36524 13142 36576
rect 14752 36564 14780 36731
rect 16390 36728 16396 36780
rect 16448 36768 16454 36780
rect 18325 36771 18383 36777
rect 16448 36740 18276 36768
rect 16448 36728 16454 36740
rect 15013 36703 15071 36709
rect 15013 36669 15025 36703
rect 15059 36700 15071 36703
rect 15059 36672 16574 36700
rect 15059 36669 15071 36672
rect 15013 36663 15071 36669
rect 16546 36632 16574 36672
rect 17126 36660 17132 36712
rect 17184 36660 17190 36712
rect 17313 36703 17371 36709
rect 17313 36669 17325 36703
rect 17359 36700 17371 36703
rect 17678 36700 17684 36712
rect 17359 36672 17684 36700
rect 17359 36669 17371 36672
rect 17313 36663 17371 36669
rect 17678 36660 17684 36672
rect 17736 36660 17742 36712
rect 18248 36700 18276 36740
rect 18325 36737 18337 36771
rect 18371 36768 18383 36771
rect 18782 36768 18788 36780
rect 18371 36740 18788 36768
rect 18371 36737 18383 36740
rect 18325 36731 18383 36737
rect 18782 36728 18788 36740
rect 18840 36728 18846 36780
rect 18601 36703 18659 36709
rect 18601 36700 18613 36703
rect 18248 36672 18613 36700
rect 18601 36669 18613 36672
rect 18647 36700 18659 36703
rect 18984 36700 19012 36876
rect 19518 36796 19524 36848
rect 19576 36796 19582 36848
rect 20456 36836 20484 36876
rect 22002 36864 22008 36916
rect 22060 36904 22066 36916
rect 22060 36876 23612 36904
rect 22060 36864 22066 36876
rect 21818 36836 21824 36848
rect 20456 36808 21824 36836
rect 21818 36796 21824 36808
rect 21876 36796 21882 36848
rect 21085 36771 21143 36777
rect 21085 36737 21097 36771
rect 21131 36737 21143 36771
rect 21085 36731 21143 36737
rect 18647 36672 19012 36700
rect 18647 36669 18659 36672
rect 18601 36663 18659 36669
rect 19886 36660 19892 36712
rect 19944 36700 19950 36712
rect 20257 36703 20315 36709
rect 20257 36700 20269 36703
rect 19944 36672 20269 36700
rect 19944 36660 19950 36672
rect 20257 36669 20269 36672
rect 20303 36669 20315 36703
rect 20257 36663 20315 36669
rect 20530 36660 20536 36712
rect 20588 36660 20594 36712
rect 20806 36660 20812 36712
rect 20864 36660 20870 36712
rect 20990 36660 20996 36712
rect 21048 36660 21054 36712
rect 16669 36635 16727 36641
rect 16669 36632 16681 36635
rect 16546 36604 16681 36632
rect 16669 36601 16681 36604
rect 16715 36601 16727 36635
rect 16669 36595 16727 36601
rect 15194 36564 15200 36576
rect 14752 36536 15200 36564
rect 15194 36524 15200 36536
rect 15252 36524 15258 36576
rect 17494 36524 17500 36576
rect 17552 36564 17558 36576
rect 17957 36567 18015 36573
rect 17957 36564 17969 36567
rect 17552 36536 17969 36564
rect 17552 36524 17558 36536
rect 17957 36533 17969 36536
rect 18003 36533 18015 36567
rect 17957 36527 18015 36533
rect 20070 36524 20076 36576
rect 20128 36564 20134 36576
rect 21100 36564 21128 36731
rect 21266 36728 21272 36780
rect 21324 36768 21330 36780
rect 22278 36768 22284 36780
rect 21324 36740 22284 36768
rect 21324 36728 21330 36740
rect 22278 36728 22284 36740
rect 22336 36728 22342 36780
rect 23584 36777 23612 36876
rect 23842 36864 23848 36916
rect 23900 36904 23906 36916
rect 24765 36907 24823 36913
rect 24765 36904 24777 36907
rect 23900 36876 24777 36904
rect 23900 36864 23906 36876
rect 24765 36873 24777 36876
rect 24811 36873 24823 36907
rect 24765 36867 24823 36873
rect 25406 36864 25412 36916
rect 25464 36904 25470 36916
rect 25593 36907 25651 36913
rect 25593 36904 25605 36907
rect 25464 36876 25605 36904
rect 25464 36864 25470 36876
rect 25593 36873 25605 36876
rect 25639 36873 25651 36907
rect 25593 36867 25651 36873
rect 24394 36796 24400 36848
rect 24452 36836 24458 36848
rect 25608 36836 25636 36867
rect 25866 36864 25872 36916
rect 25924 36904 25930 36916
rect 26053 36907 26111 36913
rect 26053 36904 26065 36907
rect 25924 36876 26065 36904
rect 25924 36864 25930 36876
rect 26053 36873 26065 36876
rect 26099 36873 26111 36907
rect 26053 36867 26111 36873
rect 26510 36864 26516 36916
rect 26568 36904 26574 36916
rect 26789 36907 26847 36913
rect 26789 36904 26801 36907
rect 26568 36876 26801 36904
rect 26568 36864 26574 36876
rect 26789 36873 26801 36876
rect 26835 36873 26847 36907
rect 29273 36907 29331 36913
rect 29273 36904 29285 36907
rect 26789 36867 26847 36873
rect 27632 36876 29285 36904
rect 26421 36839 26479 36845
rect 24452 36808 24992 36836
rect 25608 36808 26280 36836
rect 24452 36796 24458 36808
rect 23569 36771 23627 36777
rect 23569 36737 23581 36771
rect 23615 36737 23627 36771
rect 23569 36731 23627 36737
rect 24029 36771 24087 36777
rect 24029 36737 24041 36771
rect 24075 36737 24087 36771
rect 24857 36771 24915 36777
rect 24857 36768 24869 36771
rect 24029 36731 24087 36737
rect 24136 36740 24869 36768
rect 23293 36703 23351 36709
rect 23293 36669 23305 36703
rect 23339 36700 23351 36703
rect 23339 36672 23704 36700
rect 23339 36669 23351 36672
rect 23293 36663 23351 36669
rect 21450 36592 21456 36644
rect 21508 36592 21514 36644
rect 23676 36641 23704 36672
rect 23661 36635 23719 36641
rect 23661 36601 23673 36635
rect 23707 36601 23719 36635
rect 23661 36595 23719 36601
rect 20128 36536 21128 36564
rect 20128 36524 20134 36536
rect 21358 36524 21364 36576
rect 21416 36564 21422 36576
rect 21821 36567 21879 36573
rect 21821 36564 21833 36567
rect 21416 36536 21833 36564
rect 21416 36524 21422 36536
rect 21821 36533 21833 36536
rect 21867 36564 21879 36567
rect 24044 36564 24072 36731
rect 24136 36712 24164 36740
rect 24857 36737 24869 36740
rect 24903 36737 24915 36771
rect 24964 36768 24992 36808
rect 25685 36771 25743 36777
rect 25685 36768 25697 36771
rect 24964 36740 25697 36768
rect 24857 36731 24915 36737
rect 25685 36737 25697 36740
rect 25731 36737 25743 36771
rect 25685 36731 25743 36737
rect 25958 36728 25964 36780
rect 26016 36768 26022 36780
rect 26252 36777 26280 36808
rect 26421 36805 26433 36839
rect 26467 36836 26479 36839
rect 27632 36836 27660 36876
rect 29273 36873 29285 36876
rect 29319 36873 29331 36907
rect 29273 36867 29331 36873
rect 32950 36864 32956 36916
rect 33008 36904 33014 36916
rect 34790 36904 34796 36916
rect 33008 36876 34796 36904
rect 33008 36864 33014 36876
rect 34790 36864 34796 36876
rect 34848 36904 34854 36916
rect 34977 36907 35035 36913
rect 34977 36904 34989 36907
rect 34848 36876 34989 36904
rect 34848 36864 34854 36876
rect 34977 36873 34989 36876
rect 35023 36873 35035 36907
rect 34977 36867 35035 36873
rect 26467 36808 27660 36836
rect 26467 36805 26479 36808
rect 26421 36799 26479 36805
rect 27706 36796 27712 36848
rect 27764 36796 27770 36848
rect 28994 36836 29000 36848
rect 28934 36808 29000 36836
rect 28994 36796 29000 36808
rect 29052 36836 29058 36848
rect 30558 36836 30564 36848
rect 29052 36808 30564 36836
rect 29052 36796 29058 36808
rect 30558 36796 30564 36808
rect 30616 36796 30622 36848
rect 32125 36839 32183 36845
rect 32125 36836 32137 36839
rect 31726 36808 32137 36836
rect 26145 36771 26203 36777
rect 26145 36768 26157 36771
rect 26016 36740 26157 36768
rect 26016 36728 26022 36740
rect 26145 36737 26157 36740
rect 26191 36737 26203 36771
rect 26145 36731 26203 36737
rect 26238 36771 26296 36777
rect 26238 36737 26250 36771
rect 26284 36737 26296 36771
rect 26238 36731 26296 36737
rect 26510 36728 26516 36780
rect 26568 36728 26574 36780
rect 26602 36728 26608 36780
rect 26660 36777 26666 36780
rect 26660 36768 26668 36777
rect 26660 36740 26705 36768
rect 26660 36731 26668 36740
rect 26660 36728 26666 36731
rect 27062 36728 27068 36780
rect 27120 36728 27126 36780
rect 27249 36771 27307 36777
rect 27249 36737 27261 36771
rect 27295 36768 27307 36771
rect 27338 36768 27344 36780
rect 27295 36740 27344 36768
rect 27295 36737 27307 36740
rect 27249 36731 27307 36737
rect 27338 36728 27344 36740
rect 27396 36728 27402 36780
rect 29457 36771 29515 36777
rect 29457 36737 29469 36771
rect 29503 36768 29515 36771
rect 29503 36740 29684 36768
rect 29503 36737 29515 36740
rect 29457 36731 29515 36737
rect 24118 36660 24124 36712
rect 24176 36660 24182 36712
rect 24305 36703 24363 36709
rect 24305 36669 24317 36703
rect 24351 36669 24363 36703
rect 24305 36663 24363 36669
rect 24581 36703 24639 36709
rect 24581 36669 24593 36703
rect 24627 36700 24639 36703
rect 24627 36672 24900 36700
rect 24627 36669 24639 36672
rect 24581 36663 24639 36669
rect 24320 36632 24348 36663
rect 24872 36644 24900 36672
rect 25498 36660 25504 36712
rect 25556 36660 25562 36712
rect 27433 36703 27491 36709
rect 27433 36700 27445 36703
rect 26160 36672 27445 36700
rect 26160 36644 26188 36672
rect 27433 36669 27445 36672
rect 27479 36669 27491 36703
rect 29472 36700 29500 36731
rect 27433 36663 27491 36669
rect 27540 36672 29500 36700
rect 24670 36632 24676 36644
rect 24320 36604 24676 36632
rect 24670 36592 24676 36604
rect 24728 36592 24734 36644
rect 24854 36592 24860 36644
rect 24912 36592 24918 36644
rect 26142 36592 26148 36644
rect 26200 36592 26206 36644
rect 27246 36592 27252 36644
rect 27304 36592 27310 36644
rect 27338 36592 27344 36644
rect 27396 36632 27402 36644
rect 27540 36632 27568 36672
rect 29546 36660 29552 36712
rect 29604 36660 29610 36712
rect 29656 36700 29684 36740
rect 29730 36728 29736 36780
rect 29788 36728 29794 36780
rect 30374 36728 30380 36780
rect 30432 36768 30438 36780
rect 31018 36768 31024 36780
rect 30432 36740 31024 36768
rect 30432 36728 30438 36740
rect 31018 36728 31024 36740
rect 31076 36728 31082 36780
rect 31110 36728 31116 36780
rect 31168 36768 31174 36780
rect 31726 36768 31754 36808
rect 32125 36805 32137 36808
rect 32171 36805 32183 36839
rect 32125 36799 32183 36805
rect 32306 36796 32312 36848
rect 32364 36845 32370 36848
rect 32364 36839 32399 36845
rect 32387 36836 32399 36839
rect 32585 36839 32643 36845
rect 32585 36836 32597 36839
rect 32387 36808 32597 36836
rect 32387 36805 32399 36808
rect 32364 36799 32399 36805
rect 32585 36805 32597 36808
rect 32631 36836 32643 36839
rect 33410 36836 33416 36848
rect 32631 36808 33416 36836
rect 32631 36805 32643 36808
rect 32585 36799 32643 36805
rect 32364 36796 32370 36799
rect 33410 36796 33416 36808
rect 33468 36796 33474 36848
rect 33962 36796 33968 36848
rect 34020 36796 34026 36848
rect 31168 36740 31754 36768
rect 31941 36771 31999 36777
rect 31168 36728 31174 36740
rect 31941 36737 31953 36771
rect 31987 36737 31999 36771
rect 31941 36731 31999 36737
rect 31662 36700 31668 36712
rect 29656 36672 31668 36700
rect 31662 36660 31668 36672
rect 31720 36660 31726 36712
rect 31956 36700 31984 36731
rect 32030 36728 32036 36780
rect 32088 36768 32094 36780
rect 32769 36771 32827 36777
rect 32769 36768 32781 36771
rect 32088 36740 32781 36768
rect 32088 36728 32094 36740
rect 32122 36700 32128 36712
rect 31956 36672 32128 36700
rect 32122 36660 32128 36672
rect 32180 36660 32186 36712
rect 27396 36604 27568 36632
rect 27396 36592 27402 36604
rect 32416 36576 32444 36740
rect 32769 36737 32781 36740
rect 32815 36737 32827 36771
rect 32769 36731 32827 36737
rect 32861 36771 32919 36777
rect 32861 36737 32873 36771
rect 32907 36768 32919 36771
rect 33134 36768 33140 36780
rect 32907 36740 33140 36768
rect 32907 36737 32919 36740
rect 32861 36731 32919 36737
rect 33134 36728 33140 36740
rect 33192 36728 33198 36780
rect 33226 36728 33232 36780
rect 33284 36728 33290 36780
rect 33502 36660 33508 36712
rect 33560 36660 33566 36712
rect 21867 36536 24072 36564
rect 21867 36533 21879 36536
rect 21821 36527 21879 36533
rect 25222 36524 25228 36576
rect 25280 36524 25286 36576
rect 27430 36524 27436 36576
rect 27488 36564 27494 36576
rect 29181 36567 29239 36573
rect 29181 36564 29193 36567
rect 27488 36536 29193 36564
rect 27488 36524 27494 36536
rect 29181 36533 29193 36536
rect 29227 36564 29239 36567
rect 30098 36564 30104 36576
rect 29227 36536 30104 36564
rect 29227 36533 29239 36536
rect 29181 36527 29239 36533
rect 30098 36524 30104 36536
rect 30156 36524 30162 36576
rect 31294 36524 31300 36576
rect 31352 36564 31358 36576
rect 31481 36567 31539 36573
rect 31481 36564 31493 36567
rect 31352 36536 31493 36564
rect 31352 36524 31358 36536
rect 31481 36533 31493 36536
rect 31527 36533 31539 36567
rect 31481 36527 31539 36533
rect 32309 36567 32367 36573
rect 32309 36533 32321 36567
rect 32355 36564 32367 36567
rect 32398 36564 32404 36576
rect 32355 36536 32404 36564
rect 32355 36533 32367 36536
rect 32309 36527 32367 36533
rect 32398 36524 32404 36536
rect 32456 36524 32462 36576
rect 32493 36567 32551 36573
rect 32493 36533 32505 36567
rect 32539 36564 32551 36567
rect 32858 36564 32864 36576
rect 32539 36536 32864 36564
rect 32539 36533 32551 36536
rect 32493 36527 32551 36533
rect 32858 36524 32864 36536
rect 32916 36524 32922 36576
rect 33137 36567 33195 36573
rect 33137 36533 33149 36567
rect 33183 36564 33195 36567
rect 33318 36564 33324 36576
rect 33183 36536 33324 36564
rect 33183 36533 33195 36536
rect 33137 36527 33195 36533
rect 33318 36524 33324 36536
rect 33376 36524 33382 36576
rect 1104 36474 37076 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 37076 36474
rect 1104 36400 37076 36422
rect 12434 36320 12440 36372
rect 12492 36360 12498 36372
rect 12986 36360 12992 36372
rect 12492 36332 12992 36360
rect 12492 36320 12498 36332
rect 12986 36320 12992 36332
rect 13044 36360 13050 36372
rect 13173 36363 13231 36369
rect 13173 36360 13185 36363
rect 13044 36332 13185 36360
rect 13044 36320 13050 36332
rect 13173 36329 13185 36332
rect 13219 36329 13231 36363
rect 13173 36323 13231 36329
rect 14185 36363 14243 36369
rect 14185 36329 14197 36363
rect 14231 36360 14243 36363
rect 14366 36360 14372 36372
rect 14231 36332 14372 36360
rect 14231 36329 14243 36332
rect 14185 36323 14243 36329
rect 14366 36320 14372 36332
rect 14424 36320 14430 36372
rect 18506 36320 18512 36372
rect 18564 36360 18570 36372
rect 18782 36360 18788 36372
rect 18564 36332 18788 36360
rect 18564 36320 18570 36332
rect 18782 36320 18788 36332
rect 18840 36360 18846 36372
rect 18969 36363 19027 36369
rect 18969 36360 18981 36363
rect 18840 36332 18981 36360
rect 18840 36320 18846 36332
rect 18969 36329 18981 36332
rect 19015 36329 19027 36363
rect 18969 36323 19027 36329
rect 20990 36320 20996 36372
rect 21048 36360 21054 36372
rect 21729 36363 21787 36369
rect 21729 36360 21741 36363
rect 21048 36332 21741 36360
rect 21048 36320 21054 36332
rect 21729 36329 21741 36332
rect 21775 36329 21787 36363
rect 21729 36323 21787 36329
rect 21818 36320 21824 36372
rect 21876 36360 21882 36372
rect 22281 36363 22339 36369
rect 22281 36360 22293 36363
rect 21876 36332 22293 36360
rect 21876 36320 21882 36332
rect 22281 36329 22293 36332
rect 22327 36360 22339 36363
rect 25498 36360 25504 36372
rect 22327 36332 25504 36360
rect 22327 36329 22339 36332
rect 22281 36323 22339 36329
rect 25498 36320 25504 36332
rect 25556 36320 25562 36372
rect 25958 36320 25964 36372
rect 26016 36360 26022 36372
rect 26145 36363 26203 36369
rect 26145 36360 26157 36363
rect 26016 36332 26157 36360
rect 26016 36320 26022 36332
rect 26145 36329 26157 36332
rect 26191 36329 26203 36363
rect 26145 36323 26203 36329
rect 26510 36320 26516 36372
rect 26568 36360 26574 36372
rect 28537 36363 28595 36369
rect 26568 36332 28488 36360
rect 26568 36320 26574 36332
rect 24946 36252 24952 36304
rect 25004 36292 25010 36304
rect 25041 36295 25099 36301
rect 25041 36292 25053 36295
rect 25004 36264 25053 36292
rect 25004 36252 25010 36264
rect 25041 36261 25053 36264
rect 25087 36261 25099 36295
rect 25041 36255 25099 36261
rect 11698 36184 11704 36236
rect 11756 36184 11762 36236
rect 13722 36184 13728 36236
rect 13780 36224 13786 36236
rect 14829 36227 14887 36233
rect 14829 36224 14841 36227
rect 13780 36196 14841 36224
rect 13780 36184 13786 36196
rect 14829 36193 14841 36196
rect 14875 36224 14887 36227
rect 16390 36224 16396 36236
rect 14875 36196 16396 36224
rect 14875 36193 14887 36196
rect 14829 36187 14887 36193
rect 16390 36184 16396 36196
rect 16448 36184 16454 36236
rect 16482 36184 16488 36236
rect 16540 36224 16546 36236
rect 17221 36227 17279 36233
rect 17221 36224 17233 36227
rect 16540 36196 17233 36224
rect 16540 36184 16546 36196
rect 17221 36193 17233 36196
rect 17267 36193 17279 36227
rect 17221 36187 17279 36193
rect 17494 36184 17500 36236
rect 17552 36184 17558 36236
rect 20257 36227 20315 36233
rect 20257 36193 20269 36227
rect 20303 36224 20315 36227
rect 20898 36224 20904 36236
rect 20303 36196 20904 36224
rect 20303 36193 20315 36196
rect 20257 36187 20315 36193
rect 20898 36184 20904 36196
rect 20956 36184 20962 36236
rect 25406 36184 25412 36236
rect 25464 36224 25470 36236
rect 26142 36224 26148 36236
rect 25464 36196 26148 36224
rect 25464 36184 25470 36196
rect 26142 36184 26148 36196
rect 26200 36224 26206 36236
rect 26789 36227 26847 36233
rect 26789 36224 26801 36227
rect 26200 36196 26801 36224
rect 26200 36184 26206 36196
rect 26789 36193 26801 36196
rect 26835 36193 26847 36227
rect 26789 36187 26847 36193
rect 27065 36227 27123 36233
rect 27065 36193 27077 36227
rect 27111 36224 27123 36227
rect 27614 36224 27620 36236
rect 27111 36196 27620 36224
rect 27111 36193 27123 36196
rect 27065 36187 27123 36193
rect 27614 36184 27620 36196
rect 27672 36184 27678 36236
rect 11425 36159 11483 36165
rect 11425 36125 11437 36159
rect 11471 36125 11483 36159
rect 11425 36119 11483 36125
rect 11440 36020 11468 36119
rect 13078 36116 13084 36168
rect 13136 36156 13142 36168
rect 14553 36159 14611 36165
rect 14553 36156 14565 36159
rect 13136 36128 14565 36156
rect 13136 36116 13142 36128
rect 14553 36125 14565 36128
rect 14599 36125 14611 36159
rect 14553 36119 14611 36125
rect 14645 36159 14703 36165
rect 14645 36125 14657 36159
rect 14691 36156 14703 36159
rect 15470 36156 15476 36168
rect 14691 36128 15476 36156
rect 14691 36125 14703 36128
rect 14645 36119 14703 36125
rect 15470 36116 15476 36128
rect 15528 36116 15534 36168
rect 19978 36116 19984 36168
rect 20036 36116 20042 36168
rect 25317 36159 25375 36165
rect 25317 36125 25329 36159
rect 25363 36156 25375 36159
rect 25774 36156 25780 36168
rect 25363 36128 25780 36156
rect 25363 36125 25375 36128
rect 25317 36119 25375 36125
rect 25774 36116 25780 36128
rect 25832 36116 25838 36168
rect 25869 36159 25927 36165
rect 25869 36125 25881 36159
rect 25915 36125 25927 36159
rect 25869 36119 25927 36125
rect 12342 36048 12348 36100
rect 12400 36048 12406 36100
rect 19518 36088 19524 36100
rect 18722 36060 19524 36088
rect 11514 36020 11520 36032
rect 11440 35992 11520 36020
rect 11514 35980 11520 35992
rect 11572 35980 11578 36032
rect 18138 35980 18144 36032
rect 18196 36020 18202 36032
rect 18800 36020 18828 36060
rect 19518 36048 19524 36060
rect 19576 36048 19582 36100
rect 19996 36088 20024 36116
rect 20530 36088 20536 36100
rect 19996 36060 20536 36088
rect 20530 36048 20536 36060
rect 20588 36048 20594 36100
rect 21266 36048 21272 36100
rect 21324 36048 21330 36100
rect 23569 36091 23627 36097
rect 23569 36057 23581 36091
rect 23615 36088 23627 36091
rect 24762 36088 24768 36100
rect 23615 36060 24768 36088
rect 23615 36057 23627 36060
rect 23569 36051 23627 36057
rect 24762 36048 24768 36060
rect 24820 36048 24826 36100
rect 25593 36091 25651 36097
rect 25593 36088 25605 36091
rect 25424 36060 25605 36088
rect 18196 35992 18828 36020
rect 18196 35980 18202 35992
rect 24670 35980 24676 36032
rect 24728 36020 24734 36032
rect 25424 36020 25452 36060
rect 25593 36057 25605 36060
rect 25639 36088 25651 36091
rect 25884 36088 25912 36119
rect 25958 36116 25964 36168
rect 26016 36116 26022 36168
rect 28460 36156 28488 36332
rect 28537 36329 28549 36363
rect 28583 36360 28595 36363
rect 29178 36360 29184 36372
rect 28583 36332 29184 36360
rect 28583 36329 28595 36332
rect 28537 36323 28595 36329
rect 29178 36320 29184 36332
rect 29236 36320 29242 36372
rect 29546 36320 29552 36372
rect 29604 36360 29610 36372
rect 29914 36360 29920 36372
rect 29604 36332 29920 36360
rect 29604 36320 29610 36332
rect 29914 36320 29920 36332
rect 29972 36360 29978 36372
rect 30926 36360 30932 36372
rect 29972 36332 30932 36360
rect 29972 36320 29978 36332
rect 30926 36320 30932 36332
rect 30984 36320 30990 36372
rect 31018 36320 31024 36372
rect 31076 36360 31082 36372
rect 32030 36360 32036 36372
rect 31076 36332 32036 36360
rect 31076 36320 31082 36332
rect 28718 36252 28724 36304
rect 28776 36292 28782 36304
rect 28776 36264 31524 36292
rect 28776 36252 28782 36264
rect 28920 36233 28948 36264
rect 28905 36227 28963 36233
rect 28905 36193 28917 36227
rect 28951 36193 28963 36227
rect 29546 36224 29552 36236
rect 28905 36187 28963 36193
rect 29196 36196 29552 36224
rect 28718 36156 28724 36168
rect 28460 36128 28724 36156
rect 28718 36116 28724 36128
rect 28776 36156 28782 36168
rect 29196 36156 29224 36196
rect 29546 36184 29552 36196
rect 29604 36184 29610 36236
rect 30098 36184 30104 36236
rect 30156 36184 30162 36236
rect 30285 36227 30343 36233
rect 30285 36193 30297 36227
rect 30331 36224 30343 36227
rect 30466 36224 30472 36236
rect 30331 36196 30472 36224
rect 30331 36193 30343 36196
rect 30285 36187 30343 36193
rect 30466 36184 30472 36196
rect 30524 36184 30530 36236
rect 31021 36227 31079 36233
rect 31021 36224 31033 36227
rect 30576 36196 31033 36224
rect 28776 36128 29224 36156
rect 29273 36159 29331 36165
rect 28776 36116 28782 36128
rect 29273 36125 29285 36159
rect 29319 36156 29331 36159
rect 29362 36156 29368 36168
rect 29319 36128 29368 36156
rect 29319 36125 29331 36128
rect 29273 36119 29331 36125
rect 29362 36116 29368 36128
rect 29420 36116 29426 36168
rect 25639 36060 25912 36088
rect 28290 36060 28396 36088
rect 25639 36057 25651 36060
rect 25593 36051 25651 36057
rect 24728 35992 25452 36020
rect 24728 35980 24734 35992
rect 25498 35980 25504 36032
rect 25556 35980 25562 36032
rect 28368 36020 28396 36060
rect 28810 36048 28816 36100
rect 28868 36088 28874 36100
rect 30576 36088 30604 36196
rect 31021 36193 31033 36196
rect 31067 36224 31079 36227
rect 31110 36224 31116 36236
rect 31067 36196 31116 36224
rect 31067 36193 31079 36196
rect 31021 36187 31079 36193
rect 31110 36184 31116 36196
rect 31168 36184 31174 36236
rect 30745 36159 30803 36165
rect 30745 36125 30757 36159
rect 30791 36125 30803 36159
rect 30745 36119 30803 36125
rect 28868 36060 30604 36088
rect 28868 36048 28874 36060
rect 28902 36020 28908 36032
rect 28368 35992 28908 36020
rect 28902 35980 28908 35992
rect 28960 35980 28966 36032
rect 28994 35980 29000 36032
rect 29052 36020 29058 36032
rect 29641 36023 29699 36029
rect 29641 36020 29653 36023
rect 29052 35992 29653 36020
rect 29052 35980 29058 35992
rect 29641 35989 29653 35992
rect 29687 35989 29699 36023
rect 30760 36020 30788 36119
rect 30926 36116 30932 36168
rect 30984 36116 30990 36168
rect 31386 36048 31392 36100
rect 31444 36048 31450 36100
rect 31496 36088 31524 36264
rect 31588 36165 31616 36332
rect 32030 36320 32036 36332
rect 32088 36320 32094 36372
rect 33502 36320 33508 36372
rect 33560 36320 33566 36372
rect 31846 36252 31852 36304
rect 31904 36292 31910 36304
rect 34701 36295 34759 36301
rect 31904 36264 32260 36292
rect 31904 36252 31910 36264
rect 32122 36224 32128 36236
rect 31726 36196 32128 36224
rect 31573 36159 31631 36165
rect 31573 36125 31585 36159
rect 31619 36125 31631 36159
rect 31573 36119 31631 36125
rect 31726 36088 31754 36196
rect 32122 36184 32128 36196
rect 32180 36184 32186 36236
rect 32232 36165 32260 36264
rect 34701 36261 34713 36295
rect 34747 36261 34759 36295
rect 34701 36255 34759 36261
rect 32306 36184 32312 36236
rect 32364 36224 32370 36236
rect 32585 36227 32643 36233
rect 32585 36224 32597 36227
rect 32364 36196 32597 36224
rect 32364 36184 32370 36196
rect 32585 36193 32597 36196
rect 32631 36193 32643 36227
rect 34716 36224 34744 36255
rect 34790 36252 34796 36304
rect 34848 36292 34854 36304
rect 34848 36264 34928 36292
rect 34848 36252 34854 36264
rect 32585 36187 32643 36193
rect 33520 36196 34744 36224
rect 32033 36159 32091 36165
rect 32033 36125 32045 36159
rect 32079 36125 32091 36159
rect 32033 36119 32091 36125
rect 32217 36159 32275 36165
rect 32217 36125 32229 36159
rect 32263 36125 32275 36159
rect 32217 36119 32275 36125
rect 31496 36060 31754 36088
rect 31846 36048 31852 36100
rect 31904 36088 31910 36100
rect 31941 36091 31999 36097
rect 31941 36088 31953 36091
rect 31904 36060 31953 36088
rect 31904 36048 31910 36060
rect 31941 36057 31953 36060
rect 31987 36057 31999 36091
rect 31941 36051 31999 36057
rect 32048 36088 32076 36119
rect 33134 36116 33140 36168
rect 33192 36156 33198 36168
rect 33229 36159 33287 36165
rect 33229 36156 33241 36159
rect 33192 36128 33241 36156
rect 33192 36116 33198 36128
rect 33229 36125 33241 36128
rect 33275 36125 33287 36159
rect 33229 36119 33287 36125
rect 33318 36116 33324 36168
rect 33376 36116 33382 36168
rect 33520 36165 33548 36196
rect 33505 36159 33563 36165
rect 33505 36125 33517 36159
rect 33551 36125 33563 36159
rect 33505 36119 33563 36125
rect 33594 36116 33600 36168
rect 33652 36116 33658 36168
rect 33873 36159 33931 36165
rect 33873 36125 33885 36159
rect 33919 36156 33931 36159
rect 34790 36156 34796 36168
rect 33919 36128 34796 36156
rect 33919 36125 33931 36128
rect 33873 36119 33931 36125
rect 34790 36116 34796 36128
rect 34848 36116 34854 36168
rect 34900 36165 34928 36264
rect 34885 36159 34943 36165
rect 34885 36125 34897 36159
rect 34931 36125 34943 36159
rect 34885 36119 34943 36125
rect 34977 36159 35035 36165
rect 34977 36125 34989 36159
rect 35023 36125 35035 36159
rect 34977 36119 35035 36125
rect 32398 36088 32404 36100
rect 32048 36060 32404 36088
rect 32048 36020 32076 36060
rect 32398 36048 32404 36060
rect 32456 36048 32462 36100
rect 34701 36091 34759 36097
rect 34701 36088 34713 36091
rect 33520 36060 34713 36088
rect 30760 35992 32076 36020
rect 29641 35983 29699 35989
rect 32214 35980 32220 36032
rect 32272 35980 32278 36032
rect 32766 35980 32772 36032
rect 32824 35980 32830 36032
rect 32858 35980 32864 36032
rect 32916 36020 32922 36032
rect 33520 36020 33548 36060
rect 34701 36057 34713 36060
rect 34747 36057 34759 36091
rect 34701 36051 34759 36057
rect 32916 35992 33548 36020
rect 32916 35980 32922 35992
rect 34606 35980 34612 36032
rect 34664 36020 34670 36032
rect 34992 36020 35020 36119
rect 34664 35992 35020 36020
rect 34664 35980 34670 35992
rect 1104 35930 37076 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 37076 35930
rect 1104 35856 37076 35878
rect 12986 35776 12992 35828
rect 13044 35776 13050 35828
rect 18506 35776 18512 35828
rect 18564 35816 18570 35828
rect 18693 35819 18751 35825
rect 18693 35816 18705 35819
rect 18564 35788 18705 35816
rect 18564 35776 18570 35788
rect 18693 35785 18705 35788
rect 18739 35785 18751 35819
rect 18693 35779 18751 35785
rect 20898 35776 20904 35828
rect 20956 35776 20962 35828
rect 20990 35776 20996 35828
rect 21048 35816 21054 35828
rect 21269 35819 21327 35825
rect 21269 35816 21281 35819
rect 21048 35788 21281 35816
rect 21048 35776 21054 35788
rect 21269 35785 21281 35788
rect 21315 35785 21327 35819
rect 21269 35779 21327 35785
rect 21358 35776 21364 35828
rect 21416 35776 21422 35828
rect 23661 35819 23719 35825
rect 23661 35785 23673 35819
rect 23707 35816 23719 35819
rect 24118 35816 24124 35828
rect 23707 35788 24124 35816
rect 23707 35785 23719 35788
rect 23661 35779 23719 35785
rect 24118 35776 24124 35788
rect 24176 35776 24182 35828
rect 26329 35819 26387 35825
rect 26329 35785 26341 35819
rect 26375 35816 26387 35819
rect 27233 35819 27291 35825
rect 27233 35816 27245 35819
rect 26375 35788 27245 35816
rect 26375 35785 26387 35788
rect 26329 35779 26387 35785
rect 27233 35785 27245 35788
rect 27279 35816 27291 35819
rect 27279 35788 28488 35816
rect 27279 35785 27291 35788
rect 27233 35779 27291 35785
rect 16117 35751 16175 35757
rect 16117 35717 16129 35751
rect 16163 35748 16175 35751
rect 16942 35748 16948 35760
rect 16163 35720 16948 35748
rect 16163 35717 16175 35720
rect 16117 35711 16175 35717
rect 16942 35708 16948 35720
rect 17000 35708 17006 35760
rect 20806 35708 20812 35760
rect 20864 35748 20870 35760
rect 21821 35751 21879 35757
rect 21821 35748 21833 35751
rect 20864 35720 21833 35748
rect 20864 35708 20870 35720
rect 21821 35717 21833 35720
rect 21867 35717 21879 35751
rect 21821 35711 21879 35717
rect 22278 35708 22284 35760
rect 22336 35748 22342 35760
rect 25133 35751 25191 35757
rect 22336 35734 23966 35748
rect 22336 35720 23980 35734
rect 22336 35708 22342 35720
rect 11882 35640 11888 35692
rect 11940 35680 11946 35692
rect 13081 35683 13139 35689
rect 13081 35680 13093 35683
rect 11940 35652 13093 35680
rect 11940 35640 11946 35652
rect 13081 35649 13093 35652
rect 13127 35649 13139 35683
rect 13081 35643 13139 35649
rect 18601 35683 18659 35689
rect 18601 35649 18613 35683
rect 18647 35680 18659 35683
rect 19058 35680 19064 35692
rect 18647 35652 19064 35680
rect 18647 35649 18659 35652
rect 18601 35643 18659 35649
rect 19058 35640 19064 35652
rect 19116 35640 19122 35692
rect 12897 35615 12955 35621
rect 12897 35581 12909 35615
rect 12943 35612 12955 35615
rect 13722 35612 13728 35624
rect 12943 35584 13728 35612
rect 12943 35581 12955 35584
rect 12897 35575 12955 35581
rect 13722 35572 13728 35584
rect 13780 35572 13786 35624
rect 16206 35572 16212 35624
rect 16264 35572 16270 35624
rect 16390 35572 16396 35624
rect 16448 35572 16454 35624
rect 18874 35572 18880 35624
rect 18932 35612 18938 35624
rect 20254 35612 20260 35624
rect 18932 35584 20260 35612
rect 18932 35572 18938 35584
rect 20254 35572 20260 35584
rect 20312 35612 20318 35624
rect 20824 35612 20852 35708
rect 23566 35640 23572 35692
rect 23624 35640 23630 35692
rect 20312 35584 20852 35612
rect 20312 35572 20318 35584
rect 21450 35572 21456 35624
rect 21508 35572 21514 35624
rect 23952 35612 23980 35720
rect 25133 35717 25145 35751
rect 25179 35748 25191 35751
rect 25222 35748 25228 35760
rect 25179 35720 25228 35748
rect 25179 35717 25191 35720
rect 25133 35711 25191 35717
rect 25222 35708 25228 35720
rect 25280 35708 25286 35760
rect 27433 35751 27491 35757
rect 27433 35717 27445 35751
rect 27479 35717 27491 35751
rect 27433 35711 27491 35717
rect 27525 35751 27583 35757
rect 27525 35717 27537 35751
rect 27571 35748 27583 35751
rect 27614 35748 27620 35760
rect 27571 35720 27620 35748
rect 27571 35717 27583 35720
rect 27525 35711 27583 35717
rect 27448 35680 27476 35711
rect 27614 35708 27620 35720
rect 27672 35708 27678 35760
rect 27706 35680 27712 35692
rect 27448 35652 27712 35680
rect 27706 35640 27712 35652
rect 27764 35640 27770 35692
rect 27982 35640 27988 35692
rect 28040 35640 28046 35692
rect 28169 35683 28227 35689
rect 28169 35649 28181 35683
rect 28215 35649 28227 35683
rect 28169 35643 28227 35649
rect 25130 35612 25136 35624
rect 23952 35584 25136 35612
rect 25130 35572 25136 35584
rect 25188 35572 25194 35624
rect 25406 35572 25412 35624
rect 25464 35572 25470 35624
rect 26234 35572 26240 35624
rect 26292 35612 26298 35624
rect 26789 35615 26847 35621
rect 26789 35612 26801 35615
rect 26292 35584 26801 35612
rect 26292 35572 26298 35584
rect 26789 35581 26801 35584
rect 26835 35581 26847 35615
rect 26789 35575 26847 35581
rect 27246 35572 27252 35624
rect 27304 35612 27310 35624
rect 28184 35612 28212 35643
rect 27304 35584 28212 35612
rect 28261 35615 28319 35621
rect 27304 35572 27310 35584
rect 28261 35581 28273 35615
rect 28307 35581 28319 35615
rect 28460 35612 28488 35788
rect 31754 35776 31760 35828
rect 31812 35816 31818 35828
rect 32125 35819 32183 35825
rect 32125 35816 32137 35819
rect 31812 35788 32137 35816
rect 31812 35776 31818 35788
rect 32125 35785 32137 35788
rect 32171 35785 32183 35819
rect 32125 35779 32183 35785
rect 33134 35776 33140 35828
rect 33192 35816 33198 35828
rect 34238 35816 34244 35828
rect 33192 35788 34244 35816
rect 33192 35776 33198 35788
rect 34238 35776 34244 35788
rect 34296 35776 34302 35828
rect 29641 35751 29699 35757
rect 29641 35717 29653 35751
rect 29687 35748 29699 35751
rect 30101 35751 30159 35757
rect 30101 35748 30113 35751
rect 29687 35720 30113 35748
rect 29687 35717 29699 35720
rect 29641 35711 29699 35717
rect 30101 35717 30113 35720
rect 30147 35717 30159 35751
rect 30101 35711 30159 35717
rect 30558 35708 30564 35760
rect 30616 35708 30622 35760
rect 31386 35708 31392 35760
rect 31444 35748 31450 35760
rect 31444 35720 32352 35748
rect 31444 35708 31450 35720
rect 28534 35640 28540 35692
rect 28592 35680 28598 35692
rect 28905 35683 28963 35689
rect 28905 35680 28917 35683
rect 28592 35652 28917 35680
rect 28592 35640 28598 35652
rect 28905 35649 28917 35652
rect 28951 35649 28963 35683
rect 28905 35643 28963 35649
rect 29549 35683 29607 35689
rect 29549 35649 29561 35683
rect 29595 35649 29607 35683
rect 29549 35643 29607 35649
rect 28629 35615 28687 35621
rect 28629 35612 28641 35615
rect 28460 35584 28641 35612
rect 28261 35575 28319 35581
rect 28629 35581 28641 35584
rect 28675 35581 28687 35615
rect 28629 35575 28687 35581
rect 27062 35504 27068 35556
rect 27120 35544 27126 35556
rect 28276 35544 28304 35575
rect 27120 35516 28304 35544
rect 27120 35504 27126 35516
rect 13354 35436 13360 35488
rect 13412 35476 13418 35488
rect 13449 35479 13507 35485
rect 13449 35476 13461 35479
rect 13412 35448 13461 35476
rect 13412 35436 13418 35448
rect 13449 35445 13461 35448
rect 13495 35445 13507 35479
rect 13449 35439 13507 35445
rect 15470 35436 15476 35488
rect 15528 35476 15534 35488
rect 15749 35479 15807 35485
rect 15749 35476 15761 35479
rect 15528 35448 15761 35476
rect 15528 35436 15534 35448
rect 15749 35445 15761 35448
rect 15795 35445 15807 35479
rect 15749 35439 15807 35445
rect 17586 35436 17592 35488
rect 17644 35476 17650 35488
rect 18233 35479 18291 35485
rect 18233 35476 18245 35479
rect 17644 35448 18245 35476
rect 17644 35436 17650 35448
rect 18233 35445 18245 35448
rect 18279 35445 18291 35479
rect 18233 35439 18291 35445
rect 27249 35479 27307 35485
rect 27249 35445 27261 35479
rect 27295 35476 27307 35479
rect 27430 35476 27436 35488
rect 27295 35448 27436 35476
rect 27295 35445 27307 35448
rect 27249 35439 27307 35445
rect 27430 35436 27436 35448
rect 27488 35436 27494 35488
rect 27706 35436 27712 35488
rect 27764 35476 27770 35488
rect 29362 35476 29368 35488
rect 27764 35448 29368 35476
rect 27764 35436 27770 35448
rect 29362 35436 29368 35448
rect 29420 35436 29426 35488
rect 29564 35476 29592 35643
rect 29730 35640 29736 35692
rect 29788 35640 29794 35692
rect 29822 35640 29828 35692
rect 29880 35640 29886 35692
rect 31570 35640 31576 35692
rect 31628 35680 31634 35692
rect 31665 35683 31723 35689
rect 31665 35680 31677 35683
rect 31628 35652 31677 35680
rect 31628 35640 31634 35652
rect 31665 35649 31677 35652
rect 31711 35649 31723 35683
rect 31665 35643 31723 35649
rect 31754 35640 31760 35692
rect 31812 35680 31818 35692
rect 31849 35683 31907 35689
rect 31849 35680 31861 35683
rect 31812 35652 31861 35680
rect 31812 35640 31818 35652
rect 31849 35649 31861 35652
rect 31895 35649 31907 35683
rect 31849 35643 31907 35649
rect 31941 35683 31999 35689
rect 31941 35649 31953 35683
rect 31987 35680 31999 35683
rect 32214 35680 32220 35692
rect 31987 35652 32220 35680
rect 31987 35649 31999 35652
rect 31941 35643 31999 35649
rect 31665 35547 31723 35553
rect 31665 35544 31677 35547
rect 31128 35516 31677 35544
rect 31128 35476 31156 35516
rect 31665 35513 31677 35516
rect 31711 35513 31723 35547
rect 31665 35507 31723 35513
rect 31846 35504 31852 35556
rect 31904 35544 31910 35556
rect 31956 35544 31984 35643
rect 32214 35640 32220 35652
rect 32272 35640 32278 35692
rect 32324 35624 32352 35720
rect 32306 35572 32312 35624
rect 32364 35612 32370 35624
rect 32585 35615 32643 35621
rect 32585 35612 32597 35615
rect 32364 35584 32597 35612
rect 32364 35572 32370 35584
rect 32585 35581 32597 35584
rect 32631 35581 32643 35615
rect 33152 35612 33180 35776
rect 33226 35708 33232 35760
rect 33284 35748 33290 35760
rect 33962 35748 33968 35760
rect 33284 35720 33968 35748
rect 33284 35708 33290 35720
rect 33318 35640 33324 35692
rect 33376 35640 33382 35692
rect 33413 35683 33471 35689
rect 33413 35649 33425 35683
rect 33459 35649 33471 35683
rect 33413 35643 33471 35649
rect 33229 35615 33287 35621
rect 33229 35612 33241 35615
rect 33152 35584 33241 35612
rect 32585 35575 32643 35581
rect 33229 35581 33241 35584
rect 33275 35581 33287 35615
rect 33229 35575 33287 35581
rect 31904 35516 31984 35544
rect 31904 35504 31910 35516
rect 32030 35504 32036 35556
rect 32088 35544 32094 35556
rect 32217 35547 32275 35553
rect 32217 35544 32229 35547
rect 32088 35516 32229 35544
rect 32088 35504 32094 35516
rect 32217 35513 32229 35516
rect 32263 35513 32275 35547
rect 32217 35507 32275 35513
rect 32766 35504 32772 35556
rect 32824 35504 32830 35556
rect 29564 35448 31156 35476
rect 31570 35436 31576 35488
rect 31628 35436 31634 35488
rect 33042 35436 33048 35488
rect 33100 35476 33106 35488
rect 33428 35476 33456 35643
rect 33594 35640 33600 35692
rect 33652 35640 33658 35692
rect 33704 35689 33732 35720
rect 33962 35708 33968 35720
rect 34020 35708 34026 35760
rect 34054 35708 34060 35760
rect 34112 35748 34118 35760
rect 34422 35748 34428 35760
rect 34112 35720 34428 35748
rect 34112 35708 34118 35720
rect 34422 35708 34428 35720
rect 34480 35708 34486 35760
rect 33689 35683 33747 35689
rect 33689 35649 33701 35683
rect 33735 35649 33747 35683
rect 33689 35643 33747 35649
rect 33965 35615 34023 35621
rect 33965 35612 33977 35615
rect 33612 35584 33977 35612
rect 33612 35553 33640 35584
rect 33965 35581 33977 35584
rect 34011 35581 34023 35615
rect 33965 35575 34023 35581
rect 33597 35547 33655 35553
rect 33597 35513 33609 35547
rect 33643 35513 33655 35547
rect 33597 35507 33655 35513
rect 34146 35476 34152 35488
rect 33100 35448 34152 35476
rect 33100 35436 33106 35448
rect 34146 35436 34152 35448
rect 34204 35476 34210 35488
rect 35437 35479 35495 35485
rect 35437 35476 35449 35479
rect 34204 35448 35449 35476
rect 34204 35436 34210 35448
rect 35437 35445 35449 35448
rect 35483 35476 35495 35479
rect 35618 35476 35624 35488
rect 35483 35448 35624 35476
rect 35483 35445 35495 35448
rect 35437 35439 35495 35445
rect 35618 35436 35624 35448
rect 35676 35436 35682 35488
rect 1104 35386 37076 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 37076 35386
rect 1104 35312 37076 35334
rect 11882 35232 11888 35284
rect 11940 35232 11946 35284
rect 16942 35232 16948 35284
rect 17000 35232 17006 35284
rect 19058 35232 19064 35284
rect 19116 35272 19122 35284
rect 19116 35244 19748 35272
rect 19116 35232 19122 35244
rect 11514 35096 11520 35148
rect 11572 35136 11578 35148
rect 13633 35139 13691 35145
rect 13633 35136 13645 35139
rect 11572 35108 13645 35136
rect 11572 35096 11578 35108
rect 13633 35105 13645 35108
rect 13679 35136 13691 35139
rect 14182 35136 14188 35148
rect 13679 35108 14188 35136
rect 13679 35105 13691 35108
rect 13633 35099 13691 35105
rect 14182 35096 14188 35108
rect 14240 35136 14246 35148
rect 15194 35136 15200 35148
rect 14240 35108 15200 35136
rect 14240 35096 14246 35108
rect 15194 35096 15200 35108
rect 15252 35136 15258 35148
rect 17313 35139 17371 35145
rect 17313 35136 17325 35139
rect 15252 35108 17325 35136
rect 15252 35096 15258 35108
rect 17313 35105 17325 35108
rect 17359 35105 17371 35139
rect 17313 35099 17371 35105
rect 17586 35096 17592 35148
rect 17644 35096 17650 35148
rect 18138 35096 18144 35148
rect 18196 35136 18202 35148
rect 19720 35145 19748 35244
rect 19904 35244 22094 35272
rect 19705 35139 19763 35145
rect 18196 35108 18828 35136
rect 18196 35096 18202 35108
rect 12342 34960 12348 35012
rect 12400 34960 12406 35012
rect 13354 34960 13360 35012
rect 13412 34960 13418 35012
rect 15470 34960 15476 35012
rect 15528 34960 15534 35012
rect 15562 34960 15568 35012
rect 15620 35000 15626 35012
rect 18800 35000 18828 35108
rect 19705 35105 19717 35139
rect 19751 35105 19763 35139
rect 19705 35099 19763 35105
rect 19794 35096 19800 35148
rect 19852 35096 19858 35148
rect 18874 35028 18880 35080
rect 18932 35068 18938 35080
rect 19904 35068 19932 35244
rect 18932 35040 19932 35068
rect 18932 35028 18938 35040
rect 19518 35000 19524 35012
rect 15620 34972 15962 35000
rect 18800 34986 19524 35000
rect 18814 34972 19524 34986
rect 15620 34960 15626 34972
rect 15856 34932 15884 34972
rect 16390 34932 16396 34944
rect 15856 34904 16396 34932
rect 16390 34892 16396 34904
rect 16448 34932 16454 34944
rect 18892 34932 18920 34972
rect 19518 34960 19524 34972
rect 19576 34960 19582 35012
rect 16448 34904 18920 34932
rect 16448 34892 16454 34904
rect 19150 34892 19156 34944
rect 19208 34932 19214 34944
rect 19245 34935 19303 34941
rect 19245 34932 19257 34935
rect 19208 34904 19257 34932
rect 19208 34892 19214 34904
rect 19245 34901 19257 34904
rect 19291 34901 19303 34935
rect 19245 34895 19303 34901
rect 19613 34935 19671 34941
rect 19613 34901 19625 34935
rect 19659 34932 19671 34935
rect 20530 34932 20536 34944
rect 19659 34904 20536 34932
rect 19659 34901 19671 34904
rect 19613 34895 19671 34901
rect 20530 34892 20536 34904
rect 20588 34892 20594 34944
rect 22066 34932 22094 35244
rect 25958 35232 25964 35284
rect 26016 35272 26022 35284
rect 26145 35275 26203 35281
rect 26145 35272 26157 35275
rect 26016 35244 26157 35272
rect 26016 35232 26022 35244
rect 26145 35241 26157 35244
rect 26191 35241 26203 35275
rect 26145 35235 26203 35241
rect 26234 35232 26240 35284
rect 26292 35272 26298 35284
rect 26292 35244 28580 35272
rect 26292 35232 26298 35244
rect 25406 35136 25412 35148
rect 24412 35108 25412 35136
rect 24412 35080 24440 35108
rect 25406 35096 25412 35108
rect 25464 35136 25470 35148
rect 27985 35139 28043 35145
rect 27985 35136 27997 35139
rect 25464 35108 27997 35136
rect 25464 35096 25470 35108
rect 27985 35105 27997 35108
rect 28031 35105 28043 35139
rect 27985 35099 28043 35105
rect 28552 35136 28580 35244
rect 29730 35232 29736 35284
rect 29788 35272 29794 35284
rect 31481 35275 31539 35281
rect 31481 35272 31493 35275
rect 29788 35244 31493 35272
rect 29788 35232 29794 35244
rect 31481 35241 31493 35244
rect 31527 35241 31539 35275
rect 31481 35235 31539 35241
rect 33594 35232 33600 35284
rect 33652 35272 33658 35284
rect 35805 35275 35863 35281
rect 35805 35272 35817 35275
rect 33652 35244 35817 35272
rect 33652 35232 33658 35244
rect 35805 35241 35817 35244
rect 35851 35241 35863 35275
rect 35805 35235 35863 35241
rect 28626 35164 28632 35216
rect 28684 35204 28690 35216
rect 31297 35207 31355 35213
rect 28684 35176 31248 35204
rect 28684 35164 28690 35176
rect 29549 35139 29607 35145
rect 29549 35136 29561 35139
rect 28552 35108 29561 35136
rect 24394 35028 24400 35080
rect 24452 35028 24458 35080
rect 28077 35071 28135 35077
rect 28077 35068 28089 35071
rect 28000 35040 28089 35068
rect 24673 35003 24731 35009
rect 24673 34969 24685 35003
rect 24719 35000 24731 35003
rect 24946 35000 24952 35012
rect 24719 34972 24952 35000
rect 24719 34969 24731 34972
rect 24673 34963 24731 34969
rect 24946 34960 24952 34972
rect 25004 34960 25010 35012
rect 25130 34960 25136 35012
rect 25188 34960 25194 35012
rect 25958 34960 25964 35012
rect 26016 35000 26022 35012
rect 27709 35003 27767 35009
rect 26016 34972 26542 35000
rect 26016 34960 26022 34972
rect 27709 34969 27721 35003
rect 27755 35000 27767 35003
rect 28000 35000 28028 35040
rect 28077 35037 28089 35040
rect 28123 35037 28135 35071
rect 28077 35031 28135 35037
rect 28442 35028 28448 35080
rect 28500 35068 28506 35080
rect 28552 35077 28580 35108
rect 29549 35105 29561 35108
rect 29595 35105 29607 35139
rect 29549 35099 29607 35105
rect 28537 35071 28595 35077
rect 28537 35068 28549 35071
rect 28500 35040 28549 35068
rect 28500 35028 28506 35040
rect 28537 35037 28549 35040
rect 28583 35037 28595 35071
rect 28537 35031 28595 35037
rect 28718 35028 28724 35080
rect 28776 35028 28782 35080
rect 28810 35028 28816 35080
rect 28868 35028 28874 35080
rect 29178 35028 29184 35080
rect 29236 35068 29242 35080
rect 29917 35071 29975 35077
rect 29917 35068 29929 35071
rect 29236 35040 29929 35068
rect 29236 35028 29242 35040
rect 29917 35037 29929 35040
rect 29963 35068 29975 35071
rect 30193 35071 30251 35077
rect 30193 35068 30205 35071
rect 29963 35040 30205 35068
rect 29963 35037 29975 35040
rect 29917 35031 29975 35037
rect 30193 35037 30205 35040
rect 30239 35037 30251 35071
rect 30193 35031 30251 35037
rect 30466 35028 30472 35080
rect 30524 35068 30530 35080
rect 30837 35071 30895 35077
rect 30837 35068 30849 35071
rect 30524 35040 30849 35068
rect 30524 35028 30530 35040
rect 30837 35037 30849 35040
rect 30883 35037 30895 35071
rect 31220 35068 31248 35176
rect 31297 35173 31309 35207
rect 31343 35173 31355 35207
rect 31297 35167 31355 35173
rect 31312 35136 31340 35167
rect 31386 35164 31392 35216
rect 31444 35204 31450 35216
rect 31444 35176 33272 35204
rect 31444 35164 31450 35176
rect 31754 35136 31760 35148
rect 31312 35108 31760 35136
rect 31754 35096 31760 35108
rect 31812 35096 31818 35148
rect 31938 35096 31944 35148
rect 31996 35096 32002 35148
rect 32030 35096 32036 35148
rect 32088 35136 32094 35148
rect 32493 35139 32551 35145
rect 32493 35136 32505 35139
rect 32088 35108 32505 35136
rect 32088 35096 32094 35108
rect 32493 35105 32505 35108
rect 32539 35105 32551 35139
rect 32493 35099 32551 35105
rect 32585 35139 32643 35145
rect 32585 35105 32597 35139
rect 32631 35136 32643 35139
rect 32674 35136 32680 35148
rect 32631 35108 32680 35136
rect 32631 35105 32643 35108
rect 32585 35099 32643 35105
rect 31665 35071 31723 35077
rect 31665 35068 31677 35071
rect 31220 35040 31677 35068
rect 30837 35031 30895 35037
rect 31665 35037 31677 35040
rect 31711 35037 31723 35071
rect 31665 35031 31723 35037
rect 29086 35000 29092 35012
rect 27755 34972 28028 35000
rect 28092 34972 29092 35000
rect 27755 34969 27767 34972
rect 27709 34963 27767 34969
rect 28092 34932 28120 34972
rect 29086 34960 29092 34972
rect 29144 34960 29150 35012
rect 29825 35003 29883 35009
rect 29825 35000 29837 35003
rect 29656 34972 29837 35000
rect 22066 34904 28120 34932
rect 28166 34892 28172 34944
rect 28224 34932 28230 34944
rect 29656 34932 29684 34972
rect 29825 34969 29837 34972
rect 29871 34969 29883 35003
rect 29825 34963 29883 34969
rect 28224 34904 29684 34932
rect 29733 34935 29791 34941
rect 28224 34892 28230 34904
rect 29733 34901 29745 34935
rect 29779 34932 29791 34935
rect 30006 34932 30012 34944
rect 29779 34904 30012 34932
rect 29779 34901 29791 34904
rect 29733 34895 29791 34901
rect 30006 34892 30012 34904
rect 30064 34892 30070 34944
rect 30098 34892 30104 34944
rect 30156 34892 30162 34944
rect 30650 34892 30656 34944
rect 30708 34892 30714 34944
rect 31680 34932 31708 35031
rect 31846 35028 31852 35080
rect 31904 35028 31910 35080
rect 32122 35028 32128 35080
rect 32180 35068 32186 35080
rect 32217 35071 32275 35077
rect 32217 35068 32229 35071
rect 32180 35040 32229 35068
rect 32180 35028 32186 35040
rect 32217 35037 32229 35040
rect 32263 35037 32275 35071
rect 32217 35031 32275 35037
rect 32030 34960 32036 35012
rect 32088 35000 32094 35012
rect 32600 35000 32628 35099
rect 32674 35096 32680 35108
rect 32732 35096 32738 35148
rect 33244 35136 33272 35176
rect 33318 35164 33324 35216
rect 33376 35204 33382 35216
rect 34333 35207 34391 35213
rect 34333 35204 34345 35207
rect 33376 35176 34345 35204
rect 33376 35164 33382 35176
rect 34333 35173 34345 35176
rect 34379 35173 34391 35207
rect 34333 35167 34391 35173
rect 33244 35108 33364 35136
rect 33336 35080 33364 35108
rect 33502 35096 33508 35148
rect 33560 35096 33566 35148
rect 33870 35096 33876 35148
rect 33928 35096 33934 35148
rect 33137 35071 33195 35077
rect 33137 35037 33149 35071
rect 33183 35068 33195 35071
rect 33226 35068 33232 35080
rect 33183 35040 33232 35068
rect 33183 35037 33195 35040
rect 33137 35031 33195 35037
rect 33226 35028 33232 35040
rect 33284 35028 33290 35080
rect 33318 35028 33324 35080
rect 33376 35028 33382 35080
rect 33594 35028 33600 35080
rect 33652 35028 33658 35080
rect 33689 35071 33747 35077
rect 33689 35037 33701 35071
rect 33735 35037 33747 35071
rect 33689 35031 33747 35037
rect 32088 34972 32628 35000
rect 32088 34960 32094 34972
rect 33042 34960 33048 35012
rect 33100 35000 33106 35012
rect 33704 35000 33732 35031
rect 34790 35028 34796 35080
rect 34848 35028 34854 35080
rect 35526 35028 35532 35080
rect 35584 35028 35590 35080
rect 35618 35028 35624 35080
rect 35676 35028 35682 35080
rect 36081 35071 36139 35077
rect 36081 35068 36093 35071
rect 35728 35040 36093 35068
rect 33100 34972 33732 35000
rect 35161 35003 35219 35009
rect 33100 34960 33106 34972
rect 35161 34969 35173 35003
rect 35207 35000 35219 35003
rect 35728 35000 35756 35040
rect 36081 35037 36093 35040
rect 36127 35037 36139 35071
rect 36081 35031 36139 35037
rect 35207 34972 35756 35000
rect 35805 35003 35863 35009
rect 35207 34969 35219 34972
rect 35161 34963 35219 34969
rect 35805 34969 35817 35003
rect 35851 34969 35863 35003
rect 35805 34963 35863 34969
rect 31846 34932 31852 34944
rect 31680 34904 31852 34932
rect 31846 34892 31852 34904
rect 31904 34892 31910 34944
rect 33594 34892 33600 34944
rect 33652 34932 33658 34944
rect 35176 34932 35204 34963
rect 33652 34904 35204 34932
rect 35820 34932 35848 34963
rect 35897 34935 35955 34941
rect 35897 34932 35909 34935
rect 35820 34904 35909 34932
rect 33652 34892 33658 34904
rect 35897 34901 35909 34904
rect 35943 34901 35955 34935
rect 35897 34895 35955 34901
rect 1104 34842 37076 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 37076 34842
rect 1104 34768 37076 34790
rect 11882 34688 11888 34740
rect 11940 34728 11946 34740
rect 12345 34731 12403 34737
rect 12345 34728 12357 34731
rect 11940 34700 12357 34728
rect 11940 34688 11946 34700
rect 12345 34697 12357 34700
rect 12391 34697 12403 34731
rect 12345 34691 12403 34697
rect 15933 34731 15991 34737
rect 15933 34697 15945 34731
rect 15979 34728 15991 34731
rect 16206 34728 16212 34740
rect 15979 34700 16212 34728
rect 15979 34697 15991 34700
rect 15933 34691 15991 34697
rect 16206 34688 16212 34700
rect 16264 34728 16270 34740
rect 18874 34728 18880 34740
rect 16264 34700 16574 34728
rect 16264 34688 16270 34700
rect 12253 34663 12311 34669
rect 12253 34629 12265 34663
rect 12299 34660 12311 34663
rect 13173 34663 13231 34669
rect 13173 34660 13185 34663
rect 12299 34632 13185 34660
rect 12299 34629 12311 34632
rect 12253 34623 12311 34629
rect 13173 34629 13185 34632
rect 13219 34660 13231 34663
rect 13538 34660 13544 34672
rect 13219 34632 13544 34660
rect 13219 34629 13231 34632
rect 13173 34623 13231 34629
rect 13538 34620 13544 34632
rect 13596 34620 13602 34672
rect 16546 34660 16574 34700
rect 17144 34700 18880 34728
rect 16546 34632 16988 34660
rect 13078 34552 13084 34604
rect 13136 34552 13142 34604
rect 14182 34552 14188 34604
rect 14240 34552 14246 34604
rect 15562 34552 15568 34604
rect 15620 34552 15626 34604
rect 12529 34527 12587 34533
rect 12529 34493 12541 34527
rect 12575 34493 12587 34527
rect 12529 34487 12587 34493
rect 12544 34456 12572 34487
rect 13354 34484 13360 34536
rect 13412 34484 13418 34536
rect 16669 34527 16727 34533
rect 16669 34524 16681 34527
rect 16546 34496 16681 34524
rect 13814 34456 13820 34468
rect 12544 34428 13820 34456
rect 13814 34416 13820 34428
rect 13872 34416 13878 34468
rect 16546 34456 16574 34496
rect 16669 34493 16681 34496
rect 16715 34493 16727 34527
rect 16960 34524 16988 34632
rect 17144 34601 17172 34700
rect 18874 34688 18880 34700
rect 18932 34688 18938 34740
rect 19794 34688 19800 34740
rect 19852 34728 19858 34740
rect 19852 34700 20484 34728
rect 19852 34688 19858 34700
rect 19334 34660 19340 34672
rect 17236 34632 17448 34660
rect 17129 34595 17187 34601
rect 17129 34561 17141 34595
rect 17175 34561 17187 34595
rect 17129 34555 17187 34561
rect 17236 34524 17264 34632
rect 17420 34601 17448 34632
rect 18800 34632 19340 34660
rect 18800 34601 18828 34632
rect 19334 34620 19340 34632
rect 19392 34620 19398 34672
rect 19518 34620 19524 34672
rect 19576 34620 19582 34672
rect 20456 34660 20484 34700
rect 20530 34688 20536 34740
rect 20588 34688 20594 34740
rect 25409 34731 25467 34737
rect 25409 34697 25421 34731
rect 25455 34728 25467 34731
rect 25498 34728 25504 34740
rect 25455 34700 25504 34728
rect 25455 34697 25467 34700
rect 25409 34691 25467 34697
rect 25498 34688 25504 34700
rect 25556 34688 25562 34740
rect 27893 34731 27951 34737
rect 27893 34697 27905 34731
rect 27939 34697 27951 34731
rect 27893 34691 27951 34697
rect 24670 34660 24676 34672
rect 20456 34632 24676 34660
rect 24670 34620 24676 34632
rect 24728 34620 24734 34672
rect 25222 34620 25228 34672
rect 25280 34660 25286 34672
rect 25958 34660 25964 34672
rect 25280 34632 25964 34660
rect 25280 34620 25286 34632
rect 25958 34620 25964 34632
rect 26016 34620 26022 34672
rect 27525 34663 27583 34669
rect 27525 34629 27537 34663
rect 27571 34660 27583 34663
rect 27614 34660 27620 34672
rect 27571 34632 27620 34660
rect 27571 34629 27583 34632
rect 27525 34623 27583 34629
rect 27614 34620 27620 34632
rect 27672 34620 27678 34672
rect 27798 34669 27804 34672
rect 27741 34663 27804 34669
rect 27741 34629 27753 34663
rect 27787 34629 27804 34663
rect 27741 34623 27804 34629
rect 27798 34620 27804 34623
rect 27856 34620 27862 34672
rect 27908 34660 27936 34691
rect 28442 34688 28448 34740
rect 28500 34688 28506 34740
rect 28537 34731 28595 34737
rect 28537 34697 28549 34731
rect 28583 34728 28595 34731
rect 30650 34728 30656 34740
rect 28583 34700 30656 34728
rect 28583 34697 28595 34700
rect 28537 34691 28595 34697
rect 30650 34688 30656 34700
rect 30708 34688 30714 34740
rect 31846 34688 31852 34740
rect 31904 34728 31910 34740
rect 32214 34728 32220 34740
rect 31904 34700 32220 34728
rect 31904 34688 31910 34700
rect 32214 34688 32220 34700
rect 32272 34728 32278 34740
rect 32401 34731 32459 34737
rect 32401 34728 32413 34731
rect 32272 34700 32413 34728
rect 32272 34688 32278 34700
rect 32401 34697 32413 34700
rect 32447 34697 32459 34731
rect 32401 34691 32459 34697
rect 32585 34731 32643 34737
rect 32585 34697 32597 34731
rect 32631 34728 32643 34731
rect 33226 34728 33232 34740
rect 32631 34700 33232 34728
rect 32631 34697 32643 34700
rect 32585 34691 32643 34697
rect 33226 34688 33232 34700
rect 33284 34688 33290 34740
rect 33321 34731 33379 34737
rect 33321 34697 33333 34731
rect 33367 34728 33379 34731
rect 33410 34728 33416 34740
rect 33367 34700 33416 34728
rect 33367 34697 33379 34700
rect 33321 34691 33379 34697
rect 33410 34688 33416 34700
rect 33468 34688 33474 34740
rect 33597 34731 33655 34737
rect 33597 34697 33609 34731
rect 33643 34728 33655 34731
rect 34606 34728 34612 34740
rect 33643 34700 34612 34728
rect 33643 34697 33655 34700
rect 33597 34691 33655 34697
rect 34606 34688 34612 34700
rect 34664 34688 34670 34740
rect 29454 34660 29460 34672
rect 27908 34632 29460 34660
rect 29454 34620 29460 34632
rect 29512 34620 29518 34672
rect 31662 34660 31668 34672
rect 30944 34632 31668 34660
rect 30944 34604 30972 34632
rect 31662 34620 31668 34632
rect 31720 34620 31726 34672
rect 33042 34660 33048 34672
rect 32692 34632 33048 34660
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34561 17371 34595
rect 17313 34555 17371 34561
rect 17405 34595 17463 34601
rect 17405 34561 17417 34595
rect 17451 34561 17463 34595
rect 17405 34555 17463 34561
rect 18785 34595 18843 34601
rect 18785 34561 18797 34595
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 16960 34496 17264 34524
rect 17328 34524 17356 34555
rect 20622 34552 20628 34604
rect 20680 34552 20686 34604
rect 22465 34595 22523 34601
rect 22465 34561 22477 34595
rect 22511 34592 22523 34595
rect 23474 34592 23480 34604
rect 22511 34564 23480 34592
rect 22511 34561 22523 34564
rect 22465 34555 22523 34561
rect 23474 34552 23480 34564
rect 23532 34552 23538 34604
rect 25501 34595 25559 34601
rect 25501 34561 25513 34595
rect 25547 34592 25559 34595
rect 26142 34592 26148 34604
rect 25547 34564 26148 34592
rect 25547 34561 25559 34564
rect 25501 34555 25559 34561
rect 26142 34552 26148 34564
rect 26200 34552 26206 34604
rect 27985 34595 28043 34601
rect 27985 34561 27997 34595
rect 28031 34592 28043 34595
rect 28902 34592 28908 34604
rect 28031 34564 28908 34592
rect 28031 34561 28043 34564
rect 27985 34555 28043 34561
rect 28902 34552 28908 34564
rect 28960 34552 28966 34604
rect 29362 34552 29368 34604
rect 29420 34552 29426 34604
rect 29549 34595 29607 34601
rect 29549 34561 29561 34595
rect 29595 34592 29607 34595
rect 30098 34592 30104 34604
rect 29595 34564 30104 34592
rect 29595 34561 29607 34564
rect 29549 34555 29607 34561
rect 17770 34524 17776 34536
rect 17328 34496 17776 34524
rect 16669 34487 16727 34493
rect 17770 34484 17776 34496
rect 17828 34484 17834 34536
rect 19061 34527 19119 34533
rect 19061 34493 19073 34527
rect 19107 34524 19119 34527
rect 19150 34524 19156 34536
rect 19107 34496 19156 34524
rect 19107 34493 19119 34496
rect 19061 34487 19119 34493
rect 19150 34484 19156 34496
rect 19208 34484 19214 34536
rect 22554 34484 22560 34536
rect 22612 34484 22618 34536
rect 22741 34527 22799 34533
rect 22741 34493 22753 34527
rect 22787 34493 22799 34527
rect 22741 34487 22799 34493
rect 25685 34527 25743 34533
rect 25685 34493 25697 34527
rect 25731 34493 25743 34527
rect 25685 34487 25743 34493
rect 22756 34456 22784 34487
rect 24854 34456 24860 34468
rect 15856 34428 16574 34456
rect 21468 34428 24860 34456
rect 11885 34391 11943 34397
rect 11885 34357 11897 34391
rect 11931 34388 11943 34391
rect 12066 34388 12072 34400
rect 11931 34360 12072 34388
rect 11931 34357 11943 34360
rect 11885 34351 11943 34357
rect 12066 34348 12072 34360
rect 12124 34348 12130 34400
rect 12710 34348 12716 34400
rect 12768 34348 12774 34400
rect 14448 34391 14506 34397
rect 14448 34357 14460 34391
rect 14494 34388 14506 34391
rect 15856 34388 15884 34428
rect 21468 34400 21496 34428
rect 24854 34416 24860 34428
rect 24912 34456 24918 34468
rect 25700 34456 25728 34487
rect 28166 34484 28172 34536
rect 28224 34484 28230 34536
rect 28258 34484 28264 34536
rect 28316 34484 28322 34536
rect 28629 34527 28687 34533
rect 28629 34493 28641 34527
rect 28675 34524 28687 34527
rect 28994 34524 29000 34536
rect 28675 34496 28764 34524
rect 28675 34493 28687 34496
rect 28629 34487 28687 34493
rect 25774 34456 25780 34468
rect 24912 34428 25780 34456
rect 24912 34416 24918 34428
rect 25774 34416 25780 34428
rect 25832 34416 25838 34468
rect 28736 34456 28764 34496
rect 28920 34496 29000 34524
rect 28920 34456 28948 34496
rect 28994 34484 29000 34496
rect 29052 34484 29058 34536
rect 29086 34484 29092 34536
rect 29144 34484 29150 34536
rect 29270 34484 29276 34536
rect 29328 34524 29334 34536
rect 29564 34524 29592 34555
rect 30098 34552 30104 34564
rect 30156 34552 30162 34604
rect 30466 34552 30472 34604
rect 30524 34552 30530 34604
rect 30926 34552 30932 34604
rect 30984 34552 30990 34604
rect 31570 34552 31576 34604
rect 31628 34552 31634 34604
rect 31938 34552 31944 34604
rect 31996 34592 32002 34604
rect 32214 34592 32220 34604
rect 31996 34564 32220 34592
rect 31996 34552 32002 34564
rect 32214 34552 32220 34564
rect 32272 34552 32278 34604
rect 32309 34595 32367 34601
rect 32309 34561 32321 34595
rect 32355 34592 32367 34595
rect 32490 34592 32496 34604
rect 32355 34564 32496 34592
rect 32355 34561 32367 34564
rect 32309 34555 32367 34561
rect 32490 34552 32496 34564
rect 32548 34552 32554 34604
rect 32692 34601 32720 34632
rect 33042 34620 33048 34632
rect 33100 34620 33106 34672
rect 34514 34620 34520 34672
rect 34572 34660 34578 34672
rect 34572 34632 34730 34660
rect 34572 34620 34578 34632
rect 32677 34595 32735 34601
rect 32677 34561 32689 34595
rect 32723 34561 32735 34595
rect 32677 34555 32735 34561
rect 33226 34552 33232 34604
rect 33284 34552 33290 34604
rect 33410 34552 33416 34604
rect 33468 34552 33474 34604
rect 33686 34552 33692 34604
rect 33744 34552 33750 34604
rect 33962 34552 33968 34604
rect 34020 34552 34026 34604
rect 29328 34496 29592 34524
rect 29328 34484 29334 34496
rect 29730 34484 29736 34536
rect 29788 34524 29794 34536
rect 29825 34527 29883 34533
rect 29825 34524 29837 34527
rect 29788 34496 29837 34524
rect 29788 34484 29794 34496
rect 29825 34493 29837 34496
rect 29871 34493 29883 34527
rect 29825 34487 29883 34493
rect 30006 34484 30012 34536
rect 30064 34524 30070 34536
rect 30484 34524 30512 34552
rect 30064 34496 30512 34524
rect 30064 34484 30070 34496
rect 30558 34484 30564 34536
rect 30616 34524 30622 34536
rect 32030 34524 32036 34536
rect 30616 34496 32036 34524
rect 30616 34484 30622 34496
rect 32030 34484 32036 34496
rect 32088 34484 32094 34536
rect 32769 34527 32827 34533
rect 32769 34493 32781 34527
rect 32815 34524 32827 34527
rect 33428 34524 33456 34552
rect 32815 34496 33456 34524
rect 33781 34527 33839 34533
rect 32815 34493 32827 34496
rect 32769 34487 32827 34493
rect 33781 34493 33793 34527
rect 33827 34524 33839 34527
rect 34241 34527 34299 34533
rect 34241 34524 34253 34527
rect 33827 34496 34253 34524
rect 33827 34493 33839 34496
rect 33781 34487 33839 34493
rect 34241 34493 34253 34496
rect 34287 34493 34299 34527
rect 34241 34487 34299 34493
rect 34330 34484 34336 34536
rect 34388 34524 34394 34536
rect 35713 34527 35771 34533
rect 35713 34524 35725 34527
rect 34388 34496 35725 34524
rect 34388 34484 34394 34496
rect 35713 34493 35725 34496
rect 35759 34493 35771 34527
rect 35713 34487 35771 34493
rect 28736 34428 28948 34456
rect 33226 34416 33232 34468
rect 33284 34456 33290 34468
rect 33284 34428 33640 34456
rect 33284 34416 33290 34428
rect 14494 34360 15884 34388
rect 14494 34357 14506 34360
rect 14448 34351 14506 34357
rect 19610 34348 19616 34400
rect 19668 34388 19674 34400
rect 21450 34388 21456 34400
rect 19668 34360 21456 34388
rect 19668 34348 19674 34360
rect 21450 34348 21456 34360
rect 21508 34348 21514 34400
rect 22094 34348 22100 34400
rect 22152 34348 22158 34400
rect 25038 34348 25044 34400
rect 25096 34348 25102 34400
rect 27709 34391 27767 34397
rect 27709 34357 27721 34391
rect 27755 34388 27767 34391
rect 30282 34388 30288 34400
rect 27755 34360 30288 34388
rect 27755 34357 27767 34360
rect 27709 34351 27767 34357
rect 30282 34348 30288 34360
rect 30340 34348 30346 34400
rect 30466 34348 30472 34400
rect 30524 34388 30530 34400
rect 30561 34391 30619 34397
rect 30561 34388 30573 34391
rect 30524 34360 30573 34388
rect 30524 34348 30530 34360
rect 30561 34357 30573 34360
rect 30607 34357 30619 34391
rect 30561 34351 30619 34357
rect 32953 34391 33011 34397
rect 32953 34357 32965 34391
rect 32999 34388 33011 34391
rect 33042 34388 33048 34400
rect 32999 34360 33048 34388
rect 32999 34357 33011 34360
rect 32953 34351 33011 34357
rect 33042 34348 33048 34360
rect 33100 34348 33106 34400
rect 33612 34388 33640 34428
rect 34054 34388 34060 34400
rect 33612 34360 34060 34388
rect 34054 34348 34060 34360
rect 34112 34388 34118 34400
rect 34330 34388 34336 34400
rect 34112 34360 34336 34388
rect 34112 34348 34118 34360
rect 34330 34348 34336 34360
rect 34388 34348 34394 34400
rect 1104 34298 37076 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 37076 34298
rect 1104 34224 37076 34246
rect 13538 34144 13544 34196
rect 13596 34144 13602 34196
rect 14274 34144 14280 34196
rect 14332 34184 14338 34196
rect 17589 34187 17647 34193
rect 17589 34184 17601 34187
rect 14332 34156 17601 34184
rect 14332 34144 14338 34156
rect 17589 34153 17601 34156
rect 17635 34153 17647 34187
rect 17589 34147 17647 34153
rect 23293 34187 23351 34193
rect 23293 34153 23305 34187
rect 23339 34184 23351 34187
rect 23474 34184 23480 34196
rect 23339 34156 23480 34184
rect 23339 34153 23351 34156
rect 23293 34147 23351 34153
rect 23474 34144 23480 34156
rect 23532 34144 23538 34196
rect 28166 34144 28172 34196
rect 28224 34184 28230 34196
rect 28445 34187 28503 34193
rect 28445 34184 28457 34187
rect 28224 34156 28457 34184
rect 28224 34144 28230 34156
rect 28445 34153 28457 34156
rect 28491 34153 28503 34187
rect 28445 34147 28503 34153
rect 29089 34187 29147 34193
rect 29089 34153 29101 34187
rect 29135 34184 29147 34187
rect 30006 34184 30012 34196
rect 29135 34156 30012 34184
rect 29135 34153 29147 34156
rect 29089 34147 29147 34153
rect 30006 34144 30012 34156
rect 30064 34144 30070 34196
rect 31938 34184 31944 34196
rect 30852 34156 31944 34184
rect 29362 34076 29368 34128
rect 29420 34116 29426 34128
rect 29420 34088 29960 34116
rect 29420 34076 29426 34088
rect 11514 34008 11520 34060
rect 11572 34048 11578 34060
rect 11793 34051 11851 34057
rect 11793 34048 11805 34051
rect 11572 34020 11805 34048
rect 11572 34008 11578 34020
rect 11793 34017 11805 34020
rect 11839 34017 11851 34051
rect 11793 34011 11851 34017
rect 12066 34008 12072 34060
rect 12124 34008 12130 34060
rect 14182 34008 14188 34060
rect 14240 34048 14246 34060
rect 14737 34051 14795 34057
rect 14737 34048 14749 34051
rect 14240 34020 14749 34048
rect 14240 34008 14246 34020
rect 14737 34017 14749 34020
rect 14783 34017 14795 34051
rect 14737 34011 14795 34017
rect 14752 33980 14780 34011
rect 15562 34008 15568 34060
rect 15620 34048 15626 34060
rect 15620 34020 19288 34048
rect 15620 34008 15626 34020
rect 15657 33983 15715 33989
rect 15657 33980 15669 33983
rect 14752 33952 15669 33980
rect 15657 33949 15669 33952
rect 15703 33949 15715 33983
rect 15657 33943 15715 33949
rect 18141 33983 18199 33989
rect 18141 33949 18153 33983
rect 18187 33980 18199 33983
rect 18874 33980 18880 33992
rect 18187 33952 18880 33980
rect 18187 33949 18199 33952
rect 18141 33943 18199 33949
rect 18874 33940 18880 33952
rect 18932 33940 18938 33992
rect 15378 33912 15384 33924
rect 13294 33884 15384 33912
rect 12342 33804 12348 33856
rect 12400 33844 12406 33856
rect 13372 33844 13400 33884
rect 15378 33872 15384 33884
rect 15436 33872 15442 33924
rect 15562 33872 15568 33924
rect 15620 33872 15626 33924
rect 15930 33872 15936 33924
rect 15988 33872 15994 33924
rect 16390 33872 16396 33924
rect 16448 33872 16454 33924
rect 17770 33872 17776 33924
rect 17828 33912 17834 33924
rect 17865 33915 17923 33921
rect 17865 33912 17877 33915
rect 17828 33884 17877 33912
rect 17828 33872 17834 33884
rect 17865 33881 17877 33884
rect 17911 33881 17923 33915
rect 19260 33912 19288 34020
rect 19334 34008 19340 34060
rect 19392 34048 19398 34060
rect 19978 34048 19984 34060
rect 19392 34020 19984 34048
rect 19392 34008 19398 34020
rect 19978 34008 19984 34020
rect 20036 34048 20042 34060
rect 20622 34048 20628 34060
rect 20036 34020 20628 34048
rect 20036 34008 20042 34020
rect 20622 34008 20628 34020
rect 20680 34048 20686 34060
rect 24673 34051 24731 34057
rect 20680 34020 21588 34048
rect 20680 34008 20686 34020
rect 21560 33992 21588 34020
rect 24673 34017 24685 34051
rect 24719 34048 24731 34051
rect 25038 34048 25044 34060
rect 24719 34020 25044 34048
rect 24719 34017 24731 34020
rect 24673 34011 24731 34017
rect 25038 34008 25044 34020
rect 25096 34008 25102 34060
rect 25130 34008 25136 34060
rect 25188 34048 25194 34060
rect 26697 34051 26755 34057
rect 26697 34048 26709 34051
rect 25188 34020 26709 34048
rect 25188 34008 25194 34020
rect 26697 34017 26709 34020
rect 26743 34017 26755 34051
rect 26697 34011 26755 34017
rect 26973 34051 27031 34057
rect 26973 34017 26985 34051
rect 27019 34048 27031 34051
rect 28534 34048 28540 34060
rect 27019 34020 28540 34048
rect 27019 34017 27031 34020
rect 26973 34011 27031 34017
rect 28534 34008 28540 34020
rect 28592 34008 28598 34060
rect 29178 34008 29184 34060
rect 29236 34048 29242 34060
rect 29825 34051 29883 34057
rect 29825 34048 29837 34051
rect 29236 34020 29837 34048
rect 29236 34008 29242 34020
rect 29825 34017 29837 34020
rect 29871 34017 29883 34051
rect 29825 34011 29883 34017
rect 21542 33940 21548 33992
rect 21600 33940 21606 33992
rect 24394 33940 24400 33992
rect 24452 33940 24458 33992
rect 29270 33940 29276 33992
rect 29328 33940 29334 33992
rect 29362 33940 29368 33992
rect 29420 33940 29426 33992
rect 29549 33983 29607 33989
rect 29549 33949 29561 33983
rect 29595 33980 29607 33983
rect 29932 33980 29960 34088
rect 30852 33980 30880 34156
rect 31938 34144 31944 34156
rect 31996 34184 32002 34196
rect 33229 34187 33287 34193
rect 31996 34156 32812 34184
rect 31996 34144 32002 34156
rect 32784 34116 32812 34156
rect 33229 34153 33241 34187
rect 33275 34184 33287 34187
rect 33410 34184 33416 34196
rect 33275 34156 33416 34184
rect 33275 34153 33287 34156
rect 33229 34147 33287 34153
rect 33410 34144 33416 34156
rect 33468 34144 33474 34196
rect 32784 34088 33548 34116
rect 31478 34008 31484 34060
rect 31536 34048 31542 34060
rect 32766 34048 32772 34060
rect 31536 34020 32772 34048
rect 31536 34008 31542 34020
rect 32766 34008 32772 34020
rect 32824 34008 32830 34060
rect 29595 33952 30880 33980
rect 31113 33983 31171 33989
rect 29595 33949 29607 33952
rect 29549 33943 29607 33949
rect 31113 33949 31125 33983
rect 31159 33980 31171 33983
rect 31294 33980 31300 33992
rect 31159 33952 31300 33980
rect 31159 33949 31171 33952
rect 31113 33943 31171 33949
rect 31294 33940 31300 33952
rect 31352 33940 31358 33992
rect 33520 33989 33548 34088
rect 34606 34008 34612 34060
rect 34664 34048 34670 34060
rect 35253 34051 35311 34057
rect 35253 34048 35265 34051
rect 34664 34020 35265 34048
rect 34664 34008 34670 34020
rect 35253 34017 35265 34020
rect 35299 34017 35311 34051
rect 35253 34011 35311 34017
rect 35636 34020 35940 34048
rect 33505 33983 33563 33989
rect 33505 33949 33517 33983
rect 33551 33949 33563 33983
rect 33505 33943 33563 33949
rect 34330 33940 34336 33992
rect 34388 33940 34394 33992
rect 35268 33980 35296 34011
rect 35636 33989 35664 34020
rect 35621 33983 35679 33989
rect 35621 33980 35633 33983
rect 35268 33952 35633 33980
rect 35621 33949 35633 33952
rect 35667 33949 35679 33983
rect 35621 33943 35679 33949
rect 35710 33940 35716 33992
rect 35768 33940 35774 33992
rect 35912 33989 35940 34020
rect 35897 33983 35955 33989
rect 35897 33949 35909 33983
rect 35943 33949 35955 33983
rect 35897 33943 35955 33949
rect 19518 33912 19524 33924
rect 19260 33884 19524 33912
rect 17865 33875 17923 33881
rect 19518 33872 19524 33884
rect 19576 33872 19582 33924
rect 19613 33915 19671 33921
rect 19613 33881 19625 33915
rect 19659 33912 19671 33915
rect 19702 33912 19708 33924
rect 19659 33884 19708 33912
rect 19659 33881 19671 33884
rect 19613 33875 19671 33881
rect 19702 33872 19708 33884
rect 19760 33872 19766 33924
rect 21266 33912 21272 33924
rect 20838 33884 21272 33912
rect 21266 33872 21272 33884
rect 21324 33872 21330 33924
rect 21821 33915 21879 33921
rect 21821 33881 21833 33915
rect 21867 33912 21879 33915
rect 22094 33912 22100 33924
rect 21867 33884 22100 33912
rect 21867 33881 21879 33884
rect 21821 33875 21879 33881
rect 22094 33872 22100 33884
rect 22152 33872 22158 33924
rect 22204 33884 22310 33912
rect 12400 33816 13400 33844
rect 12400 33804 12406 33816
rect 17402 33804 17408 33856
rect 17460 33844 17466 33856
rect 18049 33847 18107 33853
rect 18049 33844 18061 33847
rect 17460 33816 18061 33844
rect 17460 33804 17466 33816
rect 18049 33813 18061 33816
rect 18095 33813 18107 33847
rect 18049 33807 18107 33813
rect 20622 33804 20628 33856
rect 20680 33844 20686 33856
rect 21085 33847 21143 33853
rect 21085 33844 21097 33847
rect 20680 33816 21097 33844
rect 20680 33804 20686 33816
rect 21085 33813 21097 33816
rect 21131 33813 21143 33847
rect 21284 33844 21312 33872
rect 22204 33856 22232 33884
rect 25222 33872 25228 33924
rect 25280 33872 25286 33924
rect 25958 33872 25964 33924
rect 26016 33912 26022 33924
rect 26016 33884 27462 33912
rect 26016 33872 26022 33884
rect 22186 33844 22192 33856
rect 21284 33816 22192 33844
rect 21085 33807 21143 33813
rect 22186 33804 22192 33816
rect 22244 33804 22250 33856
rect 25498 33804 25504 33856
rect 25556 33844 25562 33856
rect 26145 33847 26203 33853
rect 26145 33844 26157 33847
rect 25556 33816 26157 33844
rect 25556 33804 25562 33816
rect 26145 33813 26157 33816
rect 26191 33813 26203 33847
rect 27356 33844 27384 33884
rect 29638 33872 29644 33924
rect 29696 33912 29702 33924
rect 30561 33915 30619 33921
rect 30561 33912 30573 33915
rect 29696 33884 30573 33912
rect 29696 33872 29702 33884
rect 30561 33881 30573 33884
rect 30607 33881 30619 33915
rect 30561 33875 30619 33881
rect 31764 33915 31822 33921
rect 31764 33881 31776 33915
rect 31810 33912 31822 33915
rect 34514 33912 34520 33924
rect 31810 33884 31892 33912
rect 32982 33884 34520 33912
rect 31810 33881 31822 33884
rect 31764 33875 31822 33881
rect 30374 33844 30380 33856
rect 27356 33816 30380 33844
rect 26145 33807 26203 33813
rect 30374 33804 30380 33816
rect 30432 33844 30438 33856
rect 30650 33844 30656 33856
rect 30432 33816 30656 33844
rect 30432 33804 30438 33816
rect 30650 33804 30656 33816
rect 30708 33804 30714 33856
rect 31864 33844 31892 33884
rect 34514 33872 34520 33884
rect 34572 33872 34578 33924
rect 35250 33872 35256 33924
rect 35308 33912 35314 33924
rect 35805 33915 35863 33921
rect 35805 33912 35817 33915
rect 35308 33884 35817 33912
rect 35308 33872 35314 33884
rect 35805 33881 35817 33884
rect 35851 33881 35863 33915
rect 35805 33875 35863 33881
rect 34422 33844 34428 33856
rect 31864 33816 34428 33844
rect 34422 33804 34428 33816
rect 34480 33804 34486 33856
rect 34606 33804 34612 33856
rect 34664 33844 34670 33856
rect 34793 33847 34851 33853
rect 34793 33844 34805 33847
rect 34664 33816 34805 33844
rect 34664 33804 34670 33816
rect 34793 33813 34805 33816
rect 34839 33813 34851 33847
rect 34793 33807 34851 33813
rect 35434 33804 35440 33856
rect 35492 33804 35498 33856
rect 1104 33754 37076 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 37076 33754
rect 1104 33680 37076 33702
rect 12710 33640 12716 33652
rect 11808 33612 12716 33640
rect 11808 33581 11836 33612
rect 12710 33600 12716 33612
rect 12768 33600 12774 33652
rect 13078 33600 13084 33652
rect 13136 33640 13142 33652
rect 13265 33643 13323 33649
rect 13265 33640 13277 33643
rect 13136 33612 13277 33640
rect 13136 33600 13142 33612
rect 13265 33609 13277 33612
rect 13311 33609 13323 33643
rect 13265 33603 13323 33609
rect 15749 33643 15807 33649
rect 15749 33609 15761 33643
rect 15795 33609 15807 33643
rect 15749 33603 15807 33609
rect 11793 33575 11851 33581
rect 11793 33541 11805 33575
rect 11839 33541 11851 33575
rect 11793 33535 11851 33541
rect 12342 33532 12348 33584
rect 12400 33532 12406 33584
rect 14274 33532 14280 33584
rect 14332 33532 14338 33584
rect 15764 33572 15792 33603
rect 15930 33600 15936 33652
rect 15988 33640 15994 33652
rect 16669 33643 16727 33649
rect 16669 33640 16681 33643
rect 15988 33612 16681 33640
rect 15988 33600 15994 33612
rect 16669 33609 16681 33612
rect 16715 33609 16727 33643
rect 16669 33603 16727 33609
rect 17037 33643 17095 33649
rect 17037 33609 17049 33643
rect 17083 33640 17095 33643
rect 17402 33640 17408 33652
rect 17083 33612 17408 33640
rect 17083 33609 17095 33612
rect 17037 33603 17095 33609
rect 17402 33600 17408 33612
rect 17460 33600 17466 33652
rect 17678 33600 17684 33652
rect 17736 33640 17742 33652
rect 19610 33640 19616 33652
rect 17736 33612 19616 33640
rect 17736 33600 17742 33612
rect 19610 33600 19616 33612
rect 19668 33600 19674 33652
rect 19702 33600 19708 33652
rect 19760 33600 19766 33652
rect 20165 33643 20223 33649
rect 20165 33609 20177 33643
rect 20211 33640 20223 33643
rect 20438 33640 20444 33652
rect 20211 33612 20444 33640
rect 20211 33609 20223 33612
rect 20165 33603 20223 33609
rect 20438 33600 20444 33612
rect 20496 33600 20502 33652
rect 22189 33643 22247 33649
rect 22189 33609 22201 33643
rect 22235 33640 22247 33643
rect 22554 33640 22560 33652
rect 22235 33612 22560 33640
rect 22235 33609 22247 33612
rect 22189 33603 22247 33609
rect 22554 33600 22560 33612
rect 22612 33600 22618 33652
rect 25222 33640 25228 33652
rect 24412 33612 25228 33640
rect 17770 33572 17776 33584
rect 15764 33544 17776 33572
rect 17770 33532 17776 33544
rect 17828 33532 17834 33584
rect 19518 33532 19524 33584
rect 19576 33572 19582 33584
rect 20346 33572 20352 33584
rect 19576 33544 20352 33572
rect 19576 33532 19582 33544
rect 20346 33532 20352 33544
rect 20404 33572 20410 33584
rect 20533 33575 20591 33581
rect 20533 33572 20545 33575
rect 20404 33544 20545 33572
rect 20404 33532 20410 33544
rect 20533 33541 20545 33544
rect 20579 33541 20591 33575
rect 20533 33535 20591 33541
rect 21361 33575 21419 33581
rect 21361 33541 21373 33575
rect 21407 33572 21419 33575
rect 21542 33572 21548 33584
rect 21407 33544 21548 33572
rect 21407 33541 21419 33544
rect 21361 33535 21419 33541
rect 21542 33532 21548 33544
rect 21600 33572 21606 33584
rect 24412 33572 24440 33612
rect 25222 33600 25228 33612
rect 25280 33600 25286 33652
rect 26142 33600 26148 33652
rect 26200 33640 26206 33652
rect 26329 33643 26387 33649
rect 26329 33640 26341 33643
rect 26200 33612 26341 33640
rect 26200 33600 26206 33612
rect 26329 33609 26341 33612
rect 26375 33609 26387 33643
rect 26329 33603 26387 33609
rect 30392 33612 31754 33640
rect 25130 33572 25136 33584
rect 21600 33544 22692 33572
rect 24150 33544 24440 33572
rect 24596 33544 25136 33572
rect 21600 33532 21606 33544
rect 11514 33464 11520 33516
rect 11572 33464 11578 33516
rect 15378 33464 15384 33516
rect 15436 33504 15442 33516
rect 16390 33504 16396 33516
rect 15436 33476 16396 33504
rect 15436 33464 15442 33476
rect 16390 33464 16396 33476
rect 16448 33464 16454 33516
rect 17034 33464 17040 33516
rect 17092 33504 17098 33516
rect 17129 33507 17187 33513
rect 17129 33504 17141 33507
rect 17092 33476 17141 33504
rect 17092 33464 17098 33476
rect 17129 33473 17141 33476
rect 17175 33504 17187 33507
rect 17865 33507 17923 33513
rect 17865 33504 17877 33507
rect 17175 33476 17877 33504
rect 17175 33473 17187 33476
rect 17129 33467 17187 33473
rect 17865 33473 17877 33476
rect 17911 33473 17923 33507
rect 17865 33467 17923 33473
rect 19702 33464 19708 33516
rect 19760 33504 19766 33516
rect 20073 33507 20131 33513
rect 20073 33504 20085 33507
rect 19760 33476 20085 33504
rect 19760 33464 19766 33476
rect 20073 33473 20085 33476
rect 20119 33504 20131 33507
rect 20622 33504 20628 33516
rect 20119 33476 20628 33504
rect 20119 33473 20131 33476
rect 20073 33467 20131 33473
rect 20622 33464 20628 33476
rect 20680 33464 20686 33516
rect 21450 33464 21456 33516
rect 21508 33504 21514 33516
rect 22664 33513 22692 33544
rect 22649 33507 22707 33513
rect 21508 33476 22416 33504
rect 21508 33464 21514 33476
rect 13906 33396 13912 33448
rect 13964 33436 13970 33448
rect 14001 33439 14059 33445
rect 14001 33436 14013 33439
rect 13964 33408 14013 33436
rect 13964 33396 13970 33408
rect 14001 33405 14013 33408
rect 14047 33405 14059 33439
rect 14001 33399 14059 33405
rect 17313 33439 17371 33445
rect 17313 33405 17325 33439
rect 17359 33405 17371 33439
rect 17313 33399 17371 33405
rect 17328 33368 17356 33399
rect 17678 33396 17684 33448
rect 17736 33396 17742 33448
rect 17773 33439 17831 33445
rect 17773 33405 17785 33439
rect 17819 33436 17831 33439
rect 18046 33436 18052 33448
rect 17819 33408 18052 33436
rect 17819 33405 17831 33408
rect 17773 33399 17831 33405
rect 18046 33396 18052 33408
rect 18104 33396 18110 33448
rect 20254 33396 20260 33448
rect 20312 33396 20318 33448
rect 22278 33396 22284 33448
rect 22336 33396 22342 33448
rect 22388 33445 22416 33476
rect 22649 33473 22661 33507
rect 22695 33473 22707 33507
rect 22649 33467 22707 33473
rect 24394 33464 24400 33516
rect 24452 33504 24458 33516
rect 24596 33513 24624 33544
rect 25130 33532 25136 33544
rect 25188 33532 25194 33584
rect 25240 33572 25268 33600
rect 30392 33584 30420 33612
rect 30374 33572 30380 33584
rect 25240 33544 25346 33572
rect 27908 33544 30380 33572
rect 24581 33507 24639 33513
rect 24581 33504 24593 33507
rect 24452 33476 24593 33504
rect 24452 33464 24458 33476
rect 24581 33473 24593 33476
rect 24627 33473 24639 33507
rect 24581 33467 24639 33473
rect 27706 33464 27712 33516
rect 27764 33504 27770 33516
rect 27908 33513 27936 33544
rect 30374 33532 30380 33544
rect 30432 33532 30438 33584
rect 30650 33532 30656 33584
rect 30708 33532 30714 33584
rect 31726 33572 31754 33612
rect 33042 33600 33048 33652
rect 33100 33640 33106 33652
rect 33100 33612 33640 33640
rect 33100 33600 33106 33612
rect 32125 33575 32183 33581
rect 32125 33572 32137 33575
rect 31726 33544 32137 33572
rect 32125 33541 32137 33544
rect 32171 33541 32183 33575
rect 32125 33535 32183 33541
rect 32766 33532 32772 33584
rect 32824 33572 32830 33584
rect 32861 33575 32919 33581
rect 32861 33572 32873 33575
rect 32824 33544 32873 33572
rect 32824 33532 32830 33544
rect 32861 33541 32873 33544
rect 32907 33572 32919 33575
rect 33612 33572 33640 33612
rect 33686 33600 33692 33652
rect 33744 33640 33750 33652
rect 33781 33643 33839 33649
rect 33781 33640 33793 33643
rect 33744 33612 33793 33640
rect 33744 33600 33750 33612
rect 33781 33609 33793 33612
rect 33827 33609 33839 33643
rect 33781 33603 33839 33609
rect 34422 33600 34428 33652
rect 34480 33600 34486 33652
rect 34698 33600 34704 33652
rect 34756 33600 34762 33652
rect 34577 33575 34635 33581
rect 34577 33572 34589 33575
rect 32907 33544 33272 33572
rect 33612 33544 34589 33572
rect 32907 33541 32919 33544
rect 32861 33535 32919 33541
rect 27893 33507 27951 33513
rect 27893 33504 27905 33507
rect 27764 33476 27905 33504
rect 27764 33464 27770 33476
rect 27893 33473 27905 33476
rect 27939 33473 27951 33507
rect 27893 33467 27951 33473
rect 28169 33507 28227 33513
rect 28169 33473 28181 33507
rect 28215 33504 28227 33507
rect 28261 33507 28319 33513
rect 28261 33504 28273 33507
rect 28215 33476 28273 33504
rect 28215 33473 28227 33476
rect 28169 33467 28227 33473
rect 28261 33473 28273 33476
rect 28307 33473 28319 33507
rect 28261 33467 28319 33473
rect 28721 33507 28779 33513
rect 28721 33473 28733 33507
rect 28767 33473 28779 33507
rect 28721 33467 28779 33473
rect 28905 33507 28963 33513
rect 28905 33473 28917 33507
rect 28951 33473 28963 33507
rect 28905 33467 28963 33473
rect 22373 33439 22431 33445
rect 22373 33405 22385 33439
rect 22419 33405 22431 33439
rect 22373 33399 22431 33405
rect 22922 33396 22928 33448
rect 22980 33396 22986 33448
rect 24854 33396 24860 33448
rect 24912 33396 24918 33448
rect 26050 33396 26056 33448
rect 26108 33436 26114 33448
rect 27065 33439 27123 33445
rect 27065 33436 27077 33439
rect 26108 33408 27077 33436
rect 26108 33396 26114 33408
rect 27065 33405 27077 33408
rect 27111 33405 27123 33439
rect 27065 33399 27123 33405
rect 19794 33368 19800 33380
rect 17328 33340 19800 33368
rect 19794 33328 19800 33340
rect 19852 33328 19858 33380
rect 18233 33303 18291 33309
rect 18233 33269 18245 33303
rect 18279 33300 18291 33303
rect 18506 33300 18512 33312
rect 18279 33272 18512 33300
rect 18279 33269 18291 33272
rect 18233 33263 18291 33269
rect 18506 33260 18512 33272
rect 18564 33260 18570 33312
rect 21082 33260 21088 33312
rect 21140 33300 21146 33312
rect 21821 33303 21879 33309
rect 21821 33300 21833 33303
rect 21140 33272 21833 33300
rect 21140 33260 21146 33272
rect 21821 33269 21833 33272
rect 21867 33269 21879 33303
rect 21821 33263 21879 33269
rect 24394 33260 24400 33312
rect 24452 33260 24458 33312
rect 28074 33260 28080 33312
rect 28132 33260 28138 33312
rect 28736 33300 28764 33467
rect 28920 33368 28948 33467
rect 29362 33464 29368 33516
rect 29420 33464 29426 33516
rect 29454 33464 29460 33516
rect 29512 33464 29518 33516
rect 29638 33464 29644 33516
rect 29696 33464 29702 33516
rect 29822 33464 29828 33516
rect 29880 33464 29886 33516
rect 31386 33464 31392 33516
rect 31444 33504 31450 33516
rect 33244 33513 33272 33544
rect 34577 33541 34589 33544
rect 34623 33541 34635 33575
rect 34716 33572 34744 33600
rect 34793 33575 34851 33581
rect 34793 33572 34805 33575
rect 34716 33544 34805 33572
rect 34577 33535 34635 33541
rect 34793 33541 34805 33544
rect 34839 33541 34851 33575
rect 34793 33535 34851 33541
rect 31665 33507 31723 33513
rect 31665 33504 31677 33507
rect 31444 33476 31677 33504
rect 31444 33464 31450 33476
rect 31665 33473 31677 33476
rect 31711 33473 31723 33507
rect 31665 33467 31723 33473
rect 33229 33507 33287 33513
rect 33229 33473 33241 33507
rect 33275 33473 33287 33507
rect 33229 33467 33287 33473
rect 33502 33464 33508 33516
rect 33560 33504 33566 33516
rect 34241 33507 34299 33513
rect 34241 33504 34253 33507
rect 33560 33476 34253 33504
rect 33560 33464 33566 33476
rect 34241 33473 34253 33476
rect 34287 33473 34299 33507
rect 34241 33467 34299 33473
rect 34698 33464 34704 33516
rect 34756 33504 34762 33516
rect 35069 33507 35127 33513
rect 35069 33504 35081 33507
rect 34756 33476 35081 33504
rect 34756 33464 34762 33476
rect 35069 33473 35081 33476
rect 35115 33473 35127 33507
rect 35069 33467 35127 33473
rect 28997 33439 29055 33445
rect 28997 33405 29009 33439
rect 29043 33436 29055 33439
rect 29086 33436 29092 33448
rect 29043 33408 29092 33436
rect 29043 33405 29055 33408
rect 28997 33399 29055 33405
rect 29086 33396 29092 33408
rect 29144 33436 29150 33448
rect 29380 33436 29408 33464
rect 29144 33408 29408 33436
rect 29472 33436 29500 33464
rect 30101 33439 30159 33445
rect 30101 33436 30113 33439
rect 29472 33408 30113 33436
rect 29144 33396 29150 33408
rect 30101 33405 30113 33408
rect 30147 33405 30159 33439
rect 30101 33399 30159 33405
rect 31570 33396 31576 33448
rect 31628 33396 31634 33448
rect 33594 33396 33600 33448
rect 33652 33436 33658 33448
rect 33965 33439 34023 33445
rect 33965 33436 33977 33439
rect 33652 33408 33977 33436
rect 33652 33396 33658 33408
rect 33965 33405 33977 33408
rect 34011 33405 34023 33439
rect 33965 33399 34023 33405
rect 34054 33396 34060 33448
rect 34112 33396 34118 33448
rect 34146 33396 34152 33448
rect 34204 33396 34210 33448
rect 34790 33396 34796 33448
rect 34848 33436 34854 33448
rect 35250 33436 35256 33448
rect 34848 33408 35256 33436
rect 34848 33396 34854 33408
rect 35250 33396 35256 33408
rect 35308 33396 35314 33448
rect 29457 33371 29515 33377
rect 29457 33368 29469 33371
rect 28920 33340 29469 33368
rect 29457 33337 29469 33340
rect 29503 33337 29515 33371
rect 29457 33331 29515 33337
rect 34514 33328 34520 33380
rect 34572 33368 34578 33380
rect 34885 33371 34943 33377
rect 34885 33368 34897 33371
rect 34572 33340 34897 33368
rect 34572 33328 34578 33340
rect 34885 33337 34897 33340
rect 34931 33337 34943 33371
rect 34885 33331 34943 33337
rect 28994 33300 29000 33312
rect 28736 33272 29000 33300
rect 28994 33260 29000 33272
rect 29052 33260 29058 33312
rect 31849 33303 31907 33309
rect 31849 33269 31861 33303
rect 31895 33300 31907 33303
rect 32398 33300 32404 33312
rect 31895 33272 32404 33300
rect 31895 33269 31907 33272
rect 31849 33263 31907 33269
rect 32398 33260 32404 33272
rect 32456 33260 32462 33312
rect 34606 33260 34612 33312
rect 34664 33260 34670 33312
rect 1104 33210 37076 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 37076 33210
rect 1104 33136 37076 33158
rect 17034 33056 17040 33108
rect 17092 33056 17098 33108
rect 22554 33056 22560 33108
rect 22612 33056 22618 33108
rect 22922 33056 22928 33108
rect 22980 33096 22986 33108
rect 23109 33099 23167 33105
rect 23109 33096 23121 33099
rect 22980 33068 23121 33096
rect 22980 33056 22986 33068
rect 23109 33065 23121 33068
rect 23155 33065 23167 33099
rect 23109 33059 23167 33065
rect 24854 33056 24860 33108
rect 24912 33096 24918 33108
rect 25225 33099 25283 33105
rect 25225 33096 25237 33099
rect 24912 33068 25237 33096
rect 24912 33056 24918 33068
rect 25225 33065 25237 33068
rect 25271 33065 25283 33099
rect 25225 33059 25283 33065
rect 28534 33056 28540 33108
rect 28592 33056 28598 33108
rect 28721 33099 28779 33105
rect 28721 33065 28733 33099
rect 28767 33096 28779 33099
rect 28810 33096 28816 33108
rect 28767 33068 28816 33096
rect 28767 33065 28779 33068
rect 28721 33059 28779 33065
rect 19610 32988 19616 33040
rect 19668 33028 19674 33040
rect 24670 33028 24676 33040
rect 19668 33000 19840 33028
rect 19668 32988 19674 33000
rect 13078 32920 13084 32972
rect 13136 32960 13142 32972
rect 13173 32963 13231 32969
rect 13173 32960 13185 32963
rect 13136 32932 13185 32960
rect 13136 32920 13142 32932
rect 13173 32929 13185 32932
rect 13219 32929 13231 32963
rect 13173 32923 13231 32929
rect 13354 32920 13360 32972
rect 13412 32920 13418 32972
rect 18506 32920 18512 32972
rect 18564 32920 18570 32972
rect 19702 32920 19708 32972
rect 19760 32920 19766 32972
rect 19812 32969 19840 33000
rect 23768 33000 24676 33028
rect 19797 32963 19855 32969
rect 19797 32929 19809 32963
rect 19843 32929 19855 32963
rect 19797 32923 19855 32929
rect 21082 32920 21088 32972
rect 21140 32920 21146 32972
rect 23768 32969 23796 33000
rect 24670 32988 24676 33000
rect 24728 33028 24734 33040
rect 24728 33000 25912 33028
rect 24728 32988 24734 33000
rect 23753 32963 23811 32969
rect 23753 32929 23765 32963
rect 23799 32929 23811 32963
rect 23753 32923 23811 32929
rect 25774 32920 25780 32972
rect 25832 32920 25838 32972
rect 25884 32960 25912 33000
rect 27798 32988 27804 33040
rect 27856 33028 27862 33040
rect 28736 33028 28764 33059
rect 28810 33056 28816 33068
rect 28868 33056 28874 33108
rect 30098 33056 30104 33108
rect 30156 33056 30162 33108
rect 30282 33056 30288 33108
rect 30340 33056 30346 33108
rect 34333 33099 34391 33105
rect 34333 33065 34345 33099
rect 34379 33096 34391 33099
rect 34698 33096 34704 33108
rect 34379 33068 34704 33096
rect 34379 33065 34391 33068
rect 34333 33059 34391 33065
rect 34698 33056 34704 33068
rect 34756 33056 34762 33108
rect 29638 33028 29644 33040
rect 27856 33000 28764 33028
rect 28828 33000 29644 33028
rect 27856 32988 27862 33000
rect 28828 32960 28856 33000
rect 29638 32988 29644 33000
rect 29696 32988 29702 33040
rect 31846 33028 31852 33040
rect 30668 33000 31852 33028
rect 25884 32932 28856 32960
rect 28994 32920 29000 32972
rect 29052 32920 29058 32972
rect 30006 32920 30012 32972
rect 30064 32960 30070 32972
rect 30668 32969 30696 33000
rect 31846 32988 31852 33000
rect 31904 32988 31910 33040
rect 33594 32988 33600 33040
rect 33652 33028 33658 33040
rect 33652 33000 34376 33028
rect 33652 32988 33658 33000
rect 34348 32972 34376 33000
rect 30561 32963 30619 32969
rect 30561 32960 30573 32963
rect 30064 32932 30573 32960
rect 30064 32920 30070 32932
rect 30561 32929 30573 32932
rect 30607 32929 30619 32963
rect 30561 32923 30619 32929
rect 30653 32963 30711 32969
rect 30653 32929 30665 32963
rect 30699 32929 30711 32963
rect 30653 32923 30711 32929
rect 30745 32963 30803 32969
rect 30745 32929 30757 32963
rect 30791 32960 30803 32963
rect 31570 32960 31576 32972
rect 30791 32932 31576 32960
rect 30791 32929 30803 32932
rect 30745 32923 30803 32929
rect 31570 32920 31576 32932
rect 31628 32920 31634 32972
rect 33318 32920 33324 32972
rect 33376 32920 33382 32972
rect 34330 32920 34336 32972
rect 34388 32960 34394 32972
rect 35250 32960 35256 32972
rect 34388 32932 35256 32960
rect 34388 32920 34394 32932
rect 35250 32920 35256 32932
rect 35308 32920 35314 32972
rect 13906 32852 13912 32904
rect 13964 32892 13970 32904
rect 14829 32895 14887 32901
rect 14829 32892 14841 32895
rect 13964 32864 14841 32892
rect 13964 32852 13970 32864
rect 14829 32861 14841 32864
rect 14875 32861 14887 32895
rect 14829 32855 14887 32861
rect 18785 32895 18843 32901
rect 18785 32861 18797 32895
rect 18831 32892 18843 32895
rect 19058 32892 19064 32904
rect 18831 32864 19064 32892
rect 18831 32861 18843 32864
rect 18785 32855 18843 32861
rect 19058 32852 19064 32864
rect 19116 32892 19122 32904
rect 20165 32895 20223 32901
rect 20165 32892 20177 32895
rect 19116 32864 20177 32892
rect 19116 32852 19122 32864
rect 20165 32861 20177 32864
rect 20211 32892 20223 32895
rect 20809 32895 20867 32901
rect 20809 32892 20821 32895
rect 20211 32864 20821 32892
rect 20211 32861 20223 32864
rect 20165 32855 20223 32861
rect 20809 32861 20821 32864
rect 20855 32861 20867 32895
rect 20809 32855 20867 32861
rect 22186 32852 22192 32904
rect 22244 32852 22250 32904
rect 23477 32895 23535 32901
rect 23477 32861 23489 32895
rect 23523 32892 23535 32895
rect 23566 32892 23572 32904
rect 23523 32864 23572 32892
rect 23523 32861 23535 32864
rect 23477 32855 23535 32861
rect 23566 32852 23572 32864
rect 23624 32892 23630 32904
rect 24394 32892 24400 32904
rect 23624 32864 24400 32892
rect 23624 32852 23630 32864
rect 24394 32852 24400 32864
rect 24452 32852 24458 32904
rect 25130 32852 25136 32904
rect 25188 32892 25194 32904
rect 26050 32892 26056 32904
rect 25188 32864 26056 32892
rect 25188 32852 25194 32864
rect 26050 32852 26056 32864
rect 26108 32852 26114 32904
rect 29012 32892 29040 32920
rect 28828 32864 29040 32892
rect 16390 32784 16396 32836
rect 16448 32824 16454 32836
rect 16448 32796 17342 32824
rect 16448 32784 16454 32796
rect 18230 32784 18236 32836
rect 18288 32824 18294 32836
rect 19613 32827 19671 32833
rect 19613 32824 19625 32827
rect 18288 32796 19625 32824
rect 18288 32784 18294 32796
rect 19613 32793 19625 32796
rect 19659 32793 19671 32827
rect 19613 32787 19671 32793
rect 25593 32827 25651 32833
rect 25593 32793 25605 32827
rect 25639 32824 25651 32827
rect 26142 32824 26148 32836
rect 25639 32796 26148 32824
rect 25639 32793 25651 32796
rect 25593 32787 25651 32793
rect 26142 32784 26148 32796
rect 26200 32784 26206 32836
rect 28705 32827 28763 32833
rect 28705 32793 28717 32827
rect 28751 32824 28763 32827
rect 28828 32824 28856 32864
rect 29178 32852 29184 32904
rect 29236 32852 29242 32904
rect 29365 32895 29423 32901
rect 29365 32861 29377 32895
rect 29411 32892 29423 32895
rect 29730 32892 29736 32904
rect 29411 32864 29736 32892
rect 29411 32861 29423 32864
rect 29365 32855 29423 32861
rect 29730 32852 29736 32864
rect 29788 32852 29794 32904
rect 30190 32852 30196 32904
rect 30248 32852 30254 32904
rect 30469 32895 30527 32901
rect 30469 32861 30481 32895
rect 30515 32892 30527 32895
rect 30926 32892 30932 32904
rect 30515 32864 30932 32892
rect 30515 32861 30527 32864
rect 30469 32855 30527 32861
rect 30926 32852 30932 32864
rect 30984 32852 30990 32904
rect 31110 32852 31116 32904
rect 31168 32852 31174 32904
rect 32398 32852 32404 32904
rect 32456 32852 32462 32904
rect 33336 32892 33364 32920
rect 33873 32895 33931 32901
rect 33873 32892 33885 32895
rect 33336 32864 33885 32892
rect 33873 32861 33885 32864
rect 33919 32861 33931 32895
rect 33873 32855 33931 32861
rect 34149 32895 34207 32901
rect 34149 32861 34161 32895
rect 34195 32892 34207 32895
rect 35434 32892 35440 32904
rect 34195 32864 35440 32892
rect 34195 32861 34207 32864
rect 34149 32855 34207 32861
rect 28751 32796 28856 32824
rect 28751 32793 28763 32796
rect 28705 32787 28763 32793
rect 28902 32784 28908 32836
rect 28960 32784 28966 32836
rect 30374 32784 30380 32836
rect 30432 32824 30438 32836
rect 31389 32827 31447 32833
rect 31389 32824 31401 32827
rect 30432 32796 31401 32824
rect 30432 32784 30438 32796
rect 31389 32793 31401 32796
rect 31435 32793 31447 32827
rect 31389 32787 31447 32793
rect 31662 32784 31668 32836
rect 31720 32824 31726 32836
rect 32125 32827 32183 32833
rect 32125 32824 32137 32827
rect 31720 32796 32137 32824
rect 31720 32784 31726 32796
rect 32125 32793 32137 32796
rect 32171 32793 32183 32827
rect 32125 32787 32183 32793
rect 33226 32784 33232 32836
rect 33284 32824 33290 32836
rect 33321 32827 33379 32833
rect 33321 32824 33333 32827
rect 33284 32796 33333 32824
rect 33284 32784 33290 32796
rect 33321 32793 33333 32796
rect 33367 32793 33379 32827
rect 33888 32824 33916 32855
rect 35434 32852 35440 32864
rect 35492 32852 35498 32904
rect 35158 32824 35164 32836
rect 33888 32796 35164 32824
rect 33321 32787 33379 32793
rect 35158 32784 35164 32796
rect 35216 32784 35222 32836
rect 12066 32716 12072 32768
rect 12124 32756 12130 32768
rect 12713 32759 12771 32765
rect 12713 32756 12725 32759
rect 12124 32728 12725 32756
rect 12124 32716 12130 32728
rect 12713 32725 12725 32728
rect 12759 32725 12771 32759
rect 12713 32719 12771 32725
rect 13078 32716 13084 32768
rect 13136 32716 13142 32768
rect 19245 32759 19303 32765
rect 19245 32725 19257 32759
rect 19291 32756 19303 32759
rect 19518 32756 19524 32768
rect 19291 32728 19524 32756
rect 19291 32725 19303 32728
rect 19245 32719 19303 32725
rect 19518 32716 19524 32728
rect 19576 32716 19582 32768
rect 23474 32716 23480 32768
rect 23532 32756 23538 32768
rect 23569 32759 23627 32765
rect 23569 32756 23581 32759
rect 23532 32728 23581 32756
rect 23532 32716 23538 32728
rect 23569 32725 23581 32728
rect 23615 32725 23627 32759
rect 23569 32719 23627 32725
rect 25682 32716 25688 32768
rect 25740 32716 25746 32768
rect 28810 32716 28816 32768
rect 28868 32756 28874 32768
rect 30558 32756 30564 32768
rect 28868 32728 30564 32756
rect 28868 32716 28874 32728
rect 30558 32716 30564 32728
rect 30616 32716 30622 32768
rect 30742 32716 30748 32768
rect 30800 32756 30806 32768
rect 31021 32759 31079 32765
rect 31021 32756 31033 32759
rect 30800 32728 31033 32756
rect 30800 32716 30806 32728
rect 31021 32725 31033 32728
rect 31067 32725 31079 32759
rect 31021 32719 31079 32725
rect 33965 32759 34023 32765
rect 33965 32725 33977 32759
rect 34011 32756 34023 32759
rect 35342 32756 35348 32768
rect 34011 32728 35348 32756
rect 34011 32725 34023 32728
rect 33965 32719 34023 32725
rect 35342 32716 35348 32728
rect 35400 32716 35406 32768
rect 1104 32666 37076 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 37076 32666
rect 1104 32592 37076 32614
rect 18046 32512 18052 32564
rect 18104 32512 18110 32564
rect 22189 32555 22247 32561
rect 22189 32521 22201 32555
rect 22235 32552 22247 32555
rect 22278 32552 22284 32564
rect 22235 32524 22284 32552
rect 22235 32521 22247 32524
rect 22189 32515 22247 32521
rect 22278 32512 22284 32524
rect 22336 32512 22342 32564
rect 25774 32512 25780 32564
rect 25832 32552 25838 32564
rect 28905 32555 28963 32561
rect 25832 32524 28764 32552
rect 25832 32512 25838 32524
rect 14829 32487 14887 32493
rect 14829 32453 14841 32487
rect 14875 32484 14887 32487
rect 15562 32484 15568 32496
rect 14875 32456 15568 32484
rect 14875 32453 14887 32456
rect 14829 32447 14887 32453
rect 15562 32444 15568 32456
rect 15620 32444 15626 32496
rect 16390 32444 16396 32496
rect 16448 32484 16454 32496
rect 16448 32456 18354 32484
rect 16448 32444 16454 32456
rect 19518 32444 19524 32496
rect 19576 32444 19582 32496
rect 20346 32444 20352 32496
rect 20404 32484 20410 32496
rect 24854 32484 24860 32496
rect 20404 32456 24860 32484
rect 20404 32444 20410 32456
rect 24854 32444 24860 32456
rect 24912 32484 24918 32496
rect 25869 32487 25927 32493
rect 25869 32484 25881 32487
rect 24912 32456 25881 32484
rect 24912 32444 24918 32456
rect 25869 32453 25881 32456
rect 25915 32484 25927 32487
rect 27706 32484 27712 32496
rect 25915 32456 27712 32484
rect 25915 32453 25927 32456
rect 25869 32447 25927 32453
rect 27706 32444 27712 32456
rect 27764 32444 27770 32496
rect 27890 32444 27896 32496
rect 27948 32444 27954 32496
rect 28736 32484 28764 32524
rect 28905 32521 28917 32555
rect 28951 32552 28963 32555
rect 28994 32552 29000 32564
rect 28951 32524 29000 32552
rect 28951 32521 28963 32524
rect 28905 32515 28963 32521
rect 28994 32512 29000 32524
rect 29052 32512 29058 32564
rect 31294 32552 31300 32564
rect 29104 32524 30328 32552
rect 29104 32484 29132 32524
rect 28736 32456 29132 32484
rect 29178 32444 29184 32496
rect 29236 32484 29242 32496
rect 30161 32487 30219 32493
rect 30161 32484 30173 32487
rect 29236 32456 30173 32484
rect 29236 32444 29242 32456
rect 30161 32453 30173 32456
rect 30207 32453 30219 32487
rect 30161 32447 30219 32453
rect 14274 32376 14280 32428
rect 14332 32416 14338 32428
rect 16408 32416 16436 32444
rect 14332 32388 16436 32416
rect 14332 32376 14338 32388
rect 17034 32376 17040 32428
rect 17092 32376 17098 32428
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32416 25835 32419
rect 26050 32416 26056 32428
rect 25823 32388 26056 32416
rect 25823 32385 25835 32388
rect 25777 32379 25835 32385
rect 26050 32376 26056 32388
rect 26108 32416 26114 32428
rect 26605 32419 26663 32425
rect 26605 32416 26617 32419
rect 26108 32388 26617 32416
rect 26108 32376 26114 32388
rect 26605 32385 26617 32388
rect 26651 32416 26663 32419
rect 27157 32419 27215 32425
rect 27157 32416 27169 32419
rect 26651 32388 27169 32416
rect 26651 32385 26663 32388
rect 26605 32379 26663 32385
rect 27157 32385 27169 32388
rect 27203 32385 27215 32419
rect 27157 32379 27215 32385
rect 29733 32419 29791 32425
rect 29733 32385 29745 32419
rect 29779 32385 29791 32419
rect 29733 32379 29791 32385
rect 11606 32308 11612 32360
rect 11664 32348 11670 32360
rect 12897 32351 12955 32357
rect 12897 32348 12909 32351
rect 11664 32320 12909 32348
rect 11664 32308 11670 32320
rect 12897 32317 12909 32320
rect 12943 32317 12955 32351
rect 12897 32311 12955 32317
rect 12912 32212 12940 32311
rect 13170 32308 13176 32360
rect 13228 32308 13234 32360
rect 15286 32308 15292 32360
rect 15344 32348 15350 32360
rect 15565 32351 15623 32357
rect 15565 32348 15577 32351
rect 15344 32320 15577 32348
rect 15344 32308 15350 32320
rect 15565 32317 15577 32320
rect 15611 32317 15623 32351
rect 15565 32311 15623 32317
rect 15930 32308 15936 32360
rect 15988 32348 15994 32360
rect 17129 32351 17187 32357
rect 17129 32348 17141 32351
rect 15988 32320 17141 32348
rect 15988 32308 15994 32320
rect 17129 32317 17141 32320
rect 17175 32317 17187 32351
rect 17129 32311 17187 32317
rect 17313 32351 17371 32357
rect 17313 32317 17325 32351
rect 17359 32348 17371 32351
rect 17402 32348 17408 32360
rect 17359 32320 17408 32348
rect 17359 32317 17371 32320
rect 17313 32311 17371 32317
rect 17402 32308 17408 32320
rect 17460 32308 17466 32360
rect 19797 32351 19855 32357
rect 19797 32317 19809 32351
rect 19843 32348 19855 32351
rect 21085 32351 21143 32357
rect 21085 32348 21097 32351
rect 19843 32320 21097 32348
rect 19843 32317 19855 32320
rect 19797 32311 19855 32317
rect 21085 32317 21097 32320
rect 21131 32317 21143 32351
rect 21085 32311 21143 32317
rect 13906 32212 13912 32224
rect 12912 32184 13912 32212
rect 13906 32172 13912 32184
rect 13964 32212 13970 32224
rect 14182 32212 14188 32224
rect 13964 32184 14188 32212
rect 13964 32172 13970 32184
rect 14182 32172 14188 32184
rect 14240 32172 14246 32224
rect 14645 32215 14703 32221
rect 14645 32181 14657 32215
rect 14691 32212 14703 32215
rect 14826 32212 14832 32224
rect 14691 32184 14832 32212
rect 14691 32181 14703 32184
rect 14645 32175 14703 32181
rect 14826 32172 14832 32184
rect 14884 32172 14890 32224
rect 15562 32172 15568 32224
rect 15620 32212 15626 32224
rect 16669 32215 16727 32221
rect 16669 32212 16681 32215
rect 15620 32184 16681 32212
rect 15620 32172 15626 32184
rect 16669 32181 16681 32184
rect 16715 32181 16727 32215
rect 16669 32175 16727 32181
rect 19058 32172 19064 32224
rect 19116 32212 19122 32224
rect 19812 32212 19840 32311
rect 22094 32308 22100 32360
rect 22152 32348 22158 32360
rect 22281 32351 22339 32357
rect 22281 32348 22293 32351
rect 22152 32320 22293 32348
rect 22152 32308 22158 32320
rect 22281 32317 22293 32320
rect 22327 32317 22339 32351
rect 22281 32311 22339 32317
rect 22462 32308 22468 32360
rect 22520 32308 22526 32360
rect 27433 32351 27491 32357
rect 27433 32317 27445 32351
rect 27479 32348 27491 32351
rect 28074 32348 28080 32360
rect 27479 32320 28080 32348
rect 27479 32317 27491 32320
rect 27433 32311 27491 32317
rect 28074 32308 28080 32320
rect 28132 32308 28138 32360
rect 29748 32348 29776 32379
rect 29914 32376 29920 32428
rect 29972 32376 29978 32428
rect 30300 32416 30328 32524
rect 30392 32524 31300 32552
rect 30392 32493 30420 32524
rect 31294 32512 31300 32524
rect 31352 32512 31358 32564
rect 32858 32552 32864 32564
rect 31726 32524 32864 32552
rect 30377 32487 30435 32493
rect 30377 32453 30389 32487
rect 30423 32453 30435 32487
rect 30377 32447 30435 32453
rect 31113 32487 31171 32493
rect 31113 32453 31125 32487
rect 31159 32484 31171 32487
rect 31386 32484 31392 32496
rect 31159 32456 31392 32484
rect 31159 32453 31171 32456
rect 31113 32447 31171 32453
rect 31386 32444 31392 32456
rect 31444 32444 31450 32496
rect 31726 32484 31754 32524
rect 32858 32512 32864 32524
rect 32916 32512 32922 32564
rect 35253 32555 35311 32561
rect 35253 32552 35265 32555
rect 32968 32524 35265 32552
rect 31496 32456 31754 32484
rect 30300 32388 30696 32416
rect 29822 32348 29828 32360
rect 29748 32320 29828 32348
rect 29822 32308 29828 32320
rect 29880 32348 29886 32360
rect 30469 32351 30527 32357
rect 29880 32320 29960 32348
rect 29880 32308 29886 32320
rect 29932 32280 29960 32320
rect 30469 32317 30481 32351
rect 30515 32348 30527 32351
rect 30558 32348 30564 32360
rect 30515 32320 30564 32348
rect 30515 32317 30527 32320
rect 30469 32311 30527 32317
rect 30558 32308 30564 32320
rect 30616 32308 30622 32360
rect 30668 32348 30696 32388
rect 30742 32376 30748 32428
rect 30800 32376 30806 32428
rect 31496 32348 31524 32456
rect 31662 32376 31668 32428
rect 31720 32416 31726 32428
rect 31849 32419 31907 32425
rect 31849 32416 31861 32419
rect 31720 32388 31861 32416
rect 31720 32376 31726 32388
rect 31849 32385 31861 32388
rect 31895 32416 31907 32419
rect 31895 32388 32536 32416
rect 31895 32385 31907 32388
rect 31849 32379 31907 32385
rect 30668 32320 31524 32348
rect 32508 32348 32536 32388
rect 32582 32376 32588 32428
rect 32640 32376 32646 32428
rect 32968 32425 32996 32524
rect 35253 32521 35265 32524
rect 35299 32521 35311 32555
rect 35253 32515 35311 32521
rect 33962 32444 33968 32496
rect 34020 32444 34026 32496
rect 32953 32419 33011 32425
rect 32953 32385 32965 32419
rect 32999 32385 33011 32419
rect 32953 32379 33011 32385
rect 34422 32376 34428 32428
rect 34480 32376 34486 32428
rect 34977 32419 35035 32425
rect 34977 32385 34989 32419
rect 35023 32385 35035 32419
rect 34977 32379 35035 32385
rect 33137 32351 33195 32357
rect 33137 32348 33149 32351
rect 32508 32320 33149 32348
rect 33137 32317 33149 32320
rect 33183 32348 33195 32351
rect 33413 32351 33471 32357
rect 33183 32320 33272 32348
rect 33183 32317 33195 32320
rect 33137 32311 33195 32317
rect 30653 32283 30711 32289
rect 30653 32280 30665 32283
rect 29932 32252 30665 32280
rect 30653 32249 30665 32252
rect 30699 32249 30711 32283
rect 30653 32243 30711 32249
rect 31297 32283 31355 32289
rect 31297 32249 31309 32283
rect 31343 32280 31355 32283
rect 32306 32280 32312 32292
rect 31343 32252 32312 32280
rect 31343 32249 31355 32252
rect 31297 32243 31355 32249
rect 32306 32240 32312 32252
rect 32364 32240 32370 32292
rect 19116 32184 19840 32212
rect 19116 32172 19122 32184
rect 20990 32172 20996 32224
rect 21048 32212 21054 32224
rect 21821 32215 21879 32221
rect 21821 32212 21833 32215
rect 21048 32184 21833 32212
rect 21048 32172 21054 32184
rect 21821 32181 21833 32184
rect 21867 32181 21879 32215
rect 21821 32175 21879 32181
rect 29914 32172 29920 32224
rect 29972 32172 29978 32224
rect 30009 32215 30067 32221
rect 30009 32181 30021 32215
rect 30055 32212 30067 32215
rect 30098 32212 30104 32224
rect 30055 32184 30104 32212
rect 30055 32181 30067 32184
rect 30009 32175 30067 32181
rect 30098 32172 30104 32184
rect 30156 32172 30162 32224
rect 30193 32215 30251 32221
rect 30193 32181 30205 32215
rect 30239 32212 30251 32215
rect 30282 32212 30288 32224
rect 30239 32184 30288 32212
rect 30239 32181 30251 32184
rect 30193 32175 30251 32181
rect 30282 32172 30288 32184
rect 30340 32172 30346 32224
rect 30374 32172 30380 32224
rect 30432 32212 30438 32224
rect 30561 32215 30619 32221
rect 30561 32212 30573 32215
rect 30432 32184 30573 32212
rect 30432 32172 30438 32184
rect 30561 32181 30573 32184
rect 30607 32181 30619 32215
rect 33244 32212 33272 32320
rect 33413 32317 33425 32351
rect 33459 32348 33471 32351
rect 34440 32348 34468 32376
rect 33459 32320 34468 32348
rect 33459 32317 33471 32320
rect 33413 32311 33471 32317
rect 34606 32308 34612 32360
rect 34664 32348 34670 32360
rect 34992 32348 35020 32379
rect 35158 32376 35164 32428
rect 35216 32376 35222 32428
rect 35250 32376 35256 32428
rect 35308 32416 35314 32428
rect 35437 32419 35495 32425
rect 35437 32416 35449 32419
rect 35308 32388 35449 32416
rect 35308 32376 35314 32388
rect 35437 32385 35449 32388
rect 35483 32385 35495 32419
rect 35437 32379 35495 32385
rect 34664 32320 35020 32348
rect 34664 32308 34670 32320
rect 34514 32240 34520 32292
rect 34572 32280 34578 32292
rect 35069 32283 35127 32289
rect 35069 32280 35081 32283
rect 34572 32252 35081 32280
rect 34572 32240 34578 32252
rect 35069 32249 35081 32252
rect 35115 32249 35127 32283
rect 35069 32243 35127 32249
rect 34146 32212 34152 32224
rect 33244 32184 34152 32212
rect 30561 32175 30619 32181
rect 34146 32172 34152 32184
rect 34204 32172 34210 32224
rect 34885 32215 34943 32221
rect 34885 32181 34897 32215
rect 34931 32212 34943 32215
rect 35342 32212 35348 32224
rect 34931 32184 35348 32212
rect 34931 32181 34943 32184
rect 34885 32175 34943 32181
rect 35342 32172 35348 32184
rect 35400 32172 35406 32224
rect 1104 32122 37076 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 37076 32122
rect 1104 32048 37076 32070
rect 13078 31968 13084 32020
rect 13136 32008 13142 32020
rect 13538 32008 13544 32020
rect 13136 31980 13544 32008
rect 13136 31968 13142 31980
rect 13538 31968 13544 31980
rect 13596 31968 13602 32020
rect 17034 31968 17040 32020
rect 17092 31968 17098 32020
rect 22278 31968 22284 32020
rect 22336 32008 22342 32020
rect 22465 32011 22523 32017
rect 22465 32008 22477 32011
rect 22336 31980 22477 32008
rect 22336 31968 22342 31980
rect 22465 31977 22477 31980
rect 22511 31977 22523 32011
rect 22465 31971 22523 31977
rect 26050 31968 26056 32020
rect 26108 32008 26114 32020
rect 26108 31980 27568 32008
rect 26108 31968 26114 31980
rect 13814 31900 13820 31952
rect 13872 31940 13878 31952
rect 27433 31943 27491 31949
rect 27433 31940 27445 31943
rect 13872 31912 15056 31940
rect 13872 31900 13878 31912
rect 12066 31832 12072 31884
rect 12124 31832 12130 31884
rect 14274 31872 14280 31884
rect 13188 31844 14280 31872
rect 11606 31764 11612 31816
rect 11664 31804 11670 31816
rect 11793 31807 11851 31813
rect 11793 31804 11805 31807
rect 11664 31776 11805 31804
rect 11664 31764 11670 31776
rect 11793 31773 11805 31776
rect 11839 31773 11851 31807
rect 13188 31790 13216 31844
rect 14274 31832 14280 31844
rect 14332 31832 14338 31884
rect 14826 31832 14832 31884
rect 14884 31872 14890 31884
rect 15028 31881 15056 31912
rect 27264 31912 27445 31940
rect 14921 31875 14979 31881
rect 14921 31872 14933 31875
rect 14884 31844 14933 31872
rect 14884 31832 14890 31844
rect 14921 31841 14933 31844
rect 14967 31841 14979 31875
rect 14921 31835 14979 31841
rect 15013 31875 15071 31881
rect 15013 31841 15025 31875
rect 15059 31841 15071 31875
rect 15013 31835 15071 31841
rect 15562 31832 15568 31884
rect 15620 31832 15626 31884
rect 19058 31832 19064 31884
rect 19116 31872 19122 31884
rect 20717 31875 20775 31881
rect 20717 31872 20729 31875
rect 19116 31844 20729 31872
rect 19116 31832 19122 31844
rect 20717 31841 20729 31844
rect 20763 31841 20775 31875
rect 20717 31835 20775 31841
rect 20990 31832 20996 31884
rect 21048 31832 21054 31884
rect 22186 31832 22192 31884
rect 22244 31832 22250 31884
rect 23566 31832 23572 31884
rect 23624 31832 23630 31884
rect 23753 31875 23811 31881
rect 23753 31841 23765 31875
rect 23799 31872 23811 31875
rect 24762 31872 24768 31884
rect 23799 31844 24768 31872
rect 23799 31841 23811 31844
rect 23753 31835 23811 31841
rect 24762 31832 24768 31844
rect 24820 31872 24826 31884
rect 24949 31875 25007 31881
rect 24949 31872 24961 31875
rect 24820 31844 24961 31872
rect 24820 31832 24826 31844
rect 24949 31841 24961 31844
rect 24995 31841 25007 31875
rect 24949 31835 25007 31841
rect 25593 31875 25651 31881
rect 25593 31841 25605 31875
rect 25639 31872 25651 31875
rect 25682 31872 25688 31884
rect 25639 31844 25688 31872
rect 25639 31841 25651 31844
rect 25593 31835 25651 31841
rect 25682 31832 25688 31844
rect 25740 31872 25746 31884
rect 26970 31872 26976 31884
rect 25740 31844 26976 31872
rect 25740 31832 25746 31844
rect 26970 31832 26976 31844
rect 27028 31832 27034 31884
rect 27065 31875 27123 31881
rect 27065 31841 27077 31875
rect 27111 31872 27123 31875
rect 27264 31872 27292 31912
rect 27433 31909 27445 31912
rect 27479 31909 27491 31943
rect 27433 31903 27491 31909
rect 27111 31844 27292 31872
rect 27341 31875 27399 31881
rect 27111 31841 27123 31844
rect 27065 31835 27123 31841
rect 27341 31841 27353 31875
rect 27387 31872 27399 31875
rect 27540 31872 27568 31980
rect 27614 31968 27620 32020
rect 27672 32008 27678 32020
rect 30282 32008 30288 32020
rect 27672 31980 30288 32008
rect 27672 31968 27678 31980
rect 27387 31844 27568 31872
rect 27387 31841 27399 31844
rect 27341 31835 27399 31841
rect 27982 31832 27988 31884
rect 28040 31832 28046 31884
rect 11793 31767 11851 31773
rect 14182 31764 14188 31816
rect 14240 31804 14246 31816
rect 15286 31804 15292 31816
rect 14240 31776 15292 31804
rect 14240 31764 14246 31776
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 22204 31804 22232 31832
rect 22126 31776 22232 31804
rect 25222 31764 25228 31816
rect 25280 31804 25286 31816
rect 28905 31807 28963 31813
rect 25280 31776 25990 31804
rect 25280 31764 25286 31776
rect 28905 31773 28917 31807
rect 28951 31804 28963 31807
rect 29104 31804 29132 31980
rect 30282 31968 30288 31980
rect 30340 31968 30346 32020
rect 32582 31968 32588 32020
rect 32640 32008 32646 32020
rect 32640 31980 34744 32008
rect 32640 31968 32646 31980
rect 29914 31900 29920 31952
rect 29972 31900 29978 31952
rect 34333 31943 34391 31949
rect 34333 31909 34345 31943
rect 34379 31940 34391 31943
rect 34606 31940 34612 31952
rect 34379 31912 34612 31940
rect 34379 31909 34391 31912
rect 34333 31903 34391 31909
rect 34606 31900 34612 31912
rect 34664 31900 34670 31952
rect 29932 31872 29960 31900
rect 30745 31875 30803 31881
rect 30745 31872 30757 31875
rect 29932 31844 30757 31872
rect 30745 31841 30757 31844
rect 30791 31841 30803 31875
rect 30745 31835 30803 31841
rect 31386 31832 31392 31884
rect 31444 31872 31450 31884
rect 32585 31875 32643 31881
rect 31444 31844 32536 31872
rect 31444 31832 31450 31844
rect 28951 31776 29132 31804
rect 28951 31773 28963 31776
rect 28905 31767 28963 31773
rect 29178 31764 29184 31816
rect 29236 31764 29242 31816
rect 29365 31807 29423 31813
rect 29365 31773 29377 31807
rect 29411 31804 29423 31807
rect 29822 31804 29828 31816
rect 29411 31776 29828 31804
rect 29411 31773 29423 31776
rect 29365 31767 29423 31773
rect 29822 31764 29828 31776
rect 29880 31804 29886 31816
rect 29917 31807 29975 31813
rect 29917 31804 29929 31807
rect 29880 31776 29929 31804
rect 29880 31764 29886 31776
rect 29917 31773 29929 31776
rect 29963 31773 29975 31807
rect 29917 31767 29975 31773
rect 30098 31764 30104 31816
rect 30156 31764 30162 31816
rect 30466 31764 30472 31816
rect 30524 31764 30530 31816
rect 32508 31813 32536 31844
rect 32585 31841 32597 31875
rect 32631 31872 32643 31875
rect 34146 31872 34152 31884
rect 32631 31844 34152 31872
rect 32631 31841 32643 31844
rect 32585 31835 32643 31841
rect 34146 31832 34152 31844
rect 34204 31832 34210 31884
rect 32493 31807 32551 31813
rect 32493 31804 32505 31807
rect 32451 31776 32505 31804
rect 32493 31773 32505 31776
rect 32539 31804 32551 31807
rect 32539 31776 32628 31804
rect 32539 31773 32551 31776
rect 32493 31767 32551 31773
rect 18874 31736 18880 31748
rect 16790 31708 18880 31736
rect 14458 31628 14464 31680
rect 14516 31628 14522 31680
rect 14829 31671 14887 31677
rect 14829 31637 14841 31671
rect 14875 31668 14887 31671
rect 15930 31668 15936 31680
rect 14875 31640 15936 31668
rect 14875 31637 14887 31640
rect 14829 31631 14887 31637
rect 15930 31628 15936 31640
rect 15988 31628 15994 31680
rect 16298 31628 16304 31680
rect 16356 31668 16362 31680
rect 16868 31668 16896 31708
rect 18874 31696 18880 31708
rect 18932 31696 18938 31748
rect 23477 31739 23535 31745
rect 23477 31705 23489 31739
rect 23523 31736 23535 31739
rect 24765 31739 24823 31745
rect 23523 31708 24532 31736
rect 23523 31705 23535 31708
rect 23477 31699 23535 31705
rect 24504 31680 24532 31708
rect 24765 31705 24777 31739
rect 24811 31736 24823 31739
rect 25774 31736 25780 31748
rect 24811 31708 25780 31736
rect 24811 31705 24823 31708
rect 24765 31699 24823 31705
rect 25774 31696 25780 31708
rect 25832 31696 25838 31748
rect 26970 31696 26976 31748
rect 27028 31736 27034 31748
rect 27801 31739 27859 31745
rect 27801 31736 27813 31739
rect 27028 31708 27813 31736
rect 27028 31696 27034 31708
rect 27801 31705 27813 31708
rect 27847 31705 27859 31739
rect 27801 31699 27859 31705
rect 30650 31696 30656 31748
rect 30708 31736 30714 31748
rect 30708 31708 31234 31736
rect 30708 31696 30714 31708
rect 16356 31640 16896 31668
rect 16356 31628 16362 31640
rect 22554 31628 22560 31680
rect 22612 31668 22618 31680
rect 23109 31671 23167 31677
rect 23109 31668 23121 31671
rect 22612 31640 23121 31668
rect 22612 31628 22618 31640
rect 23109 31637 23121 31640
rect 23155 31637 23167 31671
rect 23109 31631 23167 31637
rect 24394 31628 24400 31680
rect 24452 31628 24458 31680
rect 24486 31628 24492 31680
rect 24544 31668 24550 31680
rect 24857 31671 24915 31677
rect 24857 31668 24869 31671
rect 24544 31640 24869 31668
rect 24544 31628 24550 31640
rect 24857 31637 24869 31640
rect 24903 31637 24915 31671
rect 24857 31631 24915 31637
rect 27890 31628 27896 31680
rect 27948 31628 27954 31680
rect 29825 31671 29883 31677
rect 29825 31637 29837 31671
rect 29871 31668 29883 31671
rect 30282 31668 30288 31680
rect 29871 31640 30288 31668
rect 29871 31637 29883 31640
rect 29825 31631 29883 31637
rect 30282 31628 30288 31640
rect 30340 31628 30346 31680
rect 32600 31668 32628 31776
rect 33962 31764 33968 31816
rect 34020 31764 34026 31816
rect 34716 31813 34744 31980
rect 35434 31832 35440 31884
rect 35492 31832 35498 31884
rect 34701 31807 34759 31813
rect 34701 31773 34713 31807
rect 34747 31773 34759 31807
rect 34701 31767 34759 31773
rect 32858 31696 32864 31748
rect 32916 31696 32922 31748
rect 33594 31668 33600 31680
rect 32600 31640 33600 31668
rect 33594 31628 33600 31640
rect 33652 31628 33658 31680
rect 1104 31578 37076 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 37076 31578
rect 1104 31504 37076 31526
rect 13170 31424 13176 31476
rect 13228 31464 13234 31476
rect 13357 31467 13415 31473
rect 13357 31464 13369 31467
rect 13228 31436 13369 31464
rect 13228 31424 13234 31436
rect 13357 31433 13369 31436
rect 13403 31433 13415 31467
rect 13357 31427 13415 31433
rect 13538 31424 13544 31476
rect 13596 31464 13602 31476
rect 13817 31467 13875 31473
rect 13817 31464 13829 31467
rect 13596 31436 13829 31464
rect 13596 31424 13602 31436
rect 13817 31433 13829 31436
rect 13863 31433 13875 31467
rect 14826 31464 14832 31476
rect 13817 31427 13875 31433
rect 14292 31436 14832 31464
rect 9398 31356 9404 31408
rect 9456 31356 9462 31408
rect 13725 31399 13783 31405
rect 13725 31365 13737 31399
rect 13771 31396 13783 31399
rect 14292 31396 14320 31436
rect 14826 31424 14832 31436
rect 14884 31424 14890 31476
rect 15930 31424 15936 31476
rect 15988 31424 15994 31476
rect 17034 31424 17040 31476
rect 17092 31464 17098 31476
rect 17221 31467 17279 31473
rect 17221 31464 17233 31467
rect 17092 31436 17233 31464
rect 17092 31424 17098 31436
rect 17221 31433 17233 31436
rect 17267 31433 17279 31467
rect 19058 31464 19064 31476
rect 17221 31427 17279 31433
rect 18432 31436 19064 31464
rect 13771 31368 14320 31396
rect 13771 31365 13783 31368
rect 13725 31359 13783 31365
rect 14458 31356 14464 31408
rect 14516 31356 14522 31408
rect 16298 31396 16304 31408
rect 15686 31368 16304 31396
rect 16298 31356 16304 31368
rect 16356 31356 16362 31408
rect 18432 31396 18460 31436
rect 19058 31424 19064 31436
rect 19116 31424 19122 31476
rect 21637 31467 21695 31473
rect 21637 31433 21649 31467
rect 21683 31464 21695 31467
rect 22094 31464 22100 31476
rect 21683 31436 22100 31464
rect 21683 31433 21695 31436
rect 21637 31427 21695 31433
rect 22094 31424 22100 31436
rect 22152 31424 22158 31476
rect 23937 31467 23995 31473
rect 22204 31436 22876 31464
rect 22204 31408 22232 31436
rect 18064 31368 18460 31396
rect 9953 31331 10011 31337
rect 9953 31328 9965 31331
rect 9876 31300 9965 31328
rect 8110 31220 8116 31272
rect 8168 31220 8174 31272
rect 8389 31263 8447 31269
rect 8389 31229 8401 31263
rect 8435 31260 8447 31263
rect 8938 31260 8944 31272
rect 8435 31232 8944 31260
rect 8435 31229 8447 31232
rect 8389 31223 8447 31229
rect 8938 31220 8944 31232
rect 8996 31220 9002 31272
rect 9674 31084 9680 31136
rect 9732 31124 9738 31136
rect 9876 31133 9904 31300
rect 9953 31297 9965 31300
rect 9999 31297 10011 31331
rect 9953 31291 10011 31297
rect 14182 31288 14188 31340
rect 14240 31288 14246 31340
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31328 17187 31331
rect 17954 31328 17960 31340
rect 17175 31300 17960 31328
rect 17175 31297 17187 31300
rect 17129 31291 17187 31297
rect 17954 31288 17960 31300
rect 18012 31288 18018 31340
rect 18064 31337 18092 31368
rect 18874 31356 18880 31408
rect 18932 31356 18938 31408
rect 22186 31396 22192 31408
rect 21390 31368 22192 31396
rect 22186 31356 22192 31368
rect 22244 31356 22250 31408
rect 22465 31399 22523 31405
rect 22465 31365 22477 31399
rect 22511 31396 22523 31399
rect 22554 31396 22560 31408
rect 22511 31368 22560 31396
rect 22511 31365 22523 31368
rect 22465 31359 22523 31365
rect 22554 31356 22560 31368
rect 22612 31356 22618 31408
rect 22848 31396 22876 31436
rect 23937 31433 23949 31467
rect 23983 31464 23995 31467
rect 24486 31464 24492 31476
rect 23983 31436 24492 31464
rect 23983 31433 23995 31436
rect 23937 31427 23995 31433
rect 24486 31424 24492 31436
rect 24544 31424 24550 31476
rect 25774 31424 25780 31476
rect 25832 31464 25838 31476
rect 26329 31467 26387 31473
rect 26329 31464 26341 31467
rect 25832 31436 26341 31464
rect 25832 31424 25838 31436
rect 26329 31433 26341 31436
rect 26375 31433 26387 31467
rect 26329 31427 26387 31433
rect 28813 31467 28871 31473
rect 28813 31433 28825 31467
rect 28859 31464 28871 31467
rect 28994 31464 29000 31476
rect 28859 31436 29000 31464
rect 28859 31433 28871 31436
rect 28813 31427 28871 31433
rect 28994 31424 29000 31436
rect 29052 31424 29058 31476
rect 31849 31467 31907 31473
rect 31849 31433 31861 31467
rect 31895 31464 31907 31467
rect 32858 31464 32864 31476
rect 31895 31436 32864 31464
rect 31895 31433 31907 31436
rect 31849 31427 31907 31433
rect 32858 31424 32864 31436
rect 32916 31424 32922 31476
rect 24305 31399 24363 31405
rect 22848 31368 22954 31396
rect 24305 31365 24317 31399
rect 24351 31396 24363 31399
rect 24394 31396 24400 31408
rect 24351 31368 24400 31396
rect 24351 31365 24363 31368
rect 24305 31359 24363 31365
rect 24394 31356 24400 31368
rect 24452 31356 24458 31408
rect 25314 31356 25320 31408
rect 25372 31356 25378 31408
rect 27522 31356 27528 31408
rect 27580 31396 27586 31408
rect 27706 31396 27712 31408
rect 27580 31368 27712 31396
rect 27580 31356 27586 31368
rect 27706 31356 27712 31368
rect 27764 31356 27770 31408
rect 30282 31356 30288 31408
rect 30340 31356 30346 31408
rect 33873 31399 33931 31405
rect 33873 31396 33885 31399
rect 31956 31368 33885 31396
rect 18049 31331 18107 31337
rect 18049 31297 18061 31331
rect 18095 31297 18107 31331
rect 18049 31291 18107 31297
rect 26237 31331 26295 31337
rect 26237 31297 26249 31331
rect 26283 31328 26295 31331
rect 26326 31328 26332 31340
rect 26283 31300 26332 31328
rect 26283 31297 26295 31300
rect 26237 31291 26295 31297
rect 26326 31288 26332 31300
rect 26384 31288 26390 31340
rect 13814 31220 13820 31272
rect 13872 31260 13878 31272
rect 13909 31263 13967 31269
rect 13909 31260 13921 31263
rect 13872 31232 13921 31260
rect 13872 31220 13878 31232
rect 13909 31229 13921 31232
rect 13955 31229 13967 31263
rect 13909 31223 13967 31229
rect 17402 31220 17408 31272
rect 17460 31220 17466 31272
rect 18322 31220 18328 31272
rect 18380 31220 18386 31272
rect 19058 31220 19064 31272
rect 19116 31260 19122 31272
rect 19889 31263 19947 31269
rect 19889 31260 19901 31263
rect 19116 31232 19901 31260
rect 19116 31220 19122 31232
rect 19889 31229 19901 31232
rect 19935 31229 19947 31263
rect 19889 31223 19947 31229
rect 16390 31152 16396 31204
rect 16448 31192 16454 31204
rect 17420 31192 17448 31220
rect 16448 31164 17448 31192
rect 16448 31152 16454 31164
rect 9861 31127 9919 31133
rect 9861 31124 9873 31127
rect 9732 31096 9873 31124
rect 9732 31084 9738 31096
rect 9861 31093 9873 31096
rect 9907 31093 9919 31127
rect 9861 31087 9919 31093
rect 9950 31084 9956 31136
rect 10008 31124 10014 31136
rect 10045 31127 10103 31133
rect 10045 31124 10057 31127
rect 10008 31096 10057 31124
rect 10008 31084 10014 31096
rect 10045 31093 10057 31096
rect 10091 31093 10103 31127
rect 10045 31087 10103 31093
rect 16022 31084 16028 31136
rect 16080 31124 16086 31136
rect 16761 31127 16819 31133
rect 16761 31124 16773 31127
rect 16080 31096 16773 31124
rect 16080 31084 16086 31096
rect 16761 31093 16773 31096
rect 16807 31093 16819 31127
rect 17420 31124 17448 31164
rect 19334 31124 19340 31136
rect 17420 31096 19340 31124
rect 16761 31087 16819 31093
rect 19334 31084 19340 31096
rect 19392 31084 19398 31136
rect 19610 31084 19616 31136
rect 19668 31124 19674 31136
rect 19797 31127 19855 31133
rect 19797 31124 19809 31127
rect 19668 31096 19809 31124
rect 19668 31084 19674 31096
rect 19797 31093 19809 31096
rect 19843 31093 19855 31127
rect 19904 31124 19932 31223
rect 20162 31220 20168 31272
rect 20220 31220 20226 31272
rect 22189 31263 22247 31269
rect 22189 31260 22201 31263
rect 21192 31232 22201 31260
rect 21192 31124 21220 31232
rect 22189 31229 22201 31232
rect 22235 31229 22247 31263
rect 22189 31223 22247 31229
rect 24029 31263 24087 31269
rect 24029 31229 24041 31263
rect 24075 31260 24087 31263
rect 24394 31260 24400 31272
rect 24075 31232 24400 31260
rect 24075 31229 24087 31232
rect 24029 31223 24087 31229
rect 24394 31220 24400 31232
rect 24452 31260 24458 31272
rect 25774 31260 25780 31272
rect 24452 31232 25780 31260
rect 24452 31220 24458 31232
rect 25774 31220 25780 31232
rect 25832 31260 25838 31272
rect 26050 31260 26056 31272
rect 25832 31232 26056 31260
rect 25832 31220 25838 31232
rect 26050 31220 26056 31232
rect 26108 31260 26114 31272
rect 26108 31232 26234 31260
rect 26108 31220 26114 31232
rect 26206 31192 26234 31232
rect 26510 31220 26516 31272
rect 26568 31220 26574 31272
rect 26973 31263 27031 31269
rect 26973 31229 26985 31263
rect 27019 31229 27031 31263
rect 26973 31223 27031 31229
rect 26988 31192 27016 31223
rect 27246 31220 27252 31272
rect 27304 31220 27310 31272
rect 28902 31220 28908 31272
rect 28960 31260 28966 31272
rect 29196 31260 29224 31314
rect 30558 31288 30564 31340
rect 30616 31328 30622 31340
rect 31662 31328 31668 31340
rect 30616 31300 31668 31328
rect 30616 31288 30622 31300
rect 31662 31288 31668 31300
rect 31720 31288 31726 31340
rect 31956 31337 31984 31368
rect 33873 31365 33885 31368
rect 33919 31365 33931 31399
rect 34790 31396 34796 31408
rect 33873 31359 33931 31365
rect 34348 31368 34796 31396
rect 31941 31331 31999 31337
rect 31941 31297 31953 31331
rect 31987 31297 31999 31331
rect 31941 31291 31999 31297
rect 32306 31288 32312 31340
rect 32364 31328 32370 31340
rect 34348 31337 34376 31368
rect 34790 31356 34796 31368
rect 34848 31356 34854 31408
rect 32401 31331 32459 31337
rect 32401 31328 32413 31331
rect 32364 31300 32413 31328
rect 32364 31288 32370 31300
rect 32401 31297 32413 31300
rect 32447 31297 32459 31331
rect 32401 31291 32459 31297
rect 34333 31331 34391 31337
rect 34333 31297 34345 31331
rect 34379 31297 34391 31331
rect 34333 31291 34391 31297
rect 34514 31288 34520 31340
rect 34572 31288 34578 31340
rect 34606 31288 34612 31340
rect 34664 31288 34670 31340
rect 28960 31232 29224 31260
rect 28960 31220 28966 31232
rect 29638 31220 29644 31272
rect 29696 31260 29702 31272
rect 32582 31260 32588 31272
rect 29696 31232 32588 31260
rect 29696 31220 29702 31232
rect 32582 31220 32588 31232
rect 32640 31220 32646 31272
rect 33134 31220 33140 31272
rect 33192 31220 33198 31272
rect 26206 31164 27016 31192
rect 19904 31096 21220 31124
rect 19797 31087 19855 31093
rect 25866 31084 25872 31136
rect 25924 31084 25930 31136
rect 27890 31084 27896 31136
rect 27948 31124 27954 31136
rect 28721 31127 28779 31133
rect 28721 31124 28733 31127
rect 27948 31096 28733 31124
rect 27948 31084 27954 31096
rect 28721 31093 28733 31096
rect 28767 31093 28779 31127
rect 28721 31087 28779 31093
rect 1104 31034 37076 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 37076 31034
rect 1104 30960 37076 30982
rect 8938 30880 8944 30932
rect 8996 30880 9002 30932
rect 13354 30880 13360 30932
rect 13412 30920 13418 30932
rect 16390 30920 16396 30932
rect 13412 30892 16396 30920
rect 13412 30880 13418 30892
rect 5626 30784 5632 30796
rect 3896 30756 5632 30784
rect 3510 30676 3516 30728
rect 3568 30716 3574 30728
rect 3896 30725 3924 30756
rect 5626 30744 5632 30756
rect 5684 30744 5690 30796
rect 6641 30787 6699 30793
rect 6641 30753 6653 30787
rect 6687 30784 6699 30787
rect 6733 30787 6791 30793
rect 6733 30784 6745 30787
rect 6687 30756 6745 30784
rect 6687 30753 6699 30756
rect 6641 30747 6699 30753
rect 6733 30753 6745 30756
rect 6779 30784 6791 30787
rect 8202 30784 8208 30796
rect 6779 30756 8208 30784
rect 6779 30753 6791 30756
rect 6733 30747 6791 30753
rect 8202 30744 8208 30756
rect 8260 30744 8266 30796
rect 8570 30744 8576 30796
rect 8628 30784 8634 30796
rect 13464 30793 13492 30892
rect 16390 30880 16396 30892
rect 16448 30880 16454 30932
rect 18322 30880 18328 30932
rect 18380 30920 18386 30932
rect 19245 30923 19303 30929
rect 19245 30920 19257 30923
rect 18380 30892 19257 30920
rect 18380 30880 18386 30892
rect 19245 30889 19257 30892
rect 19291 30889 19303 30923
rect 19245 30883 19303 30889
rect 20162 30880 20168 30932
rect 20220 30920 20226 30932
rect 20349 30923 20407 30929
rect 20349 30920 20361 30923
rect 20220 30892 20361 30920
rect 20220 30880 20226 30892
rect 20349 30889 20361 30892
rect 20395 30889 20407 30923
rect 20349 30883 20407 30889
rect 22462 30880 22468 30932
rect 22520 30920 22526 30932
rect 26145 30923 26203 30929
rect 22520 30892 25728 30920
rect 22520 30880 22526 30892
rect 19334 30812 19340 30864
rect 19392 30852 19398 30864
rect 20254 30852 20260 30864
rect 19392 30824 20260 30852
rect 19392 30812 19398 30824
rect 9493 30787 9551 30793
rect 9493 30784 9505 30787
rect 8628 30756 9505 30784
rect 8628 30744 8634 30756
rect 9493 30753 9505 30756
rect 9539 30753 9551 30787
rect 9493 30747 9551 30753
rect 13449 30787 13507 30793
rect 13449 30753 13461 30787
rect 13495 30753 13507 30787
rect 13449 30747 13507 30753
rect 15286 30744 15292 30796
rect 15344 30784 15350 30796
rect 15473 30787 15531 30793
rect 15473 30784 15485 30787
rect 15344 30756 15485 30784
rect 15344 30744 15350 30756
rect 15473 30753 15485 30756
rect 15519 30784 15531 30787
rect 16482 30784 16488 30796
rect 15519 30756 16488 30784
rect 15519 30753 15531 30756
rect 15473 30747 15531 30753
rect 16482 30744 16488 30756
rect 16540 30784 16546 30796
rect 17313 30787 17371 30793
rect 17313 30784 17325 30787
rect 16540 30756 17325 30784
rect 16540 30744 16546 30756
rect 17313 30753 17325 30756
rect 17359 30753 17371 30787
rect 17313 30747 17371 30753
rect 18230 30744 18236 30796
rect 18288 30784 18294 30796
rect 19904 30793 19932 30824
rect 20254 30812 20260 30824
rect 20312 30852 20318 30864
rect 22480 30852 22508 30880
rect 20312 30824 22508 30852
rect 25700 30852 25728 30892
rect 26145 30889 26157 30923
rect 26191 30920 26203 30923
rect 26326 30920 26332 30932
rect 26191 30892 26332 30920
rect 26191 30889 26203 30892
rect 26145 30883 26203 30889
rect 26326 30880 26332 30892
rect 26384 30880 26390 30932
rect 26973 30923 27031 30929
rect 26973 30889 26985 30923
rect 27019 30920 27031 30923
rect 27246 30920 27252 30932
rect 27019 30892 27252 30920
rect 27019 30889 27031 30892
rect 26973 30883 27031 30889
rect 27246 30880 27252 30892
rect 27304 30880 27310 30932
rect 29812 30923 29870 30929
rect 29812 30889 29824 30923
rect 29858 30920 29870 30923
rect 30374 30920 30380 30932
rect 29858 30892 30380 30920
rect 29858 30889 29870 30892
rect 29812 30883 29870 30889
rect 30374 30880 30380 30892
rect 30432 30880 30438 30932
rect 31110 30880 31116 30932
rect 31168 30920 31174 30932
rect 31297 30923 31355 30929
rect 31297 30920 31309 30923
rect 31168 30892 31309 30920
rect 31168 30880 31174 30892
rect 31297 30889 31309 30892
rect 31343 30889 31355 30923
rect 31297 30883 31355 30889
rect 26510 30852 26516 30864
rect 25700 30824 26516 30852
rect 20312 30812 20318 30824
rect 26510 30812 26516 30824
rect 26568 30812 26574 30864
rect 33042 30852 33048 30864
rect 32048 30824 33048 30852
rect 19061 30787 19119 30793
rect 19061 30784 19073 30787
rect 18288 30756 19073 30784
rect 18288 30744 18294 30756
rect 19061 30753 19073 30756
rect 19107 30784 19119 30787
rect 19705 30787 19763 30793
rect 19705 30784 19717 30787
rect 19107 30756 19717 30784
rect 19107 30753 19119 30756
rect 19061 30747 19119 30753
rect 19705 30753 19717 30756
rect 19751 30753 19763 30787
rect 19705 30747 19763 30753
rect 19889 30787 19947 30793
rect 19889 30753 19901 30787
rect 19935 30753 19947 30787
rect 19889 30747 19947 30753
rect 20898 30744 20904 30796
rect 20956 30744 20962 30796
rect 24673 30787 24731 30793
rect 24673 30753 24685 30787
rect 24719 30784 24731 30787
rect 25866 30784 25872 30796
rect 24719 30756 25872 30784
rect 24719 30753 24731 30756
rect 24673 30747 24731 30753
rect 25866 30744 25872 30756
rect 25924 30744 25930 30796
rect 27525 30787 27583 30793
rect 27525 30753 27537 30787
rect 27571 30784 27583 30787
rect 27982 30784 27988 30796
rect 27571 30756 27988 30784
rect 27571 30753 27583 30756
rect 27525 30747 27583 30753
rect 27982 30744 27988 30756
rect 28040 30744 28046 30796
rect 29549 30787 29607 30793
rect 29549 30753 29561 30787
rect 29595 30784 29607 30787
rect 30558 30784 30564 30796
rect 29595 30756 30564 30784
rect 29595 30753 29607 30756
rect 29549 30747 29607 30753
rect 30558 30744 30564 30756
rect 30616 30744 30622 30796
rect 32048 30793 32076 30824
rect 33042 30812 33048 30824
rect 33100 30812 33106 30864
rect 32033 30787 32091 30793
rect 32033 30753 32045 30787
rect 32079 30753 32091 30787
rect 32033 30747 32091 30753
rect 32398 30744 32404 30796
rect 32456 30784 32462 30796
rect 34977 30787 35035 30793
rect 34977 30784 34989 30787
rect 32456 30756 34989 30784
rect 32456 30744 32462 30756
rect 34977 30753 34989 30756
rect 35023 30753 35035 30787
rect 34977 30747 35035 30753
rect 3881 30719 3939 30725
rect 3881 30716 3893 30719
rect 3568 30688 3893 30716
rect 3568 30676 3574 30688
rect 3881 30685 3893 30688
rect 3927 30685 3939 30719
rect 3881 30679 3939 30685
rect 4065 30719 4123 30725
rect 4065 30685 4077 30719
rect 4111 30716 4123 30719
rect 4614 30716 4620 30728
rect 4111 30688 4620 30716
rect 4111 30685 4123 30688
rect 4065 30679 4123 30685
rect 4614 30676 4620 30688
rect 4672 30676 4678 30728
rect 9766 30676 9772 30728
rect 9824 30676 9830 30728
rect 9950 30676 9956 30728
rect 10008 30676 10014 30728
rect 19610 30676 19616 30728
rect 19668 30716 19674 30728
rect 20809 30719 20867 30725
rect 20809 30716 20821 30719
rect 19668 30688 20821 30716
rect 19668 30676 19674 30688
rect 20809 30685 20821 30688
rect 20855 30685 20867 30719
rect 20809 30679 20867 30685
rect 24394 30676 24400 30728
rect 24452 30676 24458 30728
rect 27341 30719 27399 30725
rect 27341 30685 27353 30719
rect 27387 30716 27399 30719
rect 27890 30716 27896 30728
rect 27387 30688 27896 30716
rect 27387 30685 27399 30688
rect 27341 30679 27399 30685
rect 27890 30676 27896 30688
rect 27948 30676 27954 30728
rect 31849 30719 31907 30725
rect 31849 30685 31861 30719
rect 31895 30716 31907 30719
rect 32416 30716 32444 30744
rect 31895 30688 32444 30716
rect 31895 30685 31907 30688
rect 31849 30679 31907 30685
rect 32582 30676 32588 30728
rect 32640 30676 32646 30728
rect 33594 30676 33600 30728
rect 33652 30676 33658 30728
rect 34606 30676 34612 30728
rect 34664 30716 34670 30728
rect 35069 30719 35127 30725
rect 35069 30716 35081 30719
rect 34664 30688 35081 30716
rect 34664 30676 34670 30688
rect 35069 30685 35081 30688
rect 35115 30685 35127 30719
rect 35069 30679 35127 30685
rect 35253 30719 35311 30725
rect 35253 30685 35265 30719
rect 35299 30716 35311 30719
rect 35342 30716 35348 30728
rect 35299 30688 35348 30716
rect 35299 30685 35311 30688
rect 35253 30679 35311 30685
rect 35342 30676 35348 30688
rect 35400 30676 35406 30728
rect 4706 30608 4712 30660
rect 4764 30648 4770 30660
rect 4764 30620 5198 30648
rect 4764 30608 4770 30620
rect 6362 30608 6368 30660
rect 6420 30608 6426 30660
rect 7009 30651 7067 30657
rect 7009 30617 7021 30651
rect 7055 30617 7067 30651
rect 7009 30611 7067 30617
rect 3973 30583 4031 30589
rect 3973 30549 3985 30583
rect 4019 30580 4031 30583
rect 4154 30580 4160 30592
rect 4019 30552 4160 30580
rect 4019 30549 4031 30552
rect 3973 30543 4031 30549
rect 4154 30540 4160 30552
rect 4212 30540 4218 30592
rect 4893 30583 4951 30589
rect 4893 30549 4905 30583
rect 4939 30580 4951 30583
rect 6730 30580 6736 30592
rect 4939 30552 6736 30580
rect 4939 30549 4951 30552
rect 4893 30543 4951 30549
rect 6730 30540 6736 30552
rect 6788 30540 6794 30592
rect 7024 30580 7052 30611
rect 7466 30608 7472 30660
rect 7524 30608 7530 30660
rect 9309 30651 9367 30657
rect 9309 30617 9321 30651
rect 9355 30648 9367 30651
rect 9861 30651 9919 30657
rect 9861 30648 9873 30651
rect 9355 30620 9873 30648
rect 9355 30617 9367 30620
rect 9309 30611 9367 30617
rect 9861 30617 9873 30620
rect 9907 30617 9919 30651
rect 9861 30611 9919 30617
rect 8294 30580 8300 30592
rect 7024 30552 8300 30580
rect 8294 30540 8300 30552
rect 8352 30540 8358 30592
rect 8478 30540 8484 30592
rect 8536 30540 8542 30592
rect 9401 30583 9459 30589
rect 9401 30549 9413 30583
rect 9447 30580 9459 30583
rect 9968 30580 9996 30676
rect 15749 30651 15807 30657
rect 15749 30617 15761 30651
rect 15795 30648 15807 30651
rect 16022 30648 16028 30660
rect 15795 30620 16028 30648
rect 15795 30617 15807 30620
rect 15749 30611 15807 30617
rect 16022 30608 16028 30620
rect 16080 30608 16086 30660
rect 16298 30608 16304 30660
rect 16356 30608 16362 30660
rect 17586 30608 17592 30660
rect 17644 30608 17650 30660
rect 18874 30648 18880 30660
rect 18814 30620 18880 30648
rect 18874 30608 18880 30620
rect 18932 30608 18938 30660
rect 20717 30651 20775 30657
rect 20717 30617 20729 30651
rect 20763 30648 20775 30651
rect 22094 30648 22100 30660
rect 20763 30620 22100 30648
rect 20763 30617 20775 30620
rect 20717 30611 20775 30617
rect 22094 30608 22100 30620
rect 22152 30608 22158 30660
rect 25222 30608 25228 30660
rect 25280 30608 25286 30660
rect 28902 30608 28908 30660
rect 28960 30648 28966 30660
rect 31110 30648 31116 30660
rect 28960 30620 30236 30648
rect 31050 30620 31116 30648
rect 28960 30608 28966 30620
rect 9447 30552 9996 30580
rect 9447 30549 9459 30552
rect 9401 30543 9459 30549
rect 12618 30540 12624 30592
rect 12676 30580 12682 30592
rect 12805 30583 12863 30589
rect 12805 30580 12817 30583
rect 12676 30552 12817 30580
rect 12676 30540 12682 30552
rect 12805 30549 12817 30552
rect 12851 30549 12863 30583
rect 12805 30543 12863 30549
rect 13170 30540 13176 30592
rect 13228 30540 13234 30592
rect 13265 30583 13323 30589
rect 13265 30549 13277 30583
rect 13311 30580 13323 30583
rect 13722 30580 13728 30592
rect 13311 30552 13728 30580
rect 13311 30549 13323 30552
rect 13265 30543 13323 30549
rect 13722 30540 13728 30552
rect 13780 30540 13786 30592
rect 17221 30583 17279 30589
rect 17221 30549 17233 30583
rect 17267 30580 17279 30583
rect 17954 30580 17960 30592
rect 17267 30552 17960 30580
rect 17267 30549 17279 30552
rect 17221 30543 17279 30549
rect 17954 30540 17960 30552
rect 18012 30580 18018 30592
rect 18322 30580 18328 30592
rect 18012 30552 18328 30580
rect 18012 30540 18018 30552
rect 18322 30540 18328 30552
rect 18380 30540 18386 30592
rect 18892 30580 18920 30608
rect 20806 30580 20812 30592
rect 18892 30552 20812 30580
rect 20806 30540 20812 30552
rect 20864 30540 20870 30592
rect 27433 30583 27491 30589
rect 27433 30549 27445 30583
rect 27479 30580 27491 30583
rect 27614 30580 27620 30592
rect 27479 30552 27620 30580
rect 27479 30549 27491 30552
rect 27433 30543 27491 30549
rect 27614 30540 27620 30552
rect 27672 30540 27678 30592
rect 30208 30580 30236 30620
rect 31110 30608 31116 30620
rect 31168 30648 31174 30660
rect 31570 30648 31576 30660
rect 31168 30620 31576 30648
rect 31168 30608 31174 30620
rect 31570 30608 31576 30620
rect 31628 30608 31634 30660
rect 31757 30651 31815 30657
rect 31757 30617 31769 30651
rect 31803 30648 31815 30651
rect 31938 30648 31944 30660
rect 31803 30620 31944 30648
rect 31803 30617 31815 30620
rect 31757 30611 31815 30617
rect 31938 30608 31944 30620
rect 31996 30608 32002 30660
rect 34514 30608 34520 30660
rect 34572 30648 34578 30660
rect 35713 30651 35771 30657
rect 35713 30648 35725 30651
rect 34572 30620 35725 30648
rect 34572 30608 34578 30620
rect 35713 30617 35725 30620
rect 35759 30617 35771 30651
rect 35713 30611 35771 30617
rect 31128 30580 31156 30608
rect 30208 30552 31156 30580
rect 31389 30583 31447 30589
rect 31389 30549 31401 30583
rect 31435 30580 31447 30583
rect 31478 30580 31484 30592
rect 31435 30552 31484 30580
rect 31435 30549 31447 30552
rect 31389 30543 31447 30549
rect 31478 30540 31484 30552
rect 31536 30540 31542 30592
rect 1104 30490 37076 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 37076 30490
rect 1104 30416 37076 30438
rect 4706 30376 4712 30388
rect 4080 30348 4712 30376
rect 4080 30308 4108 30348
rect 4706 30336 4712 30348
rect 4764 30376 4770 30388
rect 4764 30348 5488 30376
rect 4764 30336 4770 30348
rect 5460 30308 5488 30348
rect 6362 30336 6368 30388
rect 6420 30336 6426 30388
rect 8570 30376 8576 30388
rect 8312 30348 8576 30376
rect 5902 30308 5908 30320
rect 2746 30280 4186 30308
rect 5460 30280 5908 30308
rect 1765 30243 1823 30249
rect 1765 30209 1777 30243
rect 1811 30240 1823 30243
rect 2590 30240 2596 30252
rect 1811 30212 2596 30240
rect 1811 30209 1823 30212
rect 1765 30203 1823 30209
rect 2590 30200 2596 30212
rect 2648 30240 2654 30252
rect 2746 30240 2774 30280
rect 5902 30268 5908 30280
rect 5960 30308 5966 30320
rect 7466 30308 7472 30320
rect 5960 30280 7472 30308
rect 5960 30268 5966 30280
rect 7466 30268 7472 30280
rect 7524 30268 7530 30320
rect 8312 30317 8340 30348
rect 8570 30336 8576 30348
rect 8628 30336 8634 30388
rect 9217 30379 9275 30385
rect 9217 30345 9229 30379
rect 9263 30376 9275 30379
rect 9582 30376 9588 30388
rect 9263 30348 9588 30376
rect 9263 30345 9275 30348
rect 9217 30339 9275 30345
rect 9582 30336 9588 30348
rect 9640 30336 9646 30388
rect 16206 30376 16212 30388
rect 13924 30348 14872 30376
rect 8754 30317 8760 30320
rect 8297 30311 8355 30317
rect 8297 30277 8309 30311
rect 8343 30277 8355 30311
rect 8297 30271 8355 30277
rect 8741 30311 8760 30317
rect 8741 30277 8753 30311
rect 8741 30271 8760 30277
rect 8754 30268 8760 30271
rect 8812 30268 8818 30320
rect 8941 30311 8999 30317
rect 8941 30277 8953 30311
rect 8987 30277 8999 30311
rect 8941 30271 8999 30277
rect 9309 30311 9367 30317
rect 9309 30277 9321 30311
rect 9355 30308 9367 30311
rect 9674 30308 9680 30320
rect 9355 30280 9680 30308
rect 9355 30277 9367 30280
rect 9309 30271 9367 30277
rect 2648 30212 2774 30240
rect 2648 30200 2654 30212
rect 2958 30200 2964 30252
rect 3016 30240 3022 30252
rect 3326 30240 3332 30252
rect 3016 30212 3332 30240
rect 3016 30200 3022 30212
rect 3326 30200 3332 30212
rect 3384 30200 3390 30252
rect 5626 30200 5632 30252
rect 5684 30200 5690 30252
rect 5810 30200 5816 30252
rect 5868 30240 5874 30252
rect 6733 30243 6791 30249
rect 6733 30240 6745 30243
rect 5868 30212 6745 30240
rect 5868 30200 5874 30212
rect 6733 30209 6745 30212
rect 6779 30209 6791 30243
rect 6733 30203 6791 30209
rect 7834 30200 7840 30252
rect 7892 30240 7898 30252
rect 8021 30243 8079 30249
rect 8021 30240 8033 30243
rect 7892 30212 8033 30240
rect 7892 30200 7898 30212
rect 8021 30209 8033 30212
rect 8067 30209 8079 30243
rect 8021 30203 8079 30209
rect 8110 30200 8116 30252
rect 8168 30200 8174 30252
rect 3421 30175 3479 30181
rect 3421 30141 3433 30175
rect 3467 30141 3479 30175
rect 3421 30135 3479 30141
rect 3697 30175 3755 30181
rect 3697 30141 3709 30175
rect 3743 30172 3755 30175
rect 3786 30172 3792 30184
rect 3743 30144 3792 30172
rect 3743 30141 3755 30144
rect 3697 30135 3755 30141
rect 3436 30036 3464 30135
rect 3786 30132 3792 30144
rect 3844 30132 3850 30184
rect 5718 30132 5724 30184
rect 5776 30172 5782 30184
rect 6825 30175 6883 30181
rect 6825 30172 6837 30175
rect 5776 30144 6837 30172
rect 5776 30132 5782 30144
rect 6825 30141 6837 30144
rect 6871 30141 6883 30175
rect 6825 30135 6883 30141
rect 6917 30175 6975 30181
rect 6917 30141 6929 30175
rect 6963 30141 6975 30175
rect 6917 30135 6975 30141
rect 6730 30064 6736 30116
rect 6788 30104 6794 30116
rect 6932 30104 6960 30135
rect 6788 30076 6960 30104
rect 6788 30064 6794 30076
rect 8294 30064 8300 30116
rect 8352 30064 8358 30116
rect 8956 30104 8984 30271
rect 9674 30268 9680 30280
rect 9732 30268 9738 30320
rect 13262 30308 13268 30320
rect 13110 30280 13268 30308
rect 13262 30268 13268 30280
rect 13320 30308 13326 30320
rect 13924 30308 13952 30348
rect 14844 30308 14872 30348
rect 15212 30348 16212 30376
rect 15212 30308 15240 30348
rect 16206 30336 16212 30348
rect 16264 30336 16270 30388
rect 17586 30336 17592 30388
rect 17644 30376 17650 30388
rect 17865 30379 17923 30385
rect 17865 30376 17877 30379
rect 17644 30348 17877 30376
rect 17644 30336 17650 30348
rect 17865 30345 17877 30348
rect 17911 30345 17923 30379
rect 17865 30339 17923 30345
rect 18230 30336 18236 30388
rect 18288 30336 18294 30388
rect 18322 30336 18328 30388
rect 18380 30336 18386 30388
rect 26326 30336 26332 30388
rect 26384 30336 26390 30388
rect 32398 30336 32404 30388
rect 32456 30336 32462 30388
rect 33502 30376 33508 30388
rect 32508 30348 33508 30376
rect 13320 30280 13952 30308
rect 14766 30280 15240 30308
rect 13320 30268 13326 30280
rect 15286 30268 15292 30320
rect 15344 30308 15350 30320
rect 15344 30280 15516 30308
rect 15344 30268 15350 30280
rect 9398 30200 9404 30252
rect 9456 30200 9462 30252
rect 10413 30243 10471 30249
rect 10413 30209 10425 30243
rect 10459 30240 10471 30243
rect 10778 30240 10784 30252
rect 10459 30212 10784 30240
rect 10459 30209 10471 30212
rect 10413 30203 10471 30209
rect 10778 30200 10784 30212
rect 10836 30200 10842 30252
rect 11606 30200 11612 30252
rect 11664 30200 11670 30252
rect 15488 30249 15516 30280
rect 22186 30268 22192 30320
rect 22244 30308 22250 30320
rect 25777 30311 25835 30317
rect 22244 30280 22494 30308
rect 22244 30268 22250 30280
rect 25777 30277 25789 30311
rect 25823 30308 25835 30311
rect 30558 30308 30564 30320
rect 25823 30280 28580 30308
rect 25823 30277 25835 30280
rect 25777 30271 25835 30277
rect 15473 30243 15531 30249
rect 15473 30209 15485 30243
rect 15519 30209 15531 30243
rect 15473 30203 15531 30209
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30240 23995 30243
rect 24394 30240 24400 30252
rect 23983 30212 24400 30240
rect 23983 30209 23995 30212
rect 23937 30203 23995 30209
rect 24394 30200 24400 30212
rect 24452 30200 24458 30252
rect 26237 30243 26295 30249
rect 26237 30209 26249 30243
rect 26283 30209 26295 30243
rect 26237 30203 26295 30209
rect 9122 30132 9128 30184
rect 9180 30172 9186 30184
rect 9766 30172 9772 30184
rect 9180 30144 9772 30172
rect 9180 30132 9186 30144
rect 9766 30132 9772 30144
rect 9824 30132 9830 30184
rect 10502 30132 10508 30184
rect 10560 30132 10566 30184
rect 10597 30175 10655 30181
rect 10597 30141 10609 30175
rect 10643 30141 10655 30175
rect 10597 30135 10655 30141
rect 11885 30175 11943 30181
rect 11885 30141 11897 30175
rect 11931 30172 11943 30175
rect 12618 30172 12624 30184
rect 11931 30144 12624 30172
rect 11931 30141 11943 30144
rect 11885 30135 11943 30141
rect 9033 30107 9091 30113
rect 9033 30104 9045 30107
rect 8956 30076 9045 30104
rect 9033 30073 9045 30076
rect 9079 30104 9091 30107
rect 9214 30104 9220 30116
rect 9079 30076 9220 30104
rect 9079 30073 9091 30076
rect 9033 30067 9091 30073
rect 9214 30064 9220 30076
rect 9272 30064 9278 30116
rect 9585 30107 9643 30113
rect 9585 30073 9597 30107
rect 9631 30104 9643 30107
rect 10612 30104 10640 30135
rect 12618 30132 12624 30144
rect 12676 30132 12682 30184
rect 15194 30132 15200 30184
rect 15252 30132 15258 30184
rect 18414 30132 18420 30184
rect 18472 30172 18478 30184
rect 20898 30172 20904 30184
rect 18472 30144 20904 30172
rect 18472 30132 18478 30144
rect 20898 30132 20904 30144
rect 20956 30132 20962 30184
rect 23658 30132 23664 30184
rect 23716 30132 23722 30184
rect 25038 30132 25044 30184
rect 25096 30172 25102 30184
rect 26252 30172 26280 30203
rect 25096 30144 26280 30172
rect 25096 30132 25102 30144
rect 26510 30132 26516 30184
rect 26568 30132 26574 30184
rect 9631 30076 10640 30104
rect 24489 30107 24547 30113
rect 9631 30073 9643 30076
rect 9585 30067 9643 30073
rect 24489 30073 24501 30107
rect 24535 30104 24547 30107
rect 24854 30104 24860 30116
rect 24535 30076 24860 30104
rect 24535 30073 24547 30076
rect 24489 30067 24547 30073
rect 24854 30064 24860 30076
rect 24912 30064 24918 30116
rect 4706 30036 4712 30048
rect 3436 30008 4712 30036
rect 4706 29996 4712 30008
rect 4764 29996 4770 30048
rect 5166 29996 5172 30048
rect 5224 29996 5230 30048
rect 8478 29996 8484 30048
rect 8536 30036 8542 30048
rect 8757 30039 8815 30045
rect 8757 30036 8769 30039
rect 8536 30008 8769 30036
rect 8536 29996 8542 30008
rect 8757 30005 8769 30008
rect 8803 30036 8815 30039
rect 9490 30036 9496 30048
rect 8803 30008 9496 30036
rect 8803 30005 8815 30008
rect 8757 29999 8815 30005
rect 9490 29996 9496 30008
rect 9548 29996 9554 30048
rect 9950 29996 9956 30048
rect 10008 30036 10014 30048
rect 10045 30039 10103 30045
rect 10045 30036 10057 30039
rect 10008 30008 10057 30036
rect 10008 29996 10014 30008
rect 10045 30005 10057 30008
rect 10091 30005 10103 30039
rect 10045 29999 10103 30005
rect 12986 29996 12992 30048
rect 13044 30036 13050 30048
rect 13170 30036 13176 30048
rect 13044 30008 13176 30036
rect 13044 29996 13050 30008
rect 13170 29996 13176 30008
rect 13228 30036 13234 30048
rect 13357 30039 13415 30045
rect 13357 30036 13369 30039
rect 13228 30008 13369 30036
rect 13228 29996 13234 30008
rect 13357 30005 13369 30008
rect 13403 30005 13415 30039
rect 13357 29999 13415 30005
rect 13722 29996 13728 30048
rect 13780 29996 13786 30048
rect 22189 30039 22247 30045
rect 22189 30005 22201 30039
rect 22235 30036 22247 30039
rect 22554 30036 22560 30048
rect 22235 30008 22560 30036
rect 22235 30005 22247 30008
rect 22189 29999 22247 30005
rect 22554 29996 22560 30008
rect 22612 29996 22618 30048
rect 25866 29996 25872 30048
rect 25924 29996 25930 30048
rect 28552 30036 28580 30280
rect 30208 30280 30564 30308
rect 30208 30249 30236 30280
rect 30558 30268 30564 30280
rect 30616 30268 30622 30320
rect 30193 30243 30251 30249
rect 30193 30209 30205 30243
rect 30239 30209 30251 30243
rect 30193 30203 30251 30209
rect 31570 30200 31576 30252
rect 31628 30240 31634 30252
rect 32508 30240 32536 30348
rect 33502 30336 33508 30348
rect 33560 30376 33566 30388
rect 33962 30376 33968 30388
rect 33560 30348 33968 30376
rect 33560 30336 33566 30348
rect 33962 30336 33968 30348
rect 34020 30336 34026 30388
rect 33520 30308 33548 30336
rect 33442 30280 33548 30308
rect 33873 30311 33931 30317
rect 33873 30277 33885 30311
rect 33919 30308 33931 30311
rect 34514 30308 34520 30320
rect 33919 30280 34520 30308
rect 33919 30277 33931 30280
rect 33873 30271 33931 30277
rect 34514 30268 34520 30280
rect 34572 30268 34578 30320
rect 31628 30212 32536 30240
rect 31628 30200 31634 30212
rect 34146 30200 34152 30252
rect 34204 30200 34210 30252
rect 30469 30175 30527 30181
rect 30469 30141 30481 30175
rect 30515 30172 30527 30175
rect 31478 30172 31484 30184
rect 30515 30144 31484 30172
rect 30515 30141 30527 30144
rect 30469 30135 30527 30141
rect 31478 30132 31484 30144
rect 31536 30132 31542 30184
rect 30834 30036 30840 30048
rect 28552 30008 30840 30036
rect 30834 29996 30840 30008
rect 30892 29996 30898 30048
rect 31938 29996 31944 30048
rect 31996 29996 32002 30048
rect 1104 29946 37076 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 37076 29946
rect 1104 29872 37076 29894
rect 3786 29792 3792 29844
rect 3844 29792 3850 29844
rect 4522 29792 4528 29844
rect 4580 29832 4586 29844
rect 5166 29832 5172 29844
rect 4580 29804 5172 29832
rect 4580 29792 4586 29804
rect 5166 29792 5172 29804
rect 5224 29792 5230 29844
rect 7834 29792 7840 29844
rect 7892 29792 7898 29844
rect 8110 29792 8116 29844
rect 8168 29792 8174 29844
rect 8202 29792 8208 29844
rect 8260 29832 8266 29844
rect 8260 29804 8800 29832
rect 8260 29792 8266 29804
rect 4617 29767 4675 29773
rect 4617 29764 4629 29767
rect 3712 29736 4629 29764
rect 2133 29699 2191 29705
rect 2133 29665 2145 29699
rect 2179 29696 2191 29699
rect 3712 29696 3740 29736
rect 4617 29733 4629 29736
rect 4663 29733 4675 29767
rect 8478 29764 8484 29776
rect 4617 29727 4675 29733
rect 7944 29736 8484 29764
rect 2179 29668 3740 29696
rect 4433 29699 4491 29705
rect 2179 29665 2191 29668
rect 2133 29659 2191 29665
rect 4433 29665 4445 29699
rect 4479 29696 4491 29699
rect 4522 29696 4528 29708
rect 4479 29668 4528 29696
rect 4479 29665 4491 29668
rect 4433 29659 4491 29665
rect 4522 29656 4528 29668
rect 4580 29656 4586 29708
rect 4706 29656 4712 29708
rect 4764 29696 4770 29708
rect 5169 29699 5227 29705
rect 5169 29696 5181 29699
rect 4764 29668 5181 29696
rect 4764 29656 4770 29668
rect 5169 29665 5181 29668
rect 5215 29665 5227 29699
rect 5169 29659 5227 29665
rect 1394 29588 1400 29640
rect 1452 29628 1458 29640
rect 1857 29631 1915 29637
rect 1857 29628 1869 29631
rect 1452 29600 1869 29628
rect 1452 29588 1458 29600
rect 1857 29597 1869 29600
rect 1903 29597 1915 29631
rect 1857 29591 1915 29597
rect 4157 29631 4215 29637
rect 4157 29597 4169 29631
rect 4203 29628 4215 29631
rect 4246 29628 4252 29640
rect 4203 29600 4252 29628
rect 4203 29597 4215 29600
rect 4157 29591 4215 29597
rect 4246 29588 4252 29600
rect 4304 29628 4310 29640
rect 4614 29628 4620 29640
rect 4304 29600 4620 29628
rect 4304 29588 4310 29600
rect 4614 29588 4620 29600
rect 4672 29588 4678 29640
rect 4801 29631 4859 29637
rect 4801 29597 4813 29631
rect 4847 29597 4859 29631
rect 4801 29591 4859 29597
rect 2590 29520 2596 29572
rect 2648 29520 2654 29572
rect 4816 29560 4844 29591
rect 4890 29588 4896 29640
rect 4948 29588 4954 29640
rect 7944 29637 7972 29736
rect 8478 29724 8484 29736
rect 8536 29724 8542 29776
rect 8772 29696 8800 29804
rect 15194 29792 15200 29844
rect 15252 29832 15258 29844
rect 15289 29835 15347 29841
rect 15289 29832 15301 29835
rect 15252 29804 15301 29832
rect 15252 29792 15258 29804
rect 15289 29801 15301 29804
rect 15335 29801 15347 29835
rect 15289 29795 15347 29801
rect 27614 29792 27620 29844
rect 27672 29832 27678 29844
rect 27672 29804 28120 29832
rect 27672 29792 27678 29804
rect 24762 29724 24768 29776
rect 24820 29764 24826 29776
rect 24820 29736 25176 29764
rect 24820 29724 24826 29736
rect 9677 29699 9735 29705
rect 9677 29696 9689 29699
rect 8220 29668 8708 29696
rect 8772 29668 9689 29696
rect 8220 29637 8248 29668
rect 7745 29631 7803 29637
rect 7745 29597 7757 29631
rect 7791 29597 7803 29631
rect 7745 29591 7803 29597
rect 7929 29631 7987 29637
rect 7929 29597 7941 29631
rect 7975 29597 7987 29631
rect 7929 29591 7987 29597
rect 8021 29631 8079 29637
rect 8021 29597 8033 29631
rect 8067 29597 8079 29631
rect 8021 29591 8079 29597
rect 8205 29631 8263 29637
rect 8205 29597 8217 29631
rect 8251 29597 8263 29631
rect 8205 29591 8263 29597
rect 4264 29532 4844 29560
rect 5445 29563 5503 29569
rect 3602 29452 3608 29504
rect 3660 29452 3666 29504
rect 4154 29452 4160 29504
rect 4212 29492 4218 29504
rect 4264 29501 4292 29532
rect 5445 29529 5457 29563
rect 5491 29560 5503 29563
rect 5534 29560 5540 29572
rect 5491 29532 5540 29560
rect 5491 29529 5503 29532
rect 5445 29523 5503 29529
rect 5534 29520 5540 29532
rect 5592 29520 5598 29572
rect 5902 29520 5908 29572
rect 5960 29520 5966 29572
rect 4249 29495 4307 29501
rect 4249 29492 4261 29495
rect 4212 29464 4261 29492
rect 4212 29452 4218 29464
rect 4249 29461 4261 29464
rect 4295 29461 4307 29495
rect 4249 29455 4307 29461
rect 6086 29452 6092 29504
rect 6144 29492 6150 29504
rect 6917 29495 6975 29501
rect 6917 29492 6929 29495
rect 6144 29464 6929 29492
rect 6144 29452 6150 29464
rect 6917 29461 6929 29464
rect 6963 29461 6975 29495
rect 7760 29492 7788 29591
rect 8036 29560 8064 29591
rect 8294 29588 8300 29640
rect 8352 29588 8358 29640
rect 8478 29588 8484 29640
rect 8536 29588 8542 29640
rect 8680 29637 8708 29668
rect 9677 29665 9689 29668
rect 9723 29665 9735 29699
rect 9677 29659 9735 29665
rect 9950 29656 9956 29708
rect 10008 29656 10014 29708
rect 10410 29656 10416 29708
rect 10468 29696 10474 29708
rect 10468 29668 11376 29696
rect 10468 29656 10474 29668
rect 8665 29631 8723 29637
rect 8665 29597 8677 29631
rect 8711 29628 8723 29631
rect 9214 29628 9220 29640
rect 8711 29600 9220 29628
rect 8711 29597 8723 29600
rect 8665 29591 8723 29597
rect 9214 29588 9220 29600
rect 9272 29588 9278 29640
rect 8754 29560 8760 29572
rect 8036 29532 8760 29560
rect 8754 29520 8760 29532
rect 8812 29560 8818 29572
rect 9398 29560 9404 29572
rect 8812 29532 9404 29560
rect 8812 29520 8818 29532
rect 9398 29520 9404 29532
rect 9456 29520 9462 29572
rect 10410 29560 10416 29572
rect 9784 29532 10416 29560
rect 8478 29492 8484 29504
rect 7760 29464 8484 29492
rect 6917 29455 6975 29461
rect 8478 29452 8484 29464
rect 8536 29492 8542 29504
rect 9122 29492 9128 29504
rect 8536 29464 9128 29492
rect 8536 29452 8542 29464
rect 9122 29452 9128 29464
rect 9180 29452 9186 29504
rect 9306 29452 9312 29504
rect 9364 29492 9370 29504
rect 9493 29495 9551 29501
rect 9493 29492 9505 29495
rect 9364 29464 9505 29492
rect 9364 29452 9370 29464
rect 9493 29461 9505 29464
rect 9539 29492 9551 29495
rect 9784 29492 9812 29532
rect 10410 29520 10416 29532
rect 10468 29520 10474 29572
rect 11348 29560 11376 29668
rect 13814 29656 13820 29708
rect 13872 29696 13878 29708
rect 14642 29696 14648 29708
rect 13872 29668 14648 29696
rect 13872 29656 13878 29668
rect 14642 29656 14648 29668
rect 14700 29656 14706 29708
rect 16482 29656 16488 29708
rect 16540 29696 16546 29708
rect 17497 29699 17555 29705
rect 17497 29696 17509 29699
rect 16540 29668 17509 29696
rect 16540 29656 16546 29668
rect 17497 29665 17509 29668
rect 17543 29665 17555 29699
rect 17497 29659 17555 29665
rect 20898 29656 20904 29708
rect 20956 29696 20962 29708
rect 24780 29696 24808 29724
rect 20956 29668 24808 29696
rect 20956 29656 20962 29668
rect 25038 29656 25044 29708
rect 25096 29656 25102 29708
rect 25148 29705 25176 29736
rect 25222 29724 25228 29776
rect 25280 29764 25286 29776
rect 27709 29767 27767 29773
rect 27709 29764 27721 29767
rect 25280 29736 25636 29764
rect 25280 29724 25286 29736
rect 25133 29699 25191 29705
rect 25133 29665 25145 29699
rect 25179 29696 25191 29699
rect 25179 29668 25544 29696
rect 25179 29665 25191 29668
rect 25133 29659 25191 29665
rect 11514 29588 11520 29640
rect 11572 29588 11578 29640
rect 13262 29628 13268 29640
rect 12926 29614 13268 29628
rect 12912 29600 13268 29614
rect 11348 29532 11560 29560
rect 9539 29464 9812 29492
rect 9539 29461 9551 29464
rect 9493 29455 9551 29461
rect 10594 29452 10600 29504
rect 10652 29492 10658 29504
rect 11425 29495 11483 29501
rect 11425 29492 11437 29495
rect 10652 29464 11437 29492
rect 10652 29452 10658 29464
rect 11425 29461 11437 29464
rect 11471 29461 11483 29495
rect 11532 29492 11560 29532
rect 11790 29520 11796 29572
rect 11848 29520 11854 29572
rect 12912 29492 12940 29600
rect 13262 29588 13268 29600
rect 13320 29588 13326 29640
rect 13722 29588 13728 29640
rect 13780 29628 13786 29640
rect 14921 29631 14979 29637
rect 14921 29628 14933 29631
rect 13780 29600 14933 29628
rect 13780 29588 13786 29600
rect 14921 29597 14933 29600
rect 14967 29597 14979 29631
rect 14921 29591 14979 29597
rect 19242 29588 19248 29640
rect 19300 29588 19306 29640
rect 20806 29628 20812 29640
rect 20654 29600 20812 29628
rect 20806 29588 20812 29600
rect 20864 29628 20870 29640
rect 21177 29631 21235 29637
rect 21177 29628 21189 29631
rect 20864 29600 21189 29628
rect 20864 29588 20870 29600
rect 21177 29597 21189 29600
rect 21223 29628 21235 29631
rect 21361 29631 21419 29637
rect 21361 29628 21373 29631
rect 21223 29600 21373 29628
rect 21223 29597 21235 29600
rect 21177 29591 21235 29597
rect 21361 29597 21373 29600
rect 21407 29628 21419 29631
rect 22186 29628 22192 29640
rect 21407 29600 22192 29628
rect 21407 29597 21419 29600
rect 21361 29591 21419 29597
rect 22186 29588 22192 29600
rect 22244 29588 22250 29640
rect 23569 29631 23627 29637
rect 23569 29597 23581 29631
rect 23615 29628 23627 29631
rect 25406 29628 25412 29640
rect 23615 29600 25412 29628
rect 23615 29597 23627 29600
rect 23569 29591 23627 29597
rect 25406 29588 25412 29600
rect 25464 29588 25470 29640
rect 16206 29520 16212 29572
rect 16264 29520 16270 29572
rect 17218 29520 17224 29572
rect 17276 29520 17282 29572
rect 19518 29520 19524 29572
rect 19576 29520 19582 29572
rect 23290 29520 23296 29572
rect 23348 29520 23354 29572
rect 25130 29560 25136 29572
rect 24596 29532 25136 29560
rect 11532 29464 12940 29492
rect 11425 29455 11483 29461
rect 13262 29452 13268 29504
rect 13320 29452 13326 29504
rect 14829 29495 14887 29501
rect 14829 29461 14841 29495
rect 14875 29492 14887 29495
rect 15654 29492 15660 29504
rect 14875 29464 15660 29492
rect 14875 29461 14887 29464
rect 14829 29455 14887 29461
rect 15654 29452 15660 29464
rect 15712 29452 15718 29504
rect 15746 29452 15752 29504
rect 15804 29452 15810 29504
rect 20162 29452 20168 29504
rect 20220 29492 20226 29504
rect 20993 29495 21051 29501
rect 20993 29492 21005 29495
rect 20220 29464 21005 29492
rect 20220 29452 20226 29464
rect 20993 29461 21005 29464
rect 21039 29461 21051 29495
rect 20993 29455 21051 29461
rect 21821 29495 21879 29501
rect 21821 29461 21833 29495
rect 21867 29492 21879 29495
rect 22646 29492 22652 29504
rect 21867 29464 22652 29492
rect 21867 29461 21879 29464
rect 21821 29455 21879 29461
rect 22646 29452 22652 29464
rect 22704 29452 22710 29504
rect 24596 29501 24624 29532
rect 25130 29520 25136 29532
rect 25188 29520 25194 29572
rect 24581 29495 24639 29501
rect 24581 29461 24593 29495
rect 24627 29461 24639 29495
rect 24581 29455 24639 29461
rect 24762 29452 24768 29504
rect 24820 29492 24826 29504
rect 24949 29495 25007 29501
rect 24949 29492 24961 29495
rect 24820 29464 24961 29492
rect 24820 29452 24826 29464
rect 24949 29461 24961 29464
rect 24995 29461 25007 29495
rect 25516 29492 25544 29668
rect 25608 29560 25636 29736
rect 27448 29736 27721 29764
rect 25774 29656 25780 29708
rect 25832 29696 25838 29708
rect 25869 29699 25927 29705
rect 25869 29696 25881 29699
rect 25832 29668 25881 29696
rect 25832 29656 25838 29668
rect 25869 29665 25881 29668
rect 25915 29665 25927 29699
rect 25869 29659 25927 29665
rect 26145 29699 26203 29705
rect 26145 29665 26157 29699
rect 26191 29696 26203 29699
rect 27448 29696 27476 29736
rect 27709 29733 27721 29736
rect 27755 29733 27767 29767
rect 27709 29727 27767 29733
rect 26191 29668 27476 29696
rect 26191 29665 26203 29668
rect 26145 29659 26203 29665
rect 28092 29637 28120 29804
rect 28353 29699 28411 29705
rect 28353 29665 28365 29699
rect 28399 29696 28411 29699
rect 29086 29696 29092 29708
rect 28399 29668 29092 29696
rect 28399 29665 28411 29668
rect 28353 29659 28411 29665
rect 29086 29656 29092 29668
rect 29144 29696 29150 29708
rect 30193 29699 30251 29705
rect 30193 29696 30205 29699
rect 29144 29668 30205 29696
rect 29144 29656 29150 29668
rect 30193 29665 30205 29668
rect 30239 29696 30251 29699
rect 31021 29699 31079 29705
rect 31021 29696 31033 29699
rect 30239 29668 31033 29696
rect 30239 29665 30251 29668
rect 30193 29659 30251 29665
rect 31021 29665 31033 29668
rect 31067 29665 31079 29699
rect 33042 29696 33048 29708
rect 31021 29659 31079 29665
rect 32232 29668 33048 29696
rect 28077 29631 28135 29637
rect 28077 29597 28089 29631
rect 28123 29597 28135 29631
rect 28077 29591 28135 29597
rect 31754 29588 31760 29640
rect 31812 29628 31818 29640
rect 32232 29637 32260 29668
rect 33042 29656 33048 29668
rect 33100 29696 33106 29708
rect 33413 29699 33471 29705
rect 33413 29696 33425 29699
rect 33100 29668 33425 29696
rect 33100 29656 33106 29668
rect 33413 29665 33425 29668
rect 33459 29696 33471 29699
rect 33870 29696 33876 29708
rect 33459 29668 33876 29696
rect 33459 29665 33471 29668
rect 33413 29659 33471 29665
rect 33870 29656 33876 29668
rect 33928 29656 33934 29708
rect 32217 29631 32275 29637
rect 32217 29628 32229 29631
rect 31812 29600 32229 29628
rect 31812 29588 31818 29600
rect 32217 29597 32229 29600
rect 32263 29597 32275 29631
rect 32217 29591 32275 29597
rect 33229 29631 33287 29637
rect 33229 29597 33241 29631
rect 33275 29628 33287 29631
rect 34606 29628 34612 29640
rect 33275 29600 34612 29628
rect 33275 29597 33287 29600
rect 33229 29591 33287 29597
rect 34606 29588 34612 29600
rect 34664 29588 34670 29640
rect 26602 29560 26608 29572
rect 25608 29532 26608 29560
rect 26602 29520 26608 29532
rect 26660 29520 26666 29572
rect 27982 29560 27988 29572
rect 27448 29532 27988 29560
rect 27448 29492 27476 29532
rect 27982 29520 27988 29532
rect 28040 29520 28046 29572
rect 25516 29464 27476 29492
rect 24949 29455 25007 29461
rect 27614 29452 27620 29504
rect 27672 29492 27678 29504
rect 28169 29495 28227 29501
rect 28169 29492 28181 29495
rect 27672 29464 28181 29492
rect 27672 29452 27678 29464
rect 28169 29461 28181 29464
rect 28215 29461 28227 29495
rect 28169 29455 28227 29461
rect 29546 29452 29552 29504
rect 29604 29452 29610 29504
rect 29914 29452 29920 29504
rect 29972 29452 29978 29504
rect 30009 29495 30067 29501
rect 30009 29461 30021 29495
rect 30055 29492 30067 29495
rect 30098 29492 30104 29504
rect 30055 29464 30104 29492
rect 30055 29461 30067 29464
rect 30009 29455 30067 29461
rect 30098 29452 30104 29464
rect 30156 29452 30162 29504
rect 32490 29452 32496 29504
rect 32548 29492 32554 29504
rect 32861 29495 32919 29501
rect 32861 29492 32873 29495
rect 32548 29464 32873 29492
rect 32548 29452 32554 29464
rect 32861 29461 32873 29464
rect 32907 29461 32919 29495
rect 32861 29455 32919 29461
rect 33321 29495 33379 29501
rect 33321 29461 33333 29495
rect 33367 29492 33379 29495
rect 33410 29492 33416 29504
rect 33367 29464 33416 29492
rect 33367 29461 33379 29464
rect 33321 29455 33379 29461
rect 33410 29452 33416 29464
rect 33468 29452 33474 29504
rect 1104 29402 37076 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 37076 29402
rect 1104 29328 37076 29350
rect 3145 29291 3203 29297
rect 3145 29257 3157 29291
rect 3191 29288 3203 29291
rect 3191 29260 3924 29288
rect 3191 29257 3203 29260
rect 3145 29251 3203 29257
rect 2958 29220 2964 29232
rect 2898 29192 2964 29220
rect 2958 29180 2964 29192
rect 3016 29180 3022 29232
rect 3896 29229 3924 29260
rect 4246 29248 4252 29300
rect 4304 29248 4310 29300
rect 5445 29291 5503 29297
rect 5445 29257 5457 29291
rect 5491 29257 5503 29291
rect 5445 29251 5503 29257
rect 3881 29223 3939 29229
rect 3881 29189 3893 29223
rect 3927 29220 3939 29223
rect 3970 29220 3976 29232
rect 3927 29192 3976 29220
rect 3927 29189 3939 29192
rect 3881 29183 3939 29189
rect 3970 29180 3976 29192
rect 4028 29180 4034 29232
rect 5350 29229 5356 29232
rect 4081 29223 4139 29229
rect 4081 29220 4093 29223
rect 4080 29189 4093 29220
rect 4127 29189 4139 29223
rect 4080 29183 4139 29189
rect 5077 29223 5135 29229
rect 5077 29189 5089 29223
rect 5123 29189 5135 29223
rect 5077 29183 5135 29189
rect 5293 29223 5356 29229
rect 5293 29189 5305 29223
rect 5339 29189 5356 29223
rect 5293 29183 5356 29189
rect 1394 29044 1400 29096
rect 1452 29044 1458 29096
rect 1670 29044 1676 29096
rect 1728 29044 1734 29096
rect 2866 28976 2872 29028
rect 2924 29016 2930 29028
rect 4080 29016 4108 29183
rect 5092 29084 5120 29183
rect 5350 29180 5356 29183
rect 5408 29180 5414 29232
rect 5460 29220 5488 29251
rect 5534 29248 5540 29300
rect 5592 29248 5598 29300
rect 5902 29248 5908 29300
rect 5960 29288 5966 29300
rect 6454 29288 6460 29300
rect 5960 29260 6460 29288
rect 5960 29248 5966 29260
rect 6454 29248 6460 29260
rect 6512 29288 6518 29300
rect 7101 29291 7159 29297
rect 7101 29288 7113 29291
rect 6512 29260 7113 29288
rect 6512 29248 6518 29260
rect 7101 29257 7113 29260
rect 7147 29288 7159 29291
rect 7285 29291 7343 29297
rect 7285 29288 7297 29291
rect 7147 29260 7297 29288
rect 7147 29257 7159 29260
rect 7101 29251 7159 29257
rect 7285 29257 7297 29260
rect 7331 29257 7343 29291
rect 9306 29288 9312 29300
rect 7285 29251 7343 29257
rect 8128 29260 9312 29288
rect 5810 29220 5816 29232
rect 5460 29192 5816 29220
rect 5810 29180 5816 29192
rect 5868 29180 5874 29232
rect 7300 29220 7328 29251
rect 8128 29220 8156 29260
rect 9306 29248 9312 29260
rect 9364 29248 9370 29300
rect 10502 29248 10508 29300
rect 10560 29288 10566 29300
rect 10560 29260 10916 29288
rect 10560 29248 10566 29260
rect 9585 29223 9643 29229
rect 7300 29192 8234 29220
rect 9585 29189 9597 29223
rect 9631 29220 9643 29223
rect 9631 29192 10640 29220
rect 9631 29189 9643 29192
rect 9585 29183 9643 29189
rect 10612 29164 10640 29192
rect 10778 29180 10784 29232
rect 10836 29180 10842 29232
rect 5718 29112 5724 29164
rect 5776 29112 5782 29164
rect 5997 29155 6055 29161
rect 5997 29121 6009 29155
rect 6043 29152 6055 29155
rect 6086 29152 6092 29164
rect 6043 29124 6092 29152
rect 6043 29121 6055 29124
rect 5997 29115 6055 29121
rect 6012 29084 6040 29115
rect 6086 29112 6092 29124
rect 6144 29112 6150 29164
rect 9861 29155 9919 29161
rect 9861 29152 9873 29155
rect 9324 29124 9873 29152
rect 5092 29056 6040 29084
rect 7469 29087 7527 29093
rect 7469 29053 7481 29087
rect 7515 29084 7527 29087
rect 7515 29056 7604 29084
rect 7515 29053 7527 29056
rect 7469 29047 7527 29053
rect 2924 28988 4200 29016
rect 2924 28976 2930 28988
rect 3602 28908 3608 28960
rect 3660 28948 3666 28960
rect 4065 28951 4123 28957
rect 4065 28948 4077 28951
rect 3660 28920 4077 28948
rect 3660 28908 3666 28920
rect 4065 28917 4077 28920
rect 4111 28917 4123 28951
rect 4172 28948 4200 28988
rect 5261 28951 5319 28957
rect 5261 28948 5273 28951
rect 4172 28920 5273 28948
rect 4065 28911 4123 28917
rect 5261 28917 5273 28920
rect 5307 28917 5319 28951
rect 5261 28911 5319 28917
rect 5902 28908 5908 28960
rect 5960 28908 5966 28960
rect 7576 28948 7604 29056
rect 7742 29044 7748 29096
rect 7800 29044 7806 29096
rect 9214 28976 9220 29028
rect 9272 29016 9278 29028
rect 9324 29016 9352 29124
rect 9861 29121 9873 29124
rect 9907 29121 9919 29155
rect 9861 29115 9919 29121
rect 10594 29112 10600 29164
rect 10652 29112 10658 29164
rect 10888 29161 10916 29260
rect 11790 29248 11796 29300
rect 11848 29288 11854 29300
rect 12529 29291 12587 29297
rect 12529 29288 12541 29291
rect 11848 29260 12541 29288
rect 11848 29248 11854 29260
rect 12529 29257 12541 29260
rect 12575 29257 12587 29291
rect 12529 29251 12587 29257
rect 12897 29291 12955 29297
rect 12897 29257 12909 29291
rect 12943 29288 12955 29291
rect 13262 29288 13268 29300
rect 12943 29260 13268 29288
rect 12943 29257 12955 29260
rect 12897 29251 12955 29257
rect 13262 29248 13268 29260
rect 13320 29248 13326 29300
rect 15654 29248 15660 29300
rect 15712 29248 15718 29300
rect 17218 29248 17224 29300
rect 17276 29288 17282 29300
rect 17405 29291 17463 29297
rect 17405 29288 17417 29291
rect 17276 29260 17417 29288
rect 17276 29248 17282 29260
rect 17405 29257 17417 29260
rect 17451 29257 17463 29291
rect 17405 29251 17463 29257
rect 19518 29248 19524 29300
rect 19576 29288 19582 29300
rect 19705 29291 19763 29297
rect 19705 29288 19717 29291
rect 19576 29260 19717 29288
rect 19576 29248 19582 29260
rect 19705 29257 19717 29260
rect 19751 29257 19763 29291
rect 19705 29251 19763 29257
rect 20073 29291 20131 29297
rect 20073 29257 20085 29291
rect 20119 29288 20131 29291
rect 20162 29288 20168 29300
rect 20119 29260 20168 29288
rect 20119 29257 20131 29260
rect 20073 29251 20131 29257
rect 20162 29248 20168 29260
rect 20220 29248 20226 29300
rect 22186 29248 22192 29300
rect 22244 29288 22250 29300
rect 23293 29291 23351 29297
rect 23293 29288 23305 29291
rect 22244 29260 23305 29288
rect 22244 29248 22250 29260
rect 23293 29257 23305 29260
rect 23339 29257 23351 29291
rect 23293 29251 23351 29257
rect 12986 29180 12992 29232
rect 13044 29180 13050 29232
rect 16206 29220 16212 29232
rect 15410 29192 16212 29220
rect 16206 29180 16212 29192
rect 16264 29180 16270 29232
rect 23308 29220 23336 29251
rect 23474 29248 23480 29300
rect 23532 29288 23538 29300
rect 23661 29291 23719 29297
rect 23661 29288 23673 29291
rect 23532 29260 23673 29288
rect 23532 29248 23538 29260
rect 23661 29257 23673 29260
rect 23707 29288 23719 29291
rect 24762 29288 24768 29300
rect 23707 29260 24768 29288
rect 23707 29257 23719 29260
rect 23661 29251 23719 29257
rect 24762 29248 24768 29260
rect 24820 29248 24826 29300
rect 26602 29248 26608 29300
rect 26660 29288 26666 29300
rect 27522 29288 27528 29300
rect 26660 29260 27528 29288
rect 26660 29248 26666 29260
rect 27522 29248 27528 29260
rect 27580 29288 27586 29300
rect 28813 29291 28871 29297
rect 28813 29288 28825 29291
rect 27580 29260 28825 29288
rect 27580 29248 27586 29260
rect 28813 29257 28825 29260
rect 28859 29288 28871 29291
rect 28902 29288 28908 29300
rect 28859 29260 28908 29288
rect 28859 29257 28871 29260
rect 28813 29251 28871 29257
rect 28902 29248 28908 29260
rect 28960 29288 28966 29300
rect 28960 29260 29224 29288
rect 28960 29248 28966 29260
rect 23569 29223 23627 29229
rect 23569 29220 23581 29223
rect 23308 29192 23581 29220
rect 23569 29189 23581 29192
rect 23615 29220 23627 29223
rect 23842 29220 23848 29232
rect 23615 29192 23848 29220
rect 23615 29189 23627 29192
rect 23569 29183 23627 29189
rect 23842 29180 23848 29192
rect 23900 29220 23906 29232
rect 23900 29192 23966 29220
rect 23900 29180 23906 29192
rect 25130 29180 25136 29232
rect 25188 29180 25194 29232
rect 27540 29220 27568 29248
rect 29196 29220 29224 29260
rect 30098 29248 30104 29300
rect 30156 29248 30162 29300
rect 33965 29291 34023 29297
rect 33965 29257 33977 29291
rect 34011 29288 34023 29291
rect 34606 29288 34612 29300
rect 34011 29260 34612 29288
rect 34011 29257 34023 29260
rect 33965 29251 34023 29257
rect 34606 29248 34612 29260
rect 34664 29248 34670 29300
rect 30116 29220 30144 29248
rect 27540 29192 27738 29220
rect 29196 29192 29302 29220
rect 30116 29192 31248 29220
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29121 10747 29155
rect 10689 29115 10747 29121
rect 10873 29155 10931 29161
rect 10873 29121 10885 29155
rect 10919 29121 10931 29155
rect 10873 29115 10931 29121
rect 9674 29044 9680 29096
rect 9732 29044 9738 29096
rect 9766 29044 9772 29096
rect 9824 29084 9830 29096
rect 10704 29084 10732 29115
rect 15746 29112 15752 29164
rect 15804 29152 15810 29164
rect 17037 29155 17095 29161
rect 17037 29152 17049 29155
rect 15804 29124 17049 29152
rect 15804 29112 15810 29124
rect 17037 29121 17049 29124
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 17310 29112 17316 29164
rect 17368 29152 17374 29164
rect 18877 29155 18935 29161
rect 18877 29152 18889 29155
rect 17368 29124 18889 29152
rect 17368 29112 17374 29124
rect 18877 29121 18889 29124
rect 18923 29121 18935 29155
rect 18877 29115 18935 29121
rect 18969 29155 19027 29161
rect 18969 29121 18981 29155
rect 19015 29152 19027 29155
rect 19886 29152 19892 29164
rect 19015 29124 19892 29152
rect 19015 29121 19027 29124
rect 18969 29115 19027 29121
rect 19886 29112 19892 29124
rect 19944 29112 19950 29164
rect 20165 29155 20223 29161
rect 20165 29121 20177 29155
rect 20211 29152 20223 29155
rect 21266 29152 21272 29164
rect 20211 29124 21272 29152
rect 20211 29121 20223 29124
rect 20165 29115 20223 29121
rect 21266 29112 21272 29124
rect 21324 29112 21330 29164
rect 21361 29155 21419 29161
rect 21361 29121 21373 29155
rect 21407 29152 21419 29155
rect 22646 29152 22652 29164
rect 21407 29124 22652 29152
rect 21407 29121 21419 29124
rect 21361 29115 21419 29121
rect 22646 29112 22652 29124
rect 22704 29112 22710 29164
rect 25406 29112 25412 29164
rect 25464 29152 25470 29164
rect 26142 29152 26148 29164
rect 25464 29124 26148 29152
rect 25464 29112 25470 29124
rect 26142 29112 26148 29124
rect 26200 29152 26206 29164
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26200 29124 26985 29152
rect 26200 29112 26206 29124
rect 26973 29121 26985 29124
rect 27019 29121 27031 29155
rect 26973 29115 27031 29121
rect 9824 29056 10732 29084
rect 9824 29044 9830 29056
rect 13170 29044 13176 29096
rect 13228 29044 13234 29096
rect 13909 29087 13967 29093
rect 13909 29053 13921 29087
rect 13955 29084 13967 29087
rect 13955 29056 14044 29084
rect 13955 29053 13967 29056
rect 13909 29047 13967 29053
rect 9272 28988 9352 29016
rect 10045 29019 10103 29025
rect 9272 28976 9278 28988
rect 10045 28985 10057 29019
rect 10091 29016 10103 29019
rect 10226 29016 10232 29028
rect 10091 28988 10232 29016
rect 10091 28985 10103 28988
rect 10045 28979 10103 28985
rect 10226 28976 10232 28988
rect 10284 28976 10290 29028
rect 8202 28948 8208 28960
rect 7576 28920 8208 28948
rect 8202 28908 8208 28920
rect 8260 28908 8266 28960
rect 9582 28908 9588 28960
rect 9640 28908 9646 28960
rect 14016 28948 14044 29056
rect 14182 29044 14188 29096
rect 14240 29044 14246 29096
rect 14642 29044 14648 29096
rect 14700 29084 14706 29096
rect 16761 29087 16819 29093
rect 16761 29084 16773 29087
rect 14700 29056 16773 29084
rect 14700 29044 14706 29056
rect 16761 29053 16773 29056
rect 16807 29053 16819 29087
rect 16761 29047 16819 29053
rect 16776 29016 16804 29047
rect 16850 29044 16856 29096
rect 16908 29084 16914 29096
rect 16945 29087 17003 29093
rect 16945 29084 16957 29087
rect 16908 29056 16957 29084
rect 16908 29044 16914 29056
rect 16945 29053 16957 29056
rect 16991 29053 17003 29087
rect 16945 29047 17003 29053
rect 19153 29087 19211 29093
rect 19153 29053 19165 29087
rect 19199 29084 19211 29087
rect 20254 29084 20260 29096
rect 19199 29056 20260 29084
rect 19199 29053 19211 29056
rect 19153 29047 19211 29053
rect 20254 29044 20260 29056
rect 20312 29044 20318 29096
rect 20898 29044 20904 29096
rect 20956 29084 20962 29096
rect 21450 29084 21456 29096
rect 20956 29056 21456 29084
rect 20956 29044 20962 29056
rect 21450 29044 21456 29056
rect 21508 29044 21514 29096
rect 27246 29044 27252 29096
rect 27304 29044 27310 29096
rect 30466 29044 30472 29096
rect 30524 29044 30530 29096
rect 30745 29087 30803 29093
rect 30745 29053 30757 29087
rect 30791 29053 30803 29087
rect 30745 29047 30803 29053
rect 17954 29016 17960 29028
rect 16776 28988 17960 29016
rect 17954 28976 17960 28988
rect 18012 29016 18018 29028
rect 18414 29016 18420 29028
rect 18012 28988 18420 29016
rect 18012 28976 18018 28988
rect 18414 28976 18420 28988
rect 18472 28976 18478 29028
rect 30760 29016 30788 29047
rect 30834 29044 30840 29096
rect 30892 29044 30898 29096
rect 31220 29084 31248 29192
rect 32490 29180 32496 29232
rect 32548 29180 32554 29232
rect 33502 29180 33508 29232
rect 33560 29180 33566 29232
rect 31297 29155 31355 29161
rect 31297 29121 31309 29155
rect 31343 29152 31355 29155
rect 31386 29152 31392 29164
rect 31343 29124 31392 29152
rect 31343 29121 31355 29124
rect 31297 29115 31355 29121
rect 31386 29112 31392 29124
rect 31444 29112 31450 29164
rect 31481 29155 31539 29161
rect 31481 29121 31493 29155
rect 31527 29152 31539 29155
rect 31938 29152 31944 29164
rect 31527 29124 31944 29152
rect 31527 29121 31539 29124
rect 31481 29115 31539 29121
rect 31938 29112 31944 29124
rect 31996 29112 32002 29164
rect 31573 29087 31631 29093
rect 31573 29084 31585 29087
rect 31220 29056 31585 29084
rect 31573 29053 31585 29056
rect 31619 29053 31631 29087
rect 31573 29047 31631 29053
rect 32217 29087 32275 29093
rect 32217 29053 32229 29087
rect 32263 29053 32275 29087
rect 32217 29047 32275 29053
rect 31846 29016 31852 29028
rect 30760 28988 31852 29016
rect 31846 28976 31852 28988
rect 31904 29016 31910 29028
rect 32232 29016 32260 29047
rect 33134 29044 33140 29096
rect 33192 29084 33198 29096
rect 33520 29084 33548 29180
rect 33192 29056 33548 29084
rect 33192 29044 33198 29056
rect 31904 28988 32260 29016
rect 31904 28976 31910 28988
rect 14734 28948 14740 28960
rect 14016 28920 14740 28948
rect 14734 28908 14740 28920
rect 14792 28908 14798 28960
rect 18509 28951 18567 28957
rect 18509 28917 18521 28951
rect 18555 28948 18567 28951
rect 18782 28948 18788 28960
rect 18555 28920 18788 28948
rect 18555 28917 18567 28920
rect 18509 28911 18567 28917
rect 18782 28908 18788 28920
rect 18840 28908 18846 28960
rect 20714 28908 20720 28960
rect 20772 28948 20778 28960
rect 20901 28951 20959 28957
rect 20901 28948 20913 28951
rect 20772 28920 20913 28948
rect 20772 28908 20778 28920
rect 20901 28917 20913 28920
rect 20947 28917 20959 28951
rect 20901 28911 20959 28917
rect 27614 28908 27620 28960
rect 27672 28948 27678 28960
rect 28721 28951 28779 28957
rect 28721 28948 28733 28951
rect 27672 28920 28733 28948
rect 27672 28908 27678 28920
rect 28721 28917 28733 28920
rect 28767 28917 28779 28951
rect 28721 28911 28779 28917
rect 28994 28908 29000 28960
rect 29052 28908 29058 28960
rect 1104 28858 37076 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 37076 28858
rect 1104 28784 37076 28806
rect 1670 28704 1676 28756
rect 1728 28744 1734 28756
rect 2041 28747 2099 28753
rect 2041 28744 2053 28747
rect 1728 28716 2053 28744
rect 1728 28704 1734 28716
rect 2041 28713 2053 28716
rect 2087 28713 2099 28747
rect 4062 28744 4068 28756
rect 2041 28707 2099 28713
rect 3896 28716 4068 28744
rect 2685 28611 2743 28617
rect 2685 28577 2697 28611
rect 2731 28608 2743 28611
rect 2731 28580 3556 28608
rect 2731 28577 2743 28580
rect 2685 28571 2743 28577
rect 2409 28543 2467 28549
rect 2409 28509 2421 28543
rect 2455 28540 2467 28543
rect 2866 28540 2872 28552
rect 2455 28512 2872 28540
rect 2455 28509 2467 28512
rect 2409 28503 2467 28509
rect 2866 28500 2872 28512
rect 2924 28500 2930 28552
rect 3053 28543 3111 28549
rect 3053 28509 3065 28543
rect 3099 28509 3111 28543
rect 3528 28540 3556 28580
rect 3602 28568 3608 28620
rect 3660 28608 3666 28620
rect 3896 28617 3924 28716
rect 4062 28704 4068 28716
rect 4120 28744 4126 28756
rect 4617 28747 4675 28753
rect 4617 28744 4629 28747
rect 4120 28716 4629 28744
rect 4120 28704 4126 28716
rect 4617 28713 4629 28716
rect 4663 28713 4675 28747
rect 4617 28707 4675 28713
rect 5994 28704 6000 28756
rect 6052 28744 6058 28756
rect 6730 28744 6736 28756
rect 6052 28716 6736 28744
rect 6052 28704 6058 28716
rect 6730 28704 6736 28716
rect 6788 28704 6794 28756
rect 7742 28704 7748 28756
rect 7800 28744 7806 28756
rect 7929 28747 7987 28753
rect 7929 28744 7941 28747
rect 7800 28716 7941 28744
rect 7800 28704 7806 28716
rect 7929 28713 7941 28716
rect 7975 28713 7987 28747
rect 7929 28707 7987 28713
rect 8294 28704 8300 28756
rect 8352 28704 8358 28756
rect 14182 28704 14188 28756
rect 14240 28744 14246 28756
rect 14829 28747 14887 28753
rect 14829 28744 14841 28747
rect 14240 28716 14841 28744
rect 14240 28704 14246 28716
rect 14829 28713 14841 28716
rect 14875 28713 14887 28747
rect 14829 28707 14887 28713
rect 17310 28704 17316 28756
rect 17368 28704 17374 28756
rect 21266 28704 21272 28756
rect 21324 28744 21330 28756
rect 22189 28747 22247 28753
rect 22189 28744 22201 28747
rect 21324 28716 22201 28744
rect 21324 28704 21330 28716
rect 22189 28713 22201 28716
rect 22235 28713 22247 28747
rect 22189 28707 22247 28713
rect 23017 28747 23075 28753
rect 23017 28713 23029 28747
rect 23063 28744 23075 28747
rect 23290 28744 23296 28756
rect 23063 28716 23296 28744
rect 23063 28713 23075 28716
rect 23017 28707 23075 28713
rect 23290 28704 23296 28716
rect 23348 28704 23354 28756
rect 23658 28704 23664 28756
rect 23716 28744 23722 28756
rect 23845 28747 23903 28753
rect 23845 28744 23857 28747
rect 23716 28716 23857 28744
rect 23716 28704 23722 28716
rect 23845 28713 23857 28716
rect 23891 28713 23903 28747
rect 23845 28707 23903 28713
rect 24688 28716 26234 28744
rect 4341 28679 4399 28685
rect 4341 28645 4353 28679
rect 4387 28676 4399 28679
rect 4798 28676 4804 28688
rect 4387 28648 4804 28676
rect 4387 28645 4399 28648
rect 4341 28639 4399 28645
rect 4798 28636 4804 28648
rect 4856 28636 4862 28688
rect 3881 28611 3939 28617
rect 3881 28608 3893 28611
rect 3660 28580 3893 28608
rect 3660 28568 3666 28580
rect 3881 28577 3893 28580
rect 3927 28577 3939 28611
rect 3881 28571 3939 28577
rect 3970 28568 3976 28620
rect 4028 28608 4034 28620
rect 4028 28580 4752 28608
rect 4028 28568 4034 28580
rect 3988 28540 4016 28568
rect 3528 28512 4016 28540
rect 4065 28543 4123 28549
rect 3053 28503 3111 28509
rect 4065 28509 4077 28543
rect 4111 28509 4123 28543
rect 4065 28503 4123 28509
rect 4157 28543 4215 28549
rect 4157 28509 4169 28543
rect 4203 28540 4215 28543
rect 4614 28540 4620 28552
rect 4203 28512 4620 28540
rect 4203 28509 4215 28512
rect 4157 28503 4215 28509
rect 3068 28472 3096 28503
rect 3510 28472 3516 28484
rect 3068 28444 3516 28472
rect 3510 28432 3516 28444
rect 3568 28432 3574 28484
rect 3694 28432 3700 28484
rect 3752 28472 3758 28484
rect 4080 28472 4108 28503
rect 4614 28500 4620 28512
rect 4672 28500 4678 28552
rect 3752 28444 4108 28472
rect 4433 28475 4491 28481
rect 3752 28432 3758 28444
rect 4433 28441 4445 28475
rect 4479 28472 4491 28475
rect 4724 28472 4752 28580
rect 13170 28568 13176 28620
rect 13228 28568 13234 28620
rect 15473 28611 15531 28617
rect 15473 28577 15485 28611
rect 15519 28608 15531 28611
rect 16390 28608 16396 28620
rect 15519 28580 16396 28608
rect 15519 28577 15531 28580
rect 15473 28571 15531 28577
rect 16390 28568 16396 28580
rect 16448 28568 16454 28620
rect 18782 28568 18788 28620
rect 18840 28568 18846 28620
rect 19061 28611 19119 28617
rect 19061 28577 19073 28611
rect 19107 28608 19119 28611
rect 19242 28608 19248 28620
rect 19107 28580 19248 28608
rect 19107 28577 19119 28580
rect 19061 28571 19119 28577
rect 19242 28568 19248 28580
rect 19300 28568 19306 28620
rect 19334 28568 19340 28620
rect 19392 28608 19398 28620
rect 20073 28611 20131 28617
rect 20073 28608 20085 28611
rect 19392 28580 20085 28608
rect 19392 28568 19398 28580
rect 20073 28577 20085 28580
rect 20119 28577 20131 28611
rect 20073 28571 20131 28577
rect 20714 28568 20720 28620
rect 20772 28568 20778 28620
rect 21450 28568 21456 28620
rect 21508 28608 21514 28620
rect 22373 28611 22431 28617
rect 22373 28608 22385 28611
rect 21508 28580 22385 28608
rect 21508 28568 21514 28580
rect 22373 28577 22385 28580
rect 22419 28577 22431 28611
rect 22373 28571 22431 28577
rect 22554 28568 22560 28620
rect 22612 28568 22618 28620
rect 23293 28611 23351 28617
rect 23293 28577 23305 28611
rect 23339 28608 23351 28611
rect 24688 28608 24716 28716
rect 26206 28676 26234 28716
rect 27246 28704 27252 28756
rect 27304 28704 27310 28756
rect 29365 28747 29423 28753
rect 29365 28713 29377 28747
rect 29411 28744 29423 28747
rect 30466 28744 30472 28756
rect 29411 28716 30472 28744
rect 29411 28713 29423 28716
rect 29365 28707 29423 28713
rect 30466 28704 30472 28716
rect 30524 28704 30530 28756
rect 26510 28676 26516 28688
rect 26206 28648 26516 28676
rect 26510 28636 26516 28648
rect 26568 28676 26574 28688
rect 29086 28676 29092 28688
rect 26568 28648 29092 28676
rect 26568 28636 26574 28648
rect 23339 28580 24716 28608
rect 23339 28577 23351 28580
rect 23293 28571 23351 28577
rect 25866 28568 25872 28620
rect 25924 28568 25930 28620
rect 26142 28568 26148 28620
rect 26200 28568 26206 28620
rect 27893 28611 27951 28617
rect 27893 28577 27905 28611
rect 27939 28608 27951 28611
rect 27982 28608 27988 28620
rect 27939 28580 27988 28608
rect 27939 28577 27951 28580
rect 27893 28571 27951 28577
rect 27982 28568 27988 28580
rect 28040 28568 28046 28620
rect 28828 28617 28856 28648
rect 29086 28636 29092 28648
rect 29144 28636 29150 28688
rect 30098 28636 30104 28688
rect 30156 28636 30162 28688
rect 28813 28611 28871 28617
rect 28813 28577 28825 28611
rect 28859 28577 28871 28611
rect 28813 28571 28871 28577
rect 28905 28611 28963 28617
rect 28905 28577 28917 28611
rect 28951 28608 28963 28611
rect 29270 28608 29276 28620
rect 28951 28580 29276 28608
rect 28951 28577 28963 28580
rect 28905 28571 28963 28577
rect 29270 28568 29276 28580
rect 29328 28608 29334 28620
rect 29914 28608 29920 28620
rect 29328 28580 29920 28608
rect 29328 28568 29334 28580
rect 29914 28568 29920 28580
rect 29972 28568 29978 28620
rect 30834 28568 30840 28620
rect 30892 28608 30898 28620
rect 31573 28611 31631 28617
rect 31573 28608 31585 28611
rect 30892 28580 31585 28608
rect 30892 28568 30898 28580
rect 31573 28577 31585 28580
rect 31619 28577 31631 28611
rect 31573 28571 31631 28577
rect 33410 28568 33416 28620
rect 33468 28568 33474 28620
rect 8110 28500 8116 28552
rect 8168 28500 8174 28552
rect 8389 28543 8447 28549
rect 8389 28509 8401 28543
rect 8435 28540 8447 28543
rect 8754 28540 8760 28552
rect 8435 28512 8760 28540
rect 8435 28509 8447 28512
rect 8389 28503 8447 28509
rect 8754 28500 8760 28512
rect 8812 28500 8818 28552
rect 13081 28543 13139 28549
rect 13081 28509 13093 28543
rect 13127 28540 13139 28543
rect 13262 28540 13268 28552
rect 13127 28512 13268 28540
rect 13127 28509 13139 28512
rect 13081 28503 13139 28509
rect 13262 28500 13268 28512
rect 13320 28500 13326 28552
rect 15197 28543 15255 28549
rect 15197 28509 15209 28543
rect 15243 28540 15255 28543
rect 15654 28540 15660 28552
rect 15243 28512 15660 28540
rect 15243 28509 15255 28512
rect 15197 28503 15255 28509
rect 15654 28500 15660 28512
rect 15712 28500 15718 28552
rect 19260 28540 19288 28568
rect 20441 28543 20499 28549
rect 20441 28540 20453 28543
rect 19260 28512 20453 28540
rect 20441 28509 20453 28512
rect 20487 28509 20499 28543
rect 20441 28503 20499 28509
rect 22646 28500 22652 28552
rect 22704 28500 22710 28552
rect 23385 28543 23443 28549
rect 23385 28509 23397 28543
rect 23431 28540 23443 28543
rect 23474 28540 23480 28552
rect 23431 28512 23480 28540
rect 23431 28509 23443 28512
rect 23385 28503 23443 28509
rect 23474 28500 23480 28512
rect 23532 28500 23538 28552
rect 27614 28500 27620 28552
rect 27672 28500 27678 28552
rect 27709 28543 27767 28549
rect 27709 28509 27721 28543
rect 27755 28540 27767 28543
rect 28994 28540 29000 28552
rect 27755 28512 29000 28540
rect 27755 28509 27767 28512
rect 27709 28503 27767 28509
rect 28994 28500 29000 28512
rect 29052 28500 29058 28552
rect 31846 28500 31852 28552
rect 31904 28500 31910 28552
rect 33137 28543 33195 28549
rect 33137 28509 33149 28543
rect 33183 28509 33195 28543
rect 33137 28503 33195 28509
rect 33321 28543 33379 28549
rect 33321 28509 33333 28543
rect 33367 28540 33379 28543
rect 33962 28540 33968 28552
rect 33367 28512 33968 28540
rect 33367 28509 33379 28512
rect 33321 28503 33379 28509
rect 4479 28444 4752 28472
rect 4479 28441 4491 28444
rect 4433 28435 4491 28441
rect 5718 28432 5724 28484
rect 5776 28472 5782 28484
rect 5965 28475 6023 28481
rect 5965 28472 5977 28475
rect 5776 28444 5977 28472
rect 5776 28432 5782 28444
rect 5965 28441 5977 28444
rect 6011 28441 6023 28475
rect 5965 28435 6023 28441
rect 6086 28432 6092 28484
rect 6144 28472 6150 28484
rect 6181 28475 6239 28481
rect 6181 28472 6193 28475
rect 6144 28444 6193 28472
rect 6144 28432 6150 28444
rect 6181 28441 6193 28444
rect 6227 28441 6239 28475
rect 6181 28435 6239 28441
rect 15289 28475 15347 28481
rect 15289 28441 15301 28475
rect 15335 28472 15347 28475
rect 15746 28472 15752 28484
rect 15335 28444 15752 28472
rect 15335 28441 15347 28444
rect 15289 28435 15347 28441
rect 15746 28432 15752 28444
rect 15804 28432 15810 28484
rect 18322 28432 18328 28484
rect 18380 28432 18386 28484
rect 19886 28432 19892 28484
rect 19944 28432 19950 28484
rect 19981 28475 20039 28481
rect 19981 28441 19993 28475
rect 20027 28472 20039 28475
rect 20162 28472 20168 28484
rect 20027 28444 20168 28472
rect 20027 28441 20039 28444
rect 19981 28435 20039 28441
rect 20162 28432 20168 28444
rect 20220 28432 20226 28484
rect 20806 28432 20812 28484
rect 20864 28472 20870 28484
rect 20864 28444 21206 28472
rect 20864 28432 20870 28444
rect 23842 28432 23848 28484
rect 23900 28472 23906 28484
rect 23900 28444 24702 28472
rect 23900 28432 23906 28444
rect 30926 28432 30932 28484
rect 30984 28432 30990 28484
rect 32674 28432 32680 28484
rect 32732 28432 32738 28484
rect 33152 28472 33180 28503
rect 33962 28500 33968 28512
rect 34020 28500 34026 28552
rect 33778 28472 33784 28484
rect 33152 28444 33784 28472
rect 33778 28432 33784 28444
rect 33836 28472 33842 28484
rect 35342 28472 35348 28484
rect 33836 28444 35348 28472
rect 33836 28432 33842 28444
rect 35342 28432 35348 28444
rect 35400 28432 35406 28484
rect 2222 28364 2228 28416
rect 2280 28404 2286 28416
rect 2501 28407 2559 28413
rect 2501 28404 2513 28407
rect 2280 28376 2513 28404
rect 2280 28364 2286 28376
rect 2501 28373 2513 28376
rect 2547 28404 2559 28407
rect 2961 28407 3019 28413
rect 2961 28404 2973 28407
rect 2547 28376 2973 28404
rect 2547 28373 2559 28376
rect 2501 28367 2559 28373
rect 2961 28373 2973 28376
rect 3007 28373 3019 28407
rect 2961 28367 3019 28373
rect 4522 28364 4528 28416
rect 4580 28404 4586 28416
rect 4633 28407 4691 28413
rect 4633 28404 4645 28407
rect 4580 28376 4645 28404
rect 4580 28364 4586 28376
rect 4633 28373 4645 28376
rect 4679 28373 4691 28407
rect 4633 28367 4691 28373
rect 4801 28407 4859 28413
rect 4801 28373 4813 28407
rect 4847 28404 4859 28407
rect 5350 28404 5356 28416
rect 4847 28376 5356 28404
rect 4847 28373 4859 28376
rect 4801 28367 4859 28373
rect 5350 28364 5356 28376
rect 5408 28364 5414 28416
rect 5810 28364 5816 28416
rect 5868 28364 5874 28416
rect 11974 28364 11980 28416
rect 12032 28404 12038 28416
rect 12621 28407 12679 28413
rect 12621 28404 12633 28407
rect 12032 28376 12633 28404
rect 12032 28364 12038 28376
rect 12621 28373 12633 28376
rect 12667 28373 12679 28407
rect 12621 28367 12679 28373
rect 12989 28407 13047 28413
rect 12989 28373 13001 28407
rect 13035 28404 13047 28407
rect 13446 28404 13452 28416
rect 13035 28376 13452 28404
rect 13035 28373 13047 28376
rect 12989 28367 13047 28373
rect 13446 28364 13452 28376
rect 13504 28364 13510 28416
rect 19518 28364 19524 28416
rect 19576 28364 19582 28416
rect 22554 28364 22560 28416
rect 22612 28404 22618 28416
rect 23477 28407 23535 28413
rect 23477 28404 23489 28407
rect 22612 28376 23489 28404
rect 22612 28364 22618 28376
rect 23477 28373 23489 28376
rect 23523 28373 23535 28407
rect 23477 28367 23535 28373
rect 24397 28407 24455 28413
rect 24397 28373 24409 28407
rect 24443 28404 24455 28407
rect 25038 28404 25044 28416
rect 24443 28376 25044 28404
rect 24443 28373 24455 28376
rect 24397 28367 24455 28373
rect 25038 28364 25044 28376
rect 25096 28364 25102 28416
rect 1104 28314 37076 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 37076 28314
rect 1104 28240 37076 28262
rect 2866 28160 2872 28212
rect 2924 28200 2930 28212
rect 3053 28203 3111 28209
rect 3053 28200 3065 28203
rect 2924 28172 3065 28200
rect 2924 28160 2930 28172
rect 3053 28169 3065 28172
rect 3099 28169 3111 28203
rect 3053 28163 3111 28169
rect 5629 28203 5687 28209
rect 5629 28169 5641 28203
rect 5675 28200 5687 28203
rect 5902 28200 5908 28212
rect 5675 28172 5908 28200
rect 5675 28169 5687 28172
rect 5629 28163 5687 28169
rect 5902 28160 5908 28172
rect 5960 28160 5966 28212
rect 6086 28160 6092 28212
rect 6144 28200 6150 28212
rect 16485 28203 16543 28209
rect 6144 28172 6776 28200
rect 6144 28160 6150 28172
rect 3205 28135 3263 28141
rect 3205 28132 3217 28135
rect 2700 28104 3217 28132
rect 2222 28024 2228 28076
rect 2280 28024 2286 28076
rect 2700 28073 2728 28104
rect 3205 28101 3217 28104
rect 3251 28132 3263 28135
rect 3251 28104 3372 28132
rect 3251 28101 3263 28104
rect 3205 28095 3263 28101
rect 2685 28067 2743 28073
rect 2685 28033 2697 28067
rect 2731 28033 2743 28067
rect 2685 28027 2743 28033
rect 2869 28067 2927 28073
rect 2869 28033 2881 28067
rect 2915 28033 2927 28067
rect 2869 28027 2927 28033
rect 2961 28067 3019 28073
rect 2961 28033 2973 28067
rect 3007 28064 3019 28067
rect 3344 28064 3372 28104
rect 3418 28092 3424 28144
rect 3476 28092 3482 28144
rect 3694 28092 3700 28144
rect 3752 28132 3758 28144
rect 5258 28132 5264 28144
rect 3752 28104 5264 28132
rect 3752 28092 3758 28104
rect 5258 28092 5264 28104
rect 5316 28092 5322 28144
rect 5350 28092 5356 28144
rect 5408 28132 5414 28144
rect 5461 28135 5519 28141
rect 5461 28132 5473 28135
rect 5408 28104 5473 28132
rect 5408 28092 5414 28104
rect 5461 28101 5473 28104
rect 5507 28101 5519 28135
rect 5461 28095 5519 28101
rect 5718 28092 5724 28144
rect 5776 28092 5782 28144
rect 5920 28132 5948 28160
rect 5920 28104 6592 28132
rect 3602 28064 3608 28076
rect 3007 28036 3188 28064
rect 3344 28036 3608 28064
rect 3007 28033 3019 28036
rect 2961 28027 3019 28033
rect 2409 27999 2467 28005
rect 2409 27965 2421 27999
rect 2455 27996 2467 27999
rect 2501 27999 2559 28005
rect 2501 27996 2513 27999
rect 2455 27968 2513 27996
rect 2455 27965 2467 27968
rect 2409 27959 2467 27965
rect 2501 27965 2513 27968
rect 2547 27965 2559 27999
rect 2884 27996 2912 28027
rect 3050 27996 3056 28008
rect 2884 27968 3056 27996
rect 2501 27959 2559 27965
rect 3050 27956 3056 27968
rect 3108 27956 3114 28008
rect 3160 27872 3188 28036
rect 3602 28024 3608 28036
rect 3660 28064 3666 28076
rect 3881 28067 3939 28073
rect 3881 28064 3893 28067
rect 3660 28036 3893 28064
rect 3660 28024 3666 28036
rect 3881 28033 3893 28036
rect 3927 28033 3939 28067
rect 3881 28027 3939 28033
rect 3970 28024 3976 28076
rect 4028 28024 4034 28076
rect 4062 28024 4068 28076
rect 4120 28064 4126 28076
rect 4157 28067 4215 28073
rect 4157 28064 4169 28067
rect 4120 28036 4169 28064
rect 4120 28024 4126 28036
rect 4157 28033 4169 28036
rect 4203 28033 4215 28067
rect 4157 28027 4215 28033
rect 4522 28024 4528 28076
rect 4580 28064 4586 28076
rect 6564 28073 6592 28104
rect 6748 28073 6776 28172
rect 16485 28169 16497 28203
rect 16531 28200 16543 28203
rect 16850 28200 16856 28212
rect 16531 28172 16856 28200
rect 16531 28169 16543 28172
rect 16485 28163 16543 28169
rect 16850 28160 16856 28172
rect 16908 28160 16914 28212
rect 28169 28203 28227 28209
rect 28169 28169 28181 28203
rect 28215 28200 28227 28203
rect 29270 28200 29276 28212
rect 28215 28172 29276 28200
rect 28215 28169 28227 28172
rect 28169 28163 28227 28169
rect 29270 28160 29276 28172
rect 29328 28160 29334 28212
rect 33410 28160 33416 28212
rect 33468 28200 33474 28212
rect 33873 28203 33931 28209
rect 33873 28200 33885 28203
rect 33468 28172 33885 28200
rect 33468 28160 33474 28172
rect 33873 28169 33885 28172
rect 33919 28169 33931 28203
rect 33873 28163 33931 28169
rect 10258 28104 11284 28132
rect 5997 28067 6055 28073
rect 5997 28064 6009 28067
rect 4580 28036 6009 28064
rect 4580 28024 4586 28036
rect 5997 28033 6009 28036
rect 6043 28033 6055 28067
rect 5997 28027 6055 28033
rect 6549 28067 6607 28073
rect 6549 28033 6561 28067
rect 6595 28033 6607 28067
rect 6549 28027 6607 28033
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28033 6791 28067
rect 10781 28067 10839 28073
rect 10781 28064 10793 28067
rect 6733 28027 6791 28033
rect 10244 28036 10793 28064
rect 5902 27956 5908 28008
rect 5960 27996 5966 28008
rect 6641 27999 6699 28005
rect 6641 27996 6653 27999
rect 5960 27968 6653 27996
rect 5960 27956 5966 27968
rect 6641 27965 6653 27968
rect 6687 27965 6699 27999
rect 6641 27959 6699 27965
rect 6822 27956 6828 28008
rect 6880 27956 6886 28008
rect 8202 27956 8208 28008
rect 8260 27996 8266 28008
rect 8757 27999 8815 28005
rect 8757 27996 8769 27999
rect 8260 27968 8769 27996
rect 8260 27956 8266 27968
rect 8757 27965 8769 27968
rect 8803 27965 8815 27999
rect 8757 27959 8815 27965
rect 9030 27956 9036 28008
rect 9088 27956 9094 28008
rect 9122 27956 9128 28008
rect 9180 27996 9186 28008
rect 10244 27996 10272 28036
rect 10781 28033 10793 28036
rect 10827 28033 10839 28067
rect 10781 28027 10839 28033
rect 10965 27999 11023 28005
rect 10965 27996 10977 27999
rect 9180 27968 10272 27996
rect 10796 27968 10977 27996
rect 9180 27956 9186 27968
rect 4341 27931 4399 27937
rect 4341 27897 4353 27931
rect 4387 27928 4399 27931
rect 5626 27928 5632 27940
rect 4387 27900 5632 27928
rect 4387 27897 4399 27900
rect 4341 27891 4399 27897
rect 5626 27888 5632 27900
rect 5684 27888 5690 27940
rect 5994 27888 6000 27940
rect 6052 27928 6058 27940
rect 6365 27931 6423 27937
rect 6365 27928 6377 27931
rect 6052 27900 6377 27928
rect 6052 27888 6058 27900
rect 6365 27897 6377 27900
rect 6411 27897 6423 27931
rect 6365 27891 6423 27897
rect 10042 27888 10048 27940
rect 10100 27928 10106 27940
rect 10597 27931 10655 27937
rect 10597 27928 10609 27931
rect 10100 27900 10609 27928
rect 10100 27888 10106 27900
rect 10597 27897 10609 27900
rect 10643 27897 10655 27931
rect 10597 27891 10655 27897
rect 10796 27872 10824 27968
rect 10965 27965 10977 27968
rect 11011 27965 11023 27999
rect 11256 27996 11284 28104
rect 11974 28092 11980 28144
rect 12032 28092 12038 28144
rect 13722 28132 13728 28144
rect 13202 28118 13728 28132
rect 13188 28104 13728 28118
rect 11514 28024 11520 28076
rect 11572 28064 11578 28076
rect 11698 28064 11704 28076
rect 11572 28036 11704 28064
rect 11572 28024 11578 28036
rect 11698 28024 11704 28036
rect 11756 28024 11762 28076
rect 12434 27996 12440 28008
rect 11256 27968 12440 27996
rect 10965 27959 11023 27965
rect 12434 27956 12440 27968
rect 12492 27996 12498 28008
rect 13188 27996 13216 28104
rect 13722 28092 13728 28104
rect 13780 28092 13786 28144
rect 18230 28132 18236 28144
rect 17710 28104 18236 28132
rect 18230 28092 18236 28104
rect 18288 28092 18294 28144
rect 28902 28092 28908 28144
rect 28960 28092 28966 28144
rect 29546 28092 29552 28144
rect 29604 28132 29610 28144
rect 29641 28135 29699 28141
rect 29641 28132 29653 28135
rect 29604 28104 29653 28132
rect 29604 28092 29610 28104
rect 29641 28101 29653 28104
rect 29687 28101 29699 28135
rect 29641 28095 29699 28101
rect 32401 28135 32459 28141
rect 32401 28101 32413 28135
rect 32447 28132 32459 28135
rect 32674 28132 32680 28144
rect 32447 28104 32680 28132
rect 32447 28101 32459 28104
rect 32401 28095 32459 28101
rect 32674 28092 32680 28104
rect 32732 28092 32738 28144
rect 33134 28092 33140 28144
rect 33192 28092 33198 28144
rect 16114 28024 16120 28076
rect 16172 28024 16178 28076
rect 21361 28067 21419 28073
rect 21361 28033 21373 28067
rect 21407 28064 21419 28067
rect 22646 28064 22652 28076
rect 21407 28036 22652 28064
rect 21407 28033 21419 28036
rect 21361 28027 21419 28033
rect 22646 28024 22652 28036
rect 22704 28024 22710 28076
rect 25130 28024 25136 28076
rect 25188 28064 25194 28076
rect 26053 28067 26111 28073
rect 26053 28064 26065 28067
rect 25188 28036 26065 28064
rect 25188 28024 25194 28036
rect 26053 28033 26065 28036
rect 26099 28033 26111 28067
rect 26053 28027 26111 28033
rect 30006 28024 30012 28076
rect 30064 28064 30070 28076
rect 30469 28067 30527 28073
rect 30469 28064 30481 28067
rect 30064 28036 30481 28064
rect 30064 28024 30070 28036
rect 30469 28033 30481 28036
rect 30515 28033 30527 28067
rect 30469 28027 30527 28033
rect 30926 28024 30932 28076
rect 30984 28024 30990 28076
rect 12492 27968 13216 27996
rect 12492 27956 12498 27968
rect 14734 27956 14740 28008
rect 14792 27956 14798 28008
rect 15013 27999 15071 28005
rect 15013 27965 15025 27999
rect 15059 27996 15071 27999
rect 16298 27996 16304 28008
rect 15059 27968 16304 27996
rect 15059 27965 15071 27968
rect 15013 27959 15071 27965
rect 16298 27956 16304 27968
rect 16356 27956 16362 28008
rect 18138 27956 18144 28008
rect 18196 27956 18202 28008
rect 18417 27999 18475 28005
rect 18417 27965 18429 27999
rect 18463 27996 18475 27999
rect 19242 27996 19248 28008
rect 18463 27968 19248 27996
rect 18463 27965 18475 27968
rect 18417 27959 18475 27965
rect 19242 27956 19248 27968
rect 19300 27956 19306 28008
rect 19334 27956 19340 28008
rect 19392 27996 19398 28008
rect 19613 27999 19671 28005
rect 19613 27996 19625 27999
rect 19392 27968 19625 27996
rect 19392 27956 19398 27968
rect 19613 27965 19625 27968
rect 19659 27965 19671 27999
rect 19613 27959 19671 27965
rect 25958 27956 25964 28008
rect 26016 27996 26022 28008
rect 26145 27999 26203 28005
rect 26145 27996 26157 27999
rect 26016 27968 26157 27996
rect 26016 27956 26022 27968
rect 26145 27965 26157 27968
rect 26191 27965 26203 27999
rect 26145 27959 26203 27965
rect 26237 27999 26295 28005
rect 26237 27965 26249 27999
rect 26283 27965 26295 27999
rect 26237 27959 26295 27965
rect 29917 27999 29975 28005
rect 29917 27965 29929 27999
rect 29963 27996 29975 27999
rect 30098 27996 30104 28008
rect 29963 27968 30104 27996
rect 29963 27965 29975 27968
rect 29917 27959 29975 27965
rect 25498 27888 25504 27940
rect 25556 27928 25562 27940
rect 26252 27928 26280 27959
rect 30098 27956 30104 27968
rect 30156 27956 30162 28008
rect 30285 27999 30343 28005
rect 30285 27965 30297 27999
rect 30331 27965 30343 27999
rect 30285 27959 30343 27965
rect 30377 27999 30435 28005
rect 30377 27965 30389 27999
rect 30423 27996 30435 27999
rect 31018 27996 31024 28008
rect 30423 27968 31024 27996
rect 30423 27965 30435 27968
rect 30377 27959 30435 27965
rect 25556 27900 26280 27928
rect 30300 27928 30328 27959
rect 31018 27956 31024 27968
rect 31076 27956 31082 28008
rect 31294 27956 31300 28008
rect 31352 27996 31358 28008
rect 31665 27999 31723 28005
rect 31665 27996 31677 27999
rect 31352 27968 31677 27996
rect 31352 27956 31358 27968
rect 31665 27965 31677 27968
rect 31711 27996 31723 27999
rect 31846 27996 31852 28008
rect 31711 27968 31852 27996
rect 31711 27965 31723 27968
rect 31665 27959 31723 27965
rect 31846 27956 31852 27968
rect 31904 27996 31910 28008
rect 32125 27999 32183 28005
rect 32125 27996 32137 27999
rect 31904 27968 32137 27996
rect 31904 27956 31910 27968
rect 32125 27965 32137 27968
rect 32171 27965 32183 27999
rect 32125 27959 32183 27965
rect 30466 27928 30472 27940
rect 30300 27900 30472 27928
rect 25556 27888 25562 27900
rect 30466 27888 30472 27900
rect 30524 27928 30530 27940
rect 31754 27928 31760 27940
rect 30524 27900 31760 27928
rect 30524 27888 30530 27900
rect 31754 27888 31760 27900
rect 31812 27888 31818 27940
rect 2041 27863 2099 27869
rect 2041 27829 2053 27863
rect 2087 27860 2099 27863
rect 2130 27860 2136 27872
rect 2087 27832 2136 27860
rect 2087 27829 2099 27832
rect 2041 27823 2099 27829
rect 2130 27820 2136 27832
rect 2188 27820 2194 27872
rect 3142 27820 3148 27872
rect 3200 27860 3206 27872
rect 3237 27863 3295 27869
rect 3237 27860 3249 27863
rect 3200 27832 3249 27860
rect 3200 27820 3206 27832
rect 3237 27829 3249 27832
rect 3283 27829 3295 27863
rect 3237 27823 3295 27829
rect 4614 27820 4620 27872
rect 4672 27860 4678 27872
rect 5442 27860 5448 27872
rect 4672 27832 5448 27860
rect 4672 27820 4678 27832
rect 5442 27820 5448 27832
rect 5500 27820 5506 27872
rect 5905 27863 5963 27869
rect 5905 27829 5917 27863
rect 5951 27860 5963 27863
rect 6086 27860 6092 27872
rect 5951 27832 6092 27860
rect 5951 27829 5963 27832
rect 5905 27823 5963 27829
rect 6086 27820 6092 27832
rect 6144 27820 6150 27872
rect 6181 27863 6239 27869
rect 6181 27829 6193 27863
rect 6227 27860 6239 27863
rect 6270 27860 6276 27872
rect 6227 27832 6276 27860
rect 6227 27829 6239 27832
rect 6181 27823 6239 27829
rect 6270 27820 6276 27832
rect 6328 27820 6334 27872
rect 10505 27863 10563 27869
rect 10505 27829 10517 27863
rect 10551 27860 10563 27863
rect 10778 27860 10784 27872
rect 10551 27832 10784 27860
rect 10551 27829 10563 27832
rect 10505 27823 10563 27829
rect 10778 27820 10784 27832
rect 10836 27820 10842 27872
rect 13446 27820 13452 27872
rect 13504 27820 13510 27872
rect 15194 27820 15200 27872
rect 15252 27860 15258 27872
rect 16114 27860 16120 27872
rect 15252 27832 16120 27860
rect 15252 27820 15258 27832
rect 16114 27820 16120 27832
rect 16172 27820 16178 27872
rect 16666 27820 16672 27872
rect 16724 27820 16730 27872
rect 25685 27863 25743 27869
rect 25685 27829 25697 27863
rect 25731 27860 25743 27863
rect 25866 27860 25872 27872
rect 25731 27832 25872 27860
rect 25731 27829 25743 27832
rect 25685 27823 25743 27829
rect 25866 27820 25872 27832
rect 25924 27820 25930 27872
rect 30650 27820 30656 27872
rect 30708 27860 30714 27872
rect 30837 27863 30895 27869
rect 30837 27860 30849 27863
rect 30708 27832 30849 27860
rect 30708 27820 30714 27832
rect 30837 27829 30849 27832
rect 30883 27829 30895 27863
rect 30837 27823 30895 27829
rect 1104 27770 37076 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 37076 27770
rect 1104 27696 37076 27718
rect 2130 27665 2136 27668
rect 2120 27659 2136 27665
rect 2120 27625 2132 27659
rect 2120 27619 2136 27625
rect 2130 27616 2136 27619
rect 2188 27616 2194 27668
rect 3602 27616 3608 27668
rect 3660 27616 3666 27668
rect 4157 27659 4215 27665
rect 4157 27625 4169 27659
rect 4203 27656 4215 27659
rect 4614 27656 4620 27668
rect 4203 27628 4620 27656
rect 4203 27625 4215 27628
rect 4157 27619 4215 27625
rect 4614 27616 4620 27628
rect 4672 27616 4678 27668
rect 5718 27616 5724 27668
rect 5776 27656 5782 27668
rect 6365 27659 6423 27665
rect 6365 27656 6377 27659
rect 5776 27628 6377 27656
rect 5776 27616 5782 27628
rect 6365 27625 6377 27628
rect 6411 27656 6423 27659
rect 6822 27656 6828 27668
rect 6411 27628 6828 27656
rect 6411 27625 6423 27628
rect 6365 27619 6423 27625
rect 6822 27616 6828 27628
rect 6880 27616 6886 27668
rect 9030 27616 9036 27668
rect 9088 27656 9094 27668
rect 9493 27659 9551 27665
rect 9493 27656 9505 27659
rect 9088 27628 9505 27656
rect 9088 27616 9094 27628
rect 9493 27625 9505 27628
rect 9539 27625 9551 27659
rect 9493 27619 9551 27625
rect 18138 27616 18144 27668
rect 18196 27656 18202 27668
rect 18233 27659 18291 27665
rect 18233 27656 18245 27659
rect 18196 27628 18245 27656
rect 18196 27616 18202 27628
rect 18233 27625 18245 27628
rect 18279 27625 18291 27659
rect 19334 27656 19340 27668
rect 18233 27619 18291 27625
rect 19260 27628 19340 27656
rect 3418 27548 3424 27600
rect 3476 27588 3482 27600
rect 4062 27588 4068 27600
rect 3476 27560 4068 27588
rect 3476 27548 3482 27560
rect 4062 27548 4068 27560
rect 4120 27588 4126 27600
rect 5261 27591 5319 27597
rect 5261 27588 5273 27591
rect 4120 27560 5273 27588
rect 4120 27548 4126 27560
rect 5261 27557 5273 27560
rect 5307 27588 5319 27591
rect 6546 27588 6552 27600
rect 5307 27560 6552 27588
rect 5307 27557 5319 27560
rect 5261 27551 5319 27557
rect 6546 27548 6552 27560
rect 6604 27548 6610 27600
rect 12069 27591 12127 27597
rect 12069 27588 12081 27591
rect 11624 27560 12081 27588
rect 3142 27480 3148 27532
rect 3200 27520 3206 27532
rect 3789 27523 3847 27529
rect 3789 27520 3801 27523
rect 3200 27492 3801 27520
rect 3200 27480 3206 27492
rect 3789 27489 3801 27492
rect 3835 27489 3847 27523
rect 3789 27483 3847 27489
rect 6086 27480 6092 27532
rect 6144 27520 6150 27532
rect 7837 27523 7895 27529
rect 7837 27520 7849 27523
rect 6144 27492 7849 27520
rect 6144 27480 6150 27492
rect 7837 27489 7849 27492
rect 7883 27489 7895 27523
rect 7837 27483 7895 27489
rect 8113 27523 8171 27529
rect 8113 27489 8125 27523
rect 8159 27520 8171 27523
rect 8202 27520 8208 27532
rect 8159 27492 8208 27520
rect 8159 27489 8171 27492
rect 8113 27483 8171 27489
rect 8202 27480 8208 27492
rect 8260 27520 8266 27532
rect 8260 27492 10364 27520
rect 8260 27480 8266 27492
rect 10336 27464 10364 27492
rect 10594 27480 10600 27532
rect 10652 27520 10658 27532
rect 11624 27520 11652 27560
rect 12069 27557 12081 27560
rect 12115 27557 12127 27591
rect 12069 27551 12127 27557
rect 16298 27548 16304 27600
rect 16356 27548 16362 27600
rect 16390 27548 16396 27600
rect 16448 27588 16454 27600
rect 19260 27588 19288 27628
rect 19334 27616 19340 27628
rect 19392 27616 19398 27668
rect 19518 27665 19524 27668
rect 19508 27659 19524 27665
rect 19508 27625 19520 27659
rect 19508 27619 19524 27625
rect 19518 27616 19524 27619
rect 19576 27616 19582 27668
rect 19886 27616 19892 27668
rect 19944 27656 19950 27668
rect 25130 27656 25136 27668
rect 19944 27628 21036 27656
rect 19944 27616 19950 27628
rect 21008 27597 21036 27628
rect 24872 27628 25136 27656
rect 16448 27560 16896 27588
rect 16448 27548 16454 27560
rect 10652 27492 11652 27520
rect 10652 27480 10658 27492
rect 11790 27480 11796 27532
rect 11848 27520 11854 27532
rect 12161 27523 12219 27529
rect 12161 27520 12173 27523
rect 11848 27492 12173 27520
rect 11848 27480 11854 27492
rect 12161 27489 12173 27492
rect 12207 27520 12219 27523
rect 12802 27520 12808 27532
rect 12207 27492 12808 27520
rect 12207 27489 12219 27492
rect 12161 27483 12219 27489
rect 12802 27480 12808 27492
rect 12860 27520 12866 27532
rect 14826 27520 14832 27532
rect 12860 27492 14832 27520
rect 12860 27480 12866 27492
rect 14826 27480 14832 27492
rect 14884 27520 14890 27532
rect 14884 27492 15884 27520
rect 14884 27480 14890 27492
rect 1394 27412 1400 27464
rect 1452 27452 1458 27464
rect 1854 27452 1860 27464
rect 1452 27424 1860 27452
rect 1452 27412 1458 27424
rect 1854 27412 1860 27424
rect 1912 27412 1918 27464
rect 3602 27412 3608 27464
rect 3660 27452 3666 27464
rect 3973 27455 4031 27461
rect 3973 27452 3985 27455
rect 3660 27424 3985 27452
rect 3660 27412 3666 27424
rect 3973 27421 3985 27424
rect 4019 27421 4031 27455
rect 3973 27415 4031 27421
rect 5442 27412 5448 27464
rect 5500 27412 5506 27464
rect 5534 27412 5540 27464
rect 5592 27452 5598 27464
rect 5629 27455 5687 27461
rect 5629 27452 5641 27455
rect 5592 27424 5641 27452
rect 5592 27412 5598 27424
rect 5629 27421 5641 27424
rect 5675 27452 5687 27455
rect 5810 27452 5816 27464
rect 5675 27424 5816 27452
rect 5675 27421 5687 27424
rect 5629 27415 5687 27421
rect 5810 27412 5816 27424
rect 5868 27412 5874 27464
rect 6273 27455 6331 27461
rect 6273 27421 6285 27455
rect 6319 27421 6331 27455
rect 6273 27415 6331 27421
rect 2866 27344 2872 27396
rect 2924 27344 2930 27396
rect 6288 27384 6316 27415
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 9217 27455 9275 27461
rect 9217 27452 9229 27455
rect 9180 27424 9229 27452
rect 9180 27412 9186 27424
rect 9217 27421 9229 27424
rect 9263 27421 9275 27455
rect 9217 27415 9275 27421
rect 9401 27455 9459 27461
rect 9401 27421 9413 27455
rect 9447 27421 9459 27455
rect 9401 27415 9459 27421
rect 5828 27356 6316 27384
rect 5350 27276 5356 27328
rect 5408 27316 5414 27328
rect 5828 27325 5856 27356
rect 5537 27319 5595 27325
rect 5537 27316 5549 27319
rect 5408 27288 5549 27316
rect 5408 27276 5414 27288
rect 5537 27285 5549 27288
rect 5583 27285 5595 27319
rect 5537 27279 5595 27285
rect 5813 27319 5871 27325
rect 5813 27285 5825 27319
rect 5859 27285 5871 27319
rect 5813 27279 5871 27285
rect 6178 27276 6184 27328
rect 6236 27276 6242 27328
rect 6288 27316 6316 27356
rect 6454 27344 6460 27396
rect 6512 27384 6518 27396
rect 9416 27384 9444 27415
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 9677 27455 9735 27461
rect 9677 27452 9689 27455
rect 9640 27424 9689 27452
rect 9640 27412 9646 27424
rect 9677 27421 9689 27424
rect 9723 27421 9735 27455
rect 9677 27415 9735 27421
rect 9953 27455 10011 27461
rect 9953 27421 9965 27455
rect 9999 27452 10011 27455
rect 10042 27452 10048 27464
rect 9999 27424 10048 27452
rect 9999 27421 10011 27424
rect 9953 27415 10011 27421
rect 10042 27412 10048 27424
rect 10100 27412 10106 27464
rect 10134 27412 10140 27464
rect 10192 27412 10198 27464
rect 10318 27412 10324 27464
rect 10376 27412 10382 27464
rect 15856 27461 15884 27492
rect 16666 27480 16672 27532
rect 16724 27520 16730 27532
rect 16868 27529 16896 27560
rect 18892 27560 19288 27588
rect 20993 27591 21051 27597
rect 18892 27532 18920 27560
rect 20993 27557 21005 27591
rect 21039 27557 21051 27591
rect 24872 27588 24900 27628
rect 25130 27616 25136 27628
rect 25188 27616 25194 27668
rect 25498 27616 25504 27668
rect 25556 27656 25562 27668
rect 31039 27659 31097 27665
rect 25556 27628 26234 27656
rect 25556 27616 25562 27628
rect 20993 27551 21051 27557
rect 23768 27560 24900 27588
rect 26206 27588 26234 27628
rect 31039 27625 31051 27659
rect 31085 27656 31097 27659
rect 32122 27656 32128 27668
rect 31085 27628 32128 27656
rect 31085 27625 31097 27628
rect 31039 27619 31097 27625
rect 32122 27616 32128 27628
rect 32180 27616 32186 27668
rect 32480 27659 32538 27665
rect 32480 27625 32492 27659
rect 32526 27656 32538 27659
rect 33226 27656 33232 27668
rect 32526 27628 33232 27656
rect 32526 27625 32538 27628
rect 32480 27619 32538 27625
rect 33226 27616 33232 27628
rect 33284 27616 33290 27668
rect 33962 27616 33968 27668
rect 34020 27616 34026 27668
rect 26206 27560 27660 27588
rect 16761 27523 16819 27529
rect 16761 27520 16773 27523
rect 16724 27492 16773 27520
rect 16724 27480 16730 27492
rect 16761 27489 16773 27492
rect 16807 27489 16819 27523
rect 16761 27483 16819 27489
rect 16853 27523 16911 27529
rect 16853 27489 16865 27523
rect 16899 27489 16911 27523
rect 16853 27483 16911 27489
rect 17681 27523 17739 27529
rect 17681 27489 17693 27523
rect 17727 27520 17739 27523
rect 17954 27520 17960 27532
rect 17727 27492 17960 27520
rect 17727 27489 17739 27492
rect 17681 27483 17739 27489
rect 15841 27455 15899 27461
rect 15841 27421 15853 27455
rect 15887 27452 15899 27455
rect 16390 27452 16396 27464
rect 15887 27424 16396 27452
rect 15887 27421 15899 27424
rect 15841 27415 15899 27421
rect 16390 27412 16396 27424
rect 16448 27412 16454 27464
rect 16776 27452 16804 27483
rect 17954 27480 17960 27492
rect 18012 27520 18018 27532
rect 18874 27520 18880 27532
rect 18012 27492 18880 27520
rect 18012 27480 18018 27492
rect 18874 27480 18880 27492
rect 18932 27480 18938 27532
rect 19242 27480 19248 27532
rect 19300 27520 19306 27532
rect 21177 27523 21235 27529
rect 21177 27520 21189 27523
rect 19300 27492 21189 27520
rect 19300 27480 19306 27492
rect 21177 27489 21189 27492
rect 21223 27489 21235 27523
rect 21177 27483 21235 27489
rect 22646 27480 22652 27532
rect 22704 27520 22710 27532
rect 23768 27529 23796 27560
rect 23569 27523 23627 27529
rect 23569 27520 23581 27523
rect 22704 27492 23581 27520
rect 22704 27480 22710 27492
rect 23569 27489 23581 27492
rect 23615 27489 23627 27523
rect 23569 27483 23627 27489
rect 23753 27523 23811 27529
rect 23753 27489 23765 27523
rect 23799 27489 23811 27523
rect 23753 27483 23811 27489
rect 24854 27480 24860 27532
rect 24912 27520 24918 27532
rect 26142 27520 26148 27532
rect 24912 27492 26148 27520
rect 24912 27480 24918 27492
rect 26142 27480 26148 27492
rect 26200 27480 26206 27532
rect 27632 27529 27660 27560
rect 27617 27523 27675 27529
rect 27617 27489 27629 27523
rect 27663 27520 27675 27523
rect 28905 27523 28963 27529
rect 28905 27520 28917 27523
rect 27663 27492 28917 27520
rect 27663 27489 27675 27492
rect 27617 27483 27675 27489
rect 28905 27489 28917 27492
rect 28951 27520 28963 27523
rect 30466 27520 30472 27532
rect 28951 27492 30472 27520
rect 28951 27489 28963 27492
rect 28905 27483 28963 27489
rect 30466 27480 30472 27492
rect 30524 27480 30530 27532
rect 17865 27455 17923 27461
rect 17865 27452 17877 27455
rect 16776 27424 17877 27452
rect 17865 27421 17877 27424
rect 17911 27421 17923 27455
rect 22005 27455 22063 27461
rect 22005 27452 22017 27455
rect 17865 27415 17923 27421
rect 20916 27424 22017 27452
rect 10502 27384 10508 27396
rect 6512 27356 6670 27384
rect 9416 27356 10508 27384
rect 6512 27344 6518 27356
rect 10502 27344 10508 27356
rect 10560 27344 10566 27396
rect 10597 27387 10655 27393
rect 10597 27353 10609 27387
rect 10643 27384 10655 27387
rect 10870 27384 10876 27396
rect 10643 27356 10876 27384
rect 10643 27353 10655 27356
rect 10597 27347 10655 27353
rect 10870 27344 10876 27356
rect 10928 27344 10934 27396
rect 11054 27344 11060 27396
rect 11112 27344 11118 27396
rect 12434 27344 12440 27396
rect 12492 27344 12498 27396
rect 13722 27384 13728 27396
rect 13662 27356 13728 27384
rect 13722 27344 13728 27356
rect 13780 27384 13786 27396
rect 13780 27356 14320 27384
rect 13780 27344 13786 27356
rect 6914 27316 6920 27328
rect 6288 27288 6920 27316
rect 6914 27276 6920 27288
rect 6972 27316 6978 27328
rect 8110 27316 8116 27328
rect 6972 27288 8116 27316
rect 6972 27276 6978 27288
rect 8110 27276 8116 27288
rect 8168 27276 8174 27328
rect 9401 27319 9459 27325
rect 9401 27285 9413 27319
rect 9447 27316 9459 27319
rect 10962 27316 10968 27328
rect 9447 27288 10968 27316
rect 9447 27285 9459 27288
rect 9401 27279 9459 27285
rect 10962 27276 10968 27288
rect 11020 27276 11026 27328
rect 13354 27276 13360 27328
rect 13412 27316 13418 27328
rect 13909 27319 13967 27325
rect 13909 27316 13921 27319
rect 13412 27288 13921 27316
rect 13412 27276 13418 27288
rect 13909 27285 13921 27288
rect 13955 27285 13967 27319
rect 13909 27279 13967 27285
rect 14090 27276 14096 27328
rect 14148 27276 14154 27328
rect 14292 27316 14320 27356
rect 15102 27344 15108 27396
rect 15160 27384 15166 27396
rect 15160 27356 15240 27384
rect 15160 27344 15166 27356
rect 15212 27316 15240 27356
rect 15562 27344 15568 27396
rect 15620 27344 15626 27396
rect 16669 27387 16727 27393
rect 16669 27353 16681 27387
rect 16715 27384 16727 27387
rect 16850 27384 16856 27396
rect 16715 27356 16856 27384
rect 16715 27353 16727 27356
rect 16669 27347 16727 27353
rect 16850 27344 16856 27356
rect 16908 27344 16914 27396
rect 17310 27344 17316 27396
rect 17368 27384 17374 27396
rect 17773 27387 17831 27393
rect 17773 27384 17785 27387
rect 17368 27356 17785 27384
rect 17368 27344 17374 27356
rect 17773 27353 17785 27356
rect 17819 27353 17831 27387
rect 20806 27384 20812 27396
rect 20746 27356 20812 27384
rect 17773 27347 17831 27353
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 14292 27288 15240 27316
rect 20438 27276 20444 27328
rect 20496 27316 20502 27328
rect 20916 27316 20944 27424
rect 22005 27421 22017 27424
rect 22051 27452 22063 27455
rect 24762 27452 24768 27464
rect 22051 27424 24768 27452
rect 22051 27421 22063 27424
rect 22005 27415 22063 27421
rect 24762 27412 24768 27424
rect 24820 27412 24826 27464
rect 26970 27412 26976 27464
rect 27028 27452 27034 27464
rect 27801 27455 27859 27461
rect 27801 27452 27813 27455
rect 27028 27424 27813 27452
rect 27028 27412 27034 27424
rect 27801 27421 27813 27424
rect 27847 27421 27859 27455
rect 27801 27415 27859 27421
rect 31294 27412 31300 27464
rect 31352 27452 31358 27464
rect 32217 27455 32275 27461
rect 32217 27452 32229 27455
rect 31352 27424 32229 27452
rect 31352 27412 31358 27424
rect 32217 27421 32229 27424
rect 32263 27421 32275 27455
rect 32217 27415 32275 27421
rect 22186 27344 22192 27396
rect 22244 27384 22250 27396
rect 22557 27387 22615 27393
rect 22557 27384 22569 27387
rect 22244 27356 22569 27384
rect 22244 27344 22250 27356
rect 22557 27353 22569 27356
rect 22603 27353 22615 27387
rect 22557 27347 22615 27353
rect 23290 27344 23296 27396
rect 23348 27384 23354 27396
rect 23845 27387 23903 27393
rect 23845 27384 23857 27387
rect 23348 27356 23857 27384
rect 23348 27344 23354 27356
rect 23845 27353 23857 27356
rect 23891 27353 23903 27387
rect 23845 27347 23903 27353
rect 25130 27344 25136 27396
rect 25188 27344 25194 27396
rect 27522 27384 27528 27396
rect 26358 27356 27528 27384
rect 27522 27344 27528 27356
rect 27580 27344 27586 27396
rect 28629 27387 28687 27393
rect 28629 27384 28641 27387
rect 27724 27356 28641 27384
rect 27724 27328 27752 27356
rect 28629 27353 28641 27356
rect 28675 27353 28687 27387
rect 28629 27347 28687 27353
rect 30558 27344 30564 27396
rect 30616 27384 30622 27396
rect 30742 27384 30748 27396
rect 30616 27356 30748 27384
rect 30616 27344 30622 27356
rect 30742 27344 30748 27356
rect 30800 27344 30806 27396
rect 33134 27344 33140 27396
rect 33192 27344 33198 27396
rect 20496 27288 20944 27316
rect 20496 27276 20502 27288
rect 22094 27276 22100 27328
rect 22152 27276 22158 27328
rect 22462 27276 22468 27328
rect 22520 27276 22526 27328
rect 24213 27319 24271 27325
rect 24213 27285 24225 27319
rect 24259 27316 24271 27319
rect 25314 27316 25320 27328
rect 24259 27288 25320 27316
rect 24259 27285 24271 27288
rect 24213 27279 24271 27285
rect 25314 27276 25320 27288
rect 25372 27276 25378 27328
rect 25958 27276 25964 27328
rect 26016 27316 26022 27328
rect 26605 27319 26663 27325
rect 26605 27316 26617 27319
rect 26016 27288 26617 27316
rect 26016 27276 26022 27288
rect 26605 27285 26617 27288
rect 26651 27285 26663 27319
rect 26605 27279 26663 27285
rect 27706 27276 27712 27328
rect 27764 27276 27770 27328
rect 28166 27276 28172 27328
rect 28224 27276 28230 27328
rect 28261 27319 28319 27325
rect 28261 27285 28273 27319
rect 28307 27316 28319 27319
rect 28442 27316 28448 27328
rect 28307 27288 28448 27316
rect 28307 27285 28319 27288
rect 28261 27279 28319 27285
rect 28442 27276 28448 27288
rect 28500 27276 28506 27328
rect 28721 27319 28779 27325
rect 28721 27285 28733 27319
rect 28767 27316 28779 27319
rect 29178 27316 29184 27328
rect 28767 27288 29184 27316
rect 28767 27285 28779 27288
rect 28721 27279 28779 27285
rect 29178 27276 29184 27288
rect 29236 27276 29242 27328
rect 29549 27319 29607 27325
rect 29549 27285 29561 27319
rect 29595 27316 29607 27319
rect 31018 27316 31024 27328
rect 29595 27288 31024 27316
rect 29595 27285 29607 27288
rect 29549 27279 29607 27285
rect 31018 27276 31024 27288
rect 31076 27276 31082 27328
rect 1104 27226 37076 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 37076 27226
rect 1104 27152 37076 27174
rect 5534 27072 5540 27124
rect 5592 27121 5598 27124
rect 5592 27115 5611 27121
rect 5599 27081 5611 27115
rect 5592 27075 5611 27081
rect 6023 27115 6081 27121
rect 6023 27081 6035 27115
rect 6069 27112 6081 27115
rect 6178 27112 6184 27124
rect 6069 27084 6184 27112
rect 6069 27081 6081 27084
rect 6023 27075 6081 27081
rect 5592 27072 5598 27075
rect 6178 27072 6184 27084
rect 6236 27072 6242 27124
rect 8573 27115 8631 27121
rect 8573 27081 8585 27115
rect 8619 27112 8631 27115
rect 10413 27115 10471 27121
rect 10413 27112 10425 27115
rect 8619 27084 10425 27112
rect 8619 27081 8631 27084
rect 8573 27075 8631 27081
rect 10413 27081 10425 27084
rect 10459 27081 10471 27115
rect 10413 27075 10471 27081
rect 10686 27072 10692 27124
rect 10744 27112 10750 27124
rect 11057 27115 11115 27121
rect 11057 27112 11069 27115
rect 10744 27084 11069 27112
rect 10744 27072 10750 27084
rect 11057 27081 11069 27084
rect 11103 27081 11115 27115
rect 11057 27075 11115 27081
rect 13354 27072 13360 27124
rect 13412 27072 13418 27124
rect 13817 27115 13875 27121
rect 13817 27081 13829 27115
rect 13863 27112 13875 27115
rect 15562 27112 15568 27124
rect 13863 27084 15568 27112
rect 13863 27081 13875 27084
rect 13817 27075 13875 27081
rect 15562 27072 15568 27084
rect 15620 27072 15626 27124
rect 18693 27115 18751 27121
rect 18693 27081 18705 27115
rect 18739 27112 18751 27115
rect 19426 27112 19432 27124
rect 18739 27084 19432 27112
rect 18739 27081 18751 27084
rect 18693 27075 18751 27081
rect 19426 27072 19432 27084
rect 19484 27072 19490 27124
rect 20806 27072 20812 27124
rect 20864 27112 20870 27124
rect 20864 27084 21496 27112
rect 20864 27072 20870 27084
rect 2958 27044 2964 27056
rect 2898 27016 2964 27044
rect 2958 27004 2964 27016
rect 3016 27004 3022 27056
rect 5353 27047 5411 27053
rect 5353 27013 5365 27047
rect 5399 27044 5411 27047
rect 5442 27044 5448 27056
rect 5399 27016 5448 27044
rect 5399 27013 5411 27016
rect 5353 27007 5411 27013
rect 5442 27004 5448 27016
rect 5500 27004 5506 27056
rect 5810 27004 5816 27056
rect 5868 27004 5874 27056
rect 6503 27013 6561 27019
rect 4798 26936 4804 26988
rect 4856 26976 4862 26988
rect 4893 26979 4951 26985
rect 4893 26976 4905 26979
rect 4856 26948 4905 26976
rect 4856 26936 4862 26948
rect 4893 26945 4905 26948
rect 4939 26945 4951 26979
rect 4893 26939 4951 26945
rect 5258 26936 5264 26988
rect 5316 26976 5322 26988
rect 6503 26979 6515 27013
rect 6549 27010 6561 27013
rect 6549 26982 6684 27010
rect 6730 27004 6736 27056
rect 6788 27004 6794 27056
rect 6822 27004 6828 27056
rect 6880 27044 6886 27056
rect 6917 27047 6975 27053
rect 6917 27044 6929 27047
rect 6880 27016 6929 27044
rect 6880 27004 6886 27016
rect 6917 27013 6929 27016
rect 6963 27013 6975 27047
rect 6917 27007 6975 27013
rect 7133 27047 7191 27053
rect 7133 27013 7145 27047
rect 7179 27044 7191 27047
rect 7745 27047 7803 27053
rect 7179 27016 7696 27044
rect 7179 27013 7191 27016
rect 7133 27007 7191 27013
rect 7668 26985 7696 27016
rect 7745 27013 7757 27047
rect 7791 27044 7803 27047
rect 7791 27016 8524 27044
rect 7791 27013 7803 27016
rect 7745 27007 7803 27013
rect 6549 26979 6561 26982
rect 5316 26948 6408 26976
rect 6503 26973 6561 26979
rect 6656 26976 6684 26982
rect 7561 26979 7619 26985
rect 7561 26976 7573 26979
rect 6656 26948 7573 26976
rect 5316 26936 5322 26948
rect 1397 26911 1455 26917
rect 1397 26877 1409 26911
rect 1443 26877 1455 26911
rect 1397 26871 1455 26877
rect 1412 26772 1440 26871
rect 1670 26868 1676 26920
rect 1728 26868 1734 26920
rect 4706 26908 4712 26920
rect 2746 26880 4712 26908
rect 1854 26772 1860 26784
rect 1412 26744 1860 26772
rect 1854 26732 1860 26744
rect 1912 26772 1918 26784
rect 2746 26772 2774 26880
rect 4706 26868 4712 26880
rect 4764 26868 4770 26920
rect 5169 26911 5227 26917
rect 5169 26877 5181 26911
rect 5215 26908 5227 26911
rect 5902 26908 5908 26920
rect 5215 26880 5908 26908
rect 5215 26877 5227 26880
rect 5169 26871 5227 26877
rect 5902 26868 5908 26880
rect 5960 26868 5966 26920
rect 6380 26908 6408 26948
rect 6822 26908 6828 26920
rect 6380 26880 6828 26908
rect 5077 26843 5135 26849
rect 5077 26809 5089 26843
rect 5123 26840 5135 26843
rect 6365 26843 6423 26849
rect 6365 26840 6377 26843
rect 5123 26812 6377 26840
rect 5123 26809 5135 26812
rect 5077 26803 5135 26809
rect 6365 26809 6377 26812
rect 6411 26840 6423 26843
rect 6454 26840 6460 26852
rect 6411 26812 6460 26840
rect 6411 26809 6423 26812
rect 6365 26803 6423 26809
rect 6454 26800 6460 26812
rect 6512 26800 6518 26852
rect 1912 26744 2774 26772
rect 1912 26732 1918 26744
rect 3142 26732 3148 26784
rect 3200 26732 3206 26784
rect 4614 26732 4620 26784
rect 4672 26772 4678 26784
rect 4709 26775 4767 26781
rect 4709 26772 4721 26775
rect 4672 26744 4721 26772
rect 4672 26732 4678 26744
rect 4709 26741 4721 26744
rect 4755 26741 4767 26775
rect 4709 26735 4767 26741
rect 5350 26732 5356 26784
rect 5408 26772 5414 26784
rect 5537 26775 5595 26781
rect 5537 26772 5549 26775
rect 5408 26744 5549 26772
rect 5408 26732 5414 26744
rect 5537 26741 5549 26744
rect 5583 26741 5595 26775
rect 5537 26735 5595 26741
rect 5626 26732 5632 26784
rect 5684 26772 5690 26784
rect 5721 26775 5779 26781
rect 5721 26772 5733 26775
rect 5684 26744 5733 26772
rect 5684 26732 5690 26744
rect 5721 26741 5733 26744
rect 5767 26741 5779 26775
rect 5721 26735 5779 26741
rect 5994 26732 6000 26784
rect 6052 26732 6058 26784
rect 6086 26732 6092 26784
rect 6144 26772 6150 26784
rect 6564 26781 6592 26880
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 7116 26784 7144 26948
rect 7561 26945 7573 26948
rect 7607 26945 7619 26979
rect 7561 26939 7619 26945
rect 7653 26979 7711 26985
rect 7653 26945 7665 26979
rect 7699 26976 7711 26979
rect 8386 26976 8392 26988
rect 7699 26948 8392 26976
rect 7699 26945 7711 26948
rect 7653 26939 7711 26945
rect 8386 26936 8392 26948
rect 8444 26936 8450 26988
rect 8496 26985 8524 27016
rect 8754 27004 8760 27056
rect 8812 27044 8818 27056
rect 9582 27044 9588 27056
rect 8812 27016 9588 27044
rect 8812 27004 8818 27016
rect 9582 27004 9588 27016
rect 9640 27004 9646 27056
rect 9953 27047 10011 27053
rect 9953 27013 9965 27047
rect 9999 27013 10011 27047
rect 9953 27007 10011 27013
rect 8481 26979 8539 26985
rect 8481 26945 8493 26979
rect 8527 26976 8539 26979
rect 9490 26976 9496 26988
rect 8527 26948 9496 26976
rect 8527 26945 8539 26948
rect 8481 26939 8539 26945
rect 9490 26936 9496 26948
rect 9548 26936 9554 26988
rect 9968 26976 9996 27007
rect 10042 27004 10048 27056
rect 10100 27044 10106 27056
rect 10153 27047 10211 27053
rect 10153 27044 10165 27047
rect 10100 27016 10165 27044
rect 10100 27004 10106 27016
rect 10153 27013 10165 27016
rect 10199 27044 10211 27047
rect 10565 27047 10623 27053
rect 10565 27044 10577 27047
rect 10199 27016 10577 27044
rect 10199 27013 10211 27016
rect 10153 27007 10211 27013
rect 10565 27013 10577 27016
rect 10611 27013 10623 27047
rect 10565 27007 10623 27013
rect 10781 27047 10839 27053
rect 10781 27013 10793 27047
rect 10827 27013 10839 27047
rect 10781 27007 10839 27013
rect 10410 26976 10416 26988
rect 9968 26948 10416 26976
rect 10410 26936 10416 26948
rect 10468 26976 10474 26988
rect 10796 26976 10824 27007
rect 10962 27004 10968 27056
rect 11020 27044 11026 27056
rect 14093 27047 14151 27053
rect 11020 27016 11192 27044
rect 11020 27004 11026 27016
rect 11164 26985 11192 27016
rect 14093 27013 14105 27047
rect 14139 27044 14151 27047
rect 14734 27044 14740 27056
rect 14139 27016 14740 27044
rect 14139 27013 14151 27016
rect 14093 27007 14151 27013
rect 14734 27004 14740 27016
rect 14792 27004 14798 27056
rect 20438 27044 20444 27056
rect 15856 27016 20444 27044
rect 15856 26985 15884 27016
rect 20438 27004 20444 27016
rect 20496 27004 20502 27056
rect 20714 27004 20720 27056
rect 20772 27004 20778 27056
rect 21468 27044 21496 27084
rect 21818 27072 21824 27124
rect 21876 27112 21882 27124
rect 22462 27112 22468 27124
rect 21876 27084 22468 27112
rect 21876 27072 21882 27084
rect 22462 27072 22468 27084
rect 22520 27072 22526 27124
rect 24946 27072 24952 27124
rect 25004 27112 25010 27124
rect 25682 27112 25688 27124
rect 25004 27084 25688 27112
rect 25004 27072 25010 27084
rect 25682 27072 25688 27084
rect 25740 27112 25746 27124
rect 30926 27112 30932 27124
rect 25740 27084 30932 27112
rect 25740 27072 25746 27084
rect 30926 27072 30932 27084
rect 30984 27072 30990 27124
rect 31018 27072 31024 27124
rect 31076 27112 31082 27124
rect 31076 27084 32904 27112
rect 31076 27072 31082 27084
rect 21468 27016 22310 27044
rect 23842 27004 23848 27056
rect 23900 27044 23906 27056
rect 23900 27016 24150 27044
rect 23900 27004 23906 27016
rect 25314 27004 25320 27056
rect 25372 27004 25378 27056
rect 26142 27044 26148 27056
rect 25608 27016 26148 27044
rect 10468 26948 10824 26976
rect 10873 26979 10931 26985
rect 10468 26936 10474 26948
rect 10873 26945 10885 26979
rect 10919 26966 10931 26979
rect 11149 26979 11207 26985
rect 10919 26945 11008 26966
rect 10873 26939 11008 26945
rect 11149 26945 11161 26979
rect 11195 26945 11207 26979
rect 11149 26939 11207 26945
rect 13449 26979 13507 26985
rect 13449 26945 13461 26979
rect 13495 26945 13507 26979
rect 13449 26939 13507 26945
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26976 14887 26979
rect 15841 26979 15899 26985
rect 15841 26976 15853 26979
rect 14875 26948 15853 26976
rect 14875 26945 14887 26948
rect 14829 26939 14887 26945
rect 15841 26945 15853 26948
rect 15887 26945 15899 26979
rect 15841 26939 15899 26945
rect 10888 26938 11008 26939
rect 9858 26908 9864 26920
rect 7300 26880 9864 26908
rect 7300 26849 7328 26880
rect 9858 26868 9864 26880
rect 9916 26868 9922 26920
rect 10134 26868 10140 26920
rect 10192 26908 10198 26920
rect 10980 26908 11008 26938
rect 10192 26880 11008 26908
rect 10192 26868 10198 26880
rect 7285 26843 7343 26849
rect 7285 26809 7297 26843
rect 7331 26809 7343 26843
rect 7285 26803 7343 26809
rect 7374 26800 7380 26852
rect 7432 26800 7438 26852
rect 8110 26800 8116 26852
rect 8168 26840 8174 26852
rect 10336 26849 10364 26880
rect 13262 26868 13268 26920
rect 13320 26868 13326 26920
rect 13464 26908 13492 26939
rect 16390 26936 16396 26988
rect 16448 26936 16454 26988
rect 17681 26979 17739 26985
rect 17681 26945 17693 26979
rect 17727 26976 17739 26979
rect 17727 26948 18460 26976
rect 17727 26945 17739 26948
rect 17681 26939 17739 26945
rect 14090 26908 14096 26920
rect 13464 26880 14096 26908
rect 14090 26868 14096 26880
rect 14148 26868 14154 26920
rect 14918 26868 14924 26920
rect 14976 26908 14982 26920
rect 15013 26911 15071 26917
rect 15013 26908 15025 26911
rect 14976 26880 15025 26908
rect 14976 26868 14982 26880
rect 15013 26877 15025 26880
rect 15059 26877 15071 26911
rect 15013 26871 15071 26877
rect 17034 26868 17040 26920
rect 17092 26908 17098 26920
rect 17770 26908 17776 26920
rect 17092 26880 17776 26908
rect 17092 26868 17098 26880
rect 17770 26868 17776 26880
rect 17828 26868 17834 26920
rect 17865 26911 17923 26917
rect 17865 26877 17877 26911
rect 17911 26877 17923 26911
rect 18432 26908 18460 26948
rect 19242 26936 19248 26988
rect 19300 26976 19306 26988
rect 25608 26985 25636 27016
rect 26142 27004 26148 27016
rect 26200 27044 26206 27056
rect 26421 27047 26479 27053
rect 26421 27044 26433 27047
rect 26200 27016 26433 27044
rect 26200 27004 26206 27016
rect 26421 27013 26433 27016
rect 26467 27013 26479 27047
rect 26421 27007 26479 27013
rect 27430 27004 27436 27056
rect 27488 27004 27494 27056
rect 28166 27004 28172 27056
rect 28224 27044 28230 27056
rect 28445 27047 28503 27053
rect 28445 27044 28457 27047
rect 28224 27016 28457 27044
rect 28224 27004 28230 27016
rect 28445 27013 28457 27016
rect 28491 27013 28503 27047
rect 30374 27044 30380 27056
rect 30222 27016 30380 27044
rect 28445 27007 28503 27013
rect 30374 27004 30380 27016
rect 30432 27044 30438 27056
rect 30558 27044 30564 27056
rect 30432 27016 30564 27044
rect 30432 27004 30438 27016
rect 30558 27004 30564 27016
rect 30616 27004 30622 27056
rect 30650 27004 30656 27056
rect 30708 27004 30714 27056
rect 32122 27004 32128 27056
rect 32180 27004 32186 27056
rect 19889 26979 19947 26985
rect 19889 26976 19901 26979
rect 19300 26948 19901 26976
rect 19300 26936 19306 26948
rect 19889 26945 19901 26948
rect 19935 26945 19947 26979
rect 19889 26939 19947 26945
rect 25593 26979 25651 26985
rect 25593 26945 25605 26979
rect 25639 26945 25651 26979
rect 25593 26939 25651 26945
rect 25682 26936 25688 26988
rect 25740 26936 25746 26988
rect 31021 26979 31079 26985
rect 31021 26976 31033 26979
rect 30944 26948 31033 26976
rect 18782 26908 18788 26920
rect 18432 26880 18788 26908
rect 17865 26871 17923 26877
rect 8205 26843 8263 26849
rect 8205 26840 8217 26843
rect 8168 26812 8217 26840
rect 8168 26800 8174 26812
rect 8205 26809 8217 26812
rect 8251 26809 8263 26843
rect 8205 26803 8263 26809
rect 10321 26843 10379 26849
rect 10321 26809 10333 26843
rect 10367 26809 10379 26843
rect 10321 26803 10379 26809
rect 10870 26800 10876 26852
rect 10928 26800 10934 26852
rect 16482 26800 16488 26852
rect 16540 26840 16546 26852
rect 17880 26840 17908 26871
rect 18782 26868 18788 26880
rect 18840 26868 18846 26920
rect 18874 26868 18880 26920
rect 18932 26868 18938 26920
rect 20165 26911 20223 26917
rect 20165 26877 20177 26911
rect 20211 26908 20223 26911
rect 22094 26908 22100 26920
rect 20211 26880 22100 26908
rect 20211 26877 20223 26880
rect 20165 26871 20223 26877
rect 22094 26868 22100 26880
rect 22152 26868 22158 26920
rect 22830 26868 22836 26920
rect 22888 26908 22894 26920
rect 23477 26911 23535 26917
rect 23477 26908 23489 26911
rect 22888 26880 23489 26908
rect 22888 26868 22894 26880
rect 23477 26877 23489 26880
rect 23523 26877 23535 26911
rect 23477 26871 23535 26877
rect 23753 26911 23811 26917
rect 23753 26877 23765 26911
rect 23799 26908 23811 26911
rect 24854 26908 24860 26920
rect 23799 26880 24860 26908
rect 23799 26877 23811 26880
rect 23753 26871 23811 26877
rect 24854 26868 24860 26880
rect 24912 26868 24918 26920
rect 26510 26868 26516 26920
rect 26568 26908 26574 26920
rect 26970 26908 26976 26920
rect 26568 26880 26976 26908
rect 26568 26868 26574 26880
rect 26970 26868 26976 26880
rect 27028 26868 27034 26920
rect 28721 26911 28779 26917
rect 28721 26877 28733 26911
rect 28767 26908 28779 26911
rect 28994 26908 29000 26920
rect 28767 26880 29000 26908
rect 28767 26877 28779 26880
rect 28721 26871 28779 26877
rect 28994 26868 29000 26880
rect 29052 26868 29058 26920
rect 29178 26868 29184 26920
rect 29236 26908 29242 26920
rect 30006 26908 30012 26920
rect 29236 26880 30012 26908
rect 29236 26868 29242 26880
rect 30006 26868 30012 26880
rect 30064 26868 30070 26920
rect 30944 26917 30972 26948
rect 31021 26945 31033 26948
rect 31067 26976 31079 26979
rect 31294 26976 31300 26988
rect 31067 26948 31300 26976
rect 31067 26945 31079 26948
rect 31021 26939 31079 26945
rect 31294 26936 31300 26948
rect 31352 26936 31358 26988
rect 31386 26936 31392 26988
rect 31444 26976 31450 26988
rect 32876 26985 32904 27084
rect 33226 27072 33232 27124
rect 33284 27072 33290 27124
rect 33597 27115 33655 27121
rect 33597 27081 33609 27115
rect 33643 27112 33655 27115
rect 33962 27112 33968 27124
rect 33643 27084 33968 27112
rect 33643 27081 33655 27084
rect 33597 27075 33655 27081
rect 33962 27072 33968 27084
rect 34020 27072 34026 27124
rect 32585 26979 32643 26985
rect 32585 26976 32597 26979
rect 31444 26948 32597 26976
rect 31444 26936 31450 26948
rect 32585 26945 32597 26948
rect 32631 26945 32643 26979
rect 32585 26939 32643 26945
rect 32769 26979 32827 26985
rect 32769 26945 32781 26979
rect 32815 26945 32827 26979
rect 32769 26939 32827 26945
rect 32861 26979 32919 26985
rect 32861 26945 32873 26979
rect 32907 26945 32919 26979
rect 32861 26939 32919 26945
rect 30929 26911 30987 26917
rect 30929 26877 30941 26911
rect 30975 26877 30987 26911
rect 30929 26871 30987 26877
rect 16540 26812 17908 26840
rect 16540 26800 16546 26812
rect 6181 26775 6239 26781
rect 6181 26772 6193 26775
rect 6144 26744 6193 26772
rect 6144 26732 6150 26744
rect 6181 26741 6193 26744
rect 6227 26741 6239 26775
rect 6181 26735 6239 26741
rect 6549 26775 6607 26781
rect 6549 26741 6561 26775
rect 6595 26741 6607 26775
rect 6549 26735 6607 26741
rect 7098 26732 7104 26784
rect 7156 26732 7162 26784
rect 7929 26775 7987 26781
rect 7929 26741 7941 26775
rect 7975 26772 7987 26775
rect 8938 26772 8944 26784
rect 7975 26744 8944 26772
rect 7975 26741 7987 26744
rect 7929 26735 7987 26741
rect 8938 26732 8944 26744
rect 8996 26772 9002 26784
rect 10137 26775 10195 26781
rect 10137 26772 10149 26775
rect 8996 26744 10149 26772
rect 8996 26732 9002 26744
rect 10137 26741 10149 26744
rect 10183 26741 10195 26775
rect 10137 26735 10195 26741
rect 10597 26775 10655 26781
rect 10597 26741 10609 26775
rect 10643 26772 10655 26775
rect 10778 26772 10784 26784
rect 10643 26744 10784 26772
rect 10643 26741 10655 26744
rect 10597 26735 10655 26741
rect 10778 26732 10784 26744
rect 10836 26732 10842 26784
rect 17218 26732 17224 26784
rect 17276 26772 17282 26784
rect 17313 26775 17371 26781
rect 17313 26772 17325 26775
rect 17276 26744 17325 26772
rect 17276 26732 17282 26744
rect 17313 26741 17325 26744
rect 17359 26741 17371 26775
rect 17313 26735 17371 26741
rect 17954 26732 17960 26784
rect 18012 26772 18018 26784
rect 18325 26775 18383 26781
rect 18325 26772 18337 26775
rect 18012 26744 18337 26772
rect 18012 26732 18018 26744
rect 18325 26741 18337 26744
rect 18371 26741 18383 26775
rect 18325 26735 18383 26741
rect 21637 26775 21695 26781
rect 21637 26741 21649 26775
rect 21683 26772 21695 26775
rect 21818 26772 21824 26784
rect 21683 26744 21824 26772
rect 21683 26741 21695 26744
rect 21637 26735 21695 26741
rect 21818 26732 21824 26744
rect 21876 26732 21882 26784
rect 22005 26775 22063 26781
rect 22005 26741 22017 26775
rect 22051 26772 22063 26775
rect 22278 26772 22284 26784
rect 22051 26744 22284 26772
rect 22051 26741 22063 26744
rect 22005 26735 22063 26741
rect 22278 26732 22284 26744
rect 22336 26732 22342 26784
rect 23290 26732 23296 26784
rect 23348 26772 23354 26784
rect 23845 26775 23903 26781
rect 23845 26772 23857 26775
rect 23348 26744 23857 26772
rect 23348 26732 23354 26744
rect 23845 26741 23857 26744
rect 23891 26741 23903 26775
rect 23845 26735 23903 26741
rect 30098 26732 30104 26784
rect 30156 26772 30162 26784
rect 30944 26772 30972 26871
rect 31478 26868 31484 26920
rect 31536 26908 31542 26920
rect 32784 26908 32812 26939
rect 31536 26880 32812 26908
rect 31536 26868 31542 26880
rect 33686 26868 33692 26920
rect 33744 26868 33750 26920
rect 33870 26868 33876 26920
rect 33928 26868 33934 26920
rect 33134 26800 33140 26852
rect 33192 26840 33198 26852
rect 34054 26840 34060 26852
rect 33192 26812 34060 26840
rect 33192 26800 33198 26812
rect 34054 26800 34060 26812
rect 34112 26800 34118 26852
rect 30156 26744 30972 26772
rect 30156 26732 30162 26744
rect 1104 26682 37076 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 37076 26682
rect 1104 26608 37076 26630
rect 1670 26528 1676 26580
rect 1728 26568 1734 26580
rect 1949 26571 2007 26577
rect 1949 26568 1961 26571
rect 1728 26540 1961 26568
rect 1728 26528 1734 26540
rect 1949 26537 1961 26540
rect 1995 26537 2007 26571
rect 1949 26531 2007 26537
rect 4420 26571 4478 26577
rect 4420 26537 4432 26571
rect 4466 26568 4478 26571
rect 4614 26568 4620 26580
rect 4466 26540 4620 26568
rect 4466 26537 4478 26540
rect 4420 26531 4478 26537
rect 4614 26528 4620 26540
rect 4672 26528 4678 26580
rect 5902 26528 5908 26580
rect 5960 26528 5966 26580
rect 6362 26528 6368 26580
rect 6420 26528 6426 26580
rect 8202 26528 8208 26580
rect 8260 26568 8266 26580
rect 8297 26571 8355 26577
rect 8297 26568 8309 26571
rect 8260 26540 8309 26568
rect 8260 26528 8266 26540
rect 8297 26537 8309 26540
rect 8343 26537 8355 26571
rect 8297 26531 8355 26537
rect 8938 26528 8944 26580
rect 8996 26568 9002 26580
rect 9493 26571 9551 26577
rect 9493 26568 9505 26571
rect 8996 26540 9505 26568
rect 8996 26528 9002 26540
rect 9493 26537 9505 26540
rect 9539 26537 9551 26571
rect 9493 26531 9551 26537
rect 10045 26571 10103 26577
rect 10045 26537 10057 26571
rect 10091 26568 10103 26571
rect 10686 26568 10692 26580
rect 10091 26540 10692 26568
rect 10091 26537 10103 26540
rect 10045 26531 10103 26537
rect 5810 26460 5816 26512
rect 5868 26500 5874 26512
rect 9122 26500 9128 26512
rect 5868 26472 9128 26500
rect 5868 26460 5874 26472
rect 9122 26460 9128 26472
rect 9180 26460 9186 26512
rect 9214 26460 9220 26512
rect 9272 26460 9278 26512
rect 2593 26435 2651 26441
rect 2593 26401 2605 26435
rect 2639 26432 2651 26435
rect 3142 26432 3148 26444
rect 2639 26404 3148 26432
rect 2639 26401 2651 26404
rect 2593 26395 2651 26401
rect 3142 26392 3148 26404
rect 3200 26392 3206 26444
rect 4157 26435 4215 26441
rect 4157 26401 4169 26435
rect 4203 26432 4215 26435
rect 4522 26432 4528 26444
rect 4203 26404 4528 26432
rect 4203 26401 4215 26404
rect 4157 26395 4215 26401
rect 4522 26392 4528 26404
rect 4580 26392 4586 26444
rect 6270 26392 6276 26444
rect 6328 26432 6334 26444
rect 6457 26435 6515 26441
rect 6457 26432 6469 26435
rect 6328 26404 6469 26432
rect 6328 26392 6334 26404
rect 6457 26401 6469 26404
rect 6503 26401 6515 26435
rect 6457 26395 6515 26401
rect 6546 26392 6552 26444
rect 6604 26432 6610 26444
rect 7374 26432 7380 26444
rect 6604 26404 7380 26432
rect 6604 26392 6610 26404
rect 7374 26392 7380 26404
rect 7432 26392 7438 26444
rect 9140 26432 9168 26460
rect 9309 26435 9367 26441
rect 9309 26432 9321 26435
rect 9140 26404 9321 26432
rect 9309 26401 9321 26404
rect 9355 26401 9367 26435
rect 9508 26432 9536 26531
rect 10686 26528 10692 26540
rect 10744 26528 10750 26580
rect 12434 26528 12440 26580
rect 12492 26568 12498 26580
rect 12989 26571 13047 26577
rect 12989 26568 13001 26571
rect 12492 26540 13001 26568
rect 12492 26528 12498 26540
rect 12989 26537 13001 26540
rect 13035 26537 13047 26571
rect 12989 26531 13047 26537
rect 17770 26528 17776 26580
rect 17828 26568 17834 26580
rect 18877 26571 18935 26577
rect 18877 26568 18889 26571
rect 17828 26540 18889 26568
rect 17828 26528 17834 26540
rect 18877 26537 18889 26540
rect 18923 26537 18935 26571
rect 18877 26531 18935 26537
rect 22830 26528 22836 26580
rect 22888 26528 22894 26580
rect 24397 26571 24455 26577
rect 24397 26537 24409 26571
rect 24443 26568 24455 26571
rect 25222 26568 25228 26580
rect 24443 26540 25228 26568
rect 24443 26537 24455 26540
rect 24397 26531 24455 26537
rect 25222 26528 25228 26540
rect 25280 26528 25286 26580
rect 26973 26571 27031 26577
rect 26973 26537 26985 26571
rect 27019 26568 27031 26571
rect 27706 26568 27712 26580
rect 27019 26540 27712 26568
rect 27019 26537 27031 26540
rect 26973 26531 27031 26537
rect 27706 26528 27712 26540
rect 27764 26528 27770 26580
rect 31478 26528 31484 26580
rect 31536 26528 31542 26580
rect 13262 26460 13268 26512
rect 13320 26500 13326 26512
rect 16482 26500 16488 26512
rect 13320 26472 16488 26500
rect 13320 26460 13326 26472
rect 9508 26404 9996 26432
rect 9309 26395 9367 26401
rect 5718 26324 5724 26376
rect 5776 26364 5782 26376
rect 6641 26367 6699 26373
rect 6641 26364 6653 26367
rect 5776 26336 6653 26364
rect 5776 26324 5782 26336
rect 6641 26333 6653 26336
rect 6687 26333 6699 26367
rect 6641 26327 6699 26333
rect 8938 26324 8944 26376
rect 8996 26324 9002 26376
rect 9033 26367 9091 26373
rect 9033 26333 9045 26367
rect 9079 26364 9091 26367
rect 9585 26367 9643 26373
rect 9140 26364 9352 26366
rect 9585 26364 9597 26367
rect 9079 26338 9597 26364
rect 9079 26336 9168 26338
rect 9324 26336 9597 26338
rect 9079 26333 9091 26336
rect 9033 26327 9091 26333
rect 9585 26333 9597 26336
rect 9631 26364 9643 26367
rect 9674 26364 9680 26376
rect 9631 26336 9680 26364
rect 9631 26333 9643 26336
rect 9585 26327 9643 26333
rect 9674 26324 9680 26336
rect 9732 26324 9738 26376
rect 9968 26373 9996 26404
rect 13446 26392 13452 26444
rect 13504 26392 13510 26444
rect 13648 26441 13676 26472
rect 14752 26444 14780 26472
rect 16482 26460 16488 26472
rect 16540 26460 16546 26512
rect 21821 26503 21879 26509
rect 21821 26500 21833 26503
rect 21284 26472 21833 26500
rect 13633 26435 13691 26441
rect 13633 26401 13645 26435
rect 13679 26401 13691 26435
rect 13633 26395 13691 26401
rect 14090 26392 14096 26444
rect 14148 26432 14154 26444
rect 14553 26435 14611 26441
rect 14553 26432 14565 26435
rect 14148 26404 14565 26432
rect 14148 26392 14154 26404
rect 14553 26401 14565 26404
rect 14599 26401 14611 26435
rect 14553 26395 14611 26401
rect 14734 26392 14740 26444
rect 14792 26392 14798 26444
rect 16390 26392 16396 26444
rect 16448 26432 16454 26444
rect 17129 26435 17187 26441
rect 17129 26432 17141 26435
rect 16448 26404 17141 26432
rect 16448 26392 16454 26404
rect 17129 26401 17141 26404
rect 17175 26401 17187 26435
rect 17129 26395 17187 26401
rect 19242 26392 19248 26444
rect 19300 26432 19306 26444
rect 19981 26435 20039 26441
rect 19981 26432 19993 26435
rect 19300 26404 19993 26432
rect 19300 26392 19306 26404
rect 19981 26401 19993 26404
rect 20027 26401 20039 26435
rect 19981 26395 20039 26401
rect 20257 26435 20315 26441
rect 20257 26401 20269 26435
rect 20303 26432 20315 26435
rect 21284 26432 21312 26472
rect 21821 26469 21833 26472
rect 21867 26469 21879 26503
rect 21821 26463 21879 26469
rect 22664 26472 23428 26500
rect 22664 26444 22692 26472
rect 20303 26404 21312 26432
rect 21729 26435 21787 26441
rect 20303 26401 20315 26404
rect 20257 26395 20315 26401
rect 21729 26401 21741 26435
rect 21775 26432 21787 26435
rect 21775 26404 22094 26432
rect 21775 26401 21787 26404
rect 21729 26395 21787 26401
rect 9953 26367 10011 26373
rect 9953 26333 9965 26367
rect 9999 26333 10011 26367
rect 9953 26327 10011 26333
rect 10134 26324 10140 26376
rect 10192 26324 10198 26376
rect 10318 26324 10324 26376
rect 10376 26324 10382 26376
rect 13354 26324 13360 26376
rect 13412 26324 13418 26376
rect 14918 26324 14924 26376
rect 14976 26324 14982 26376
rect 22066 26364 22094 26404
rect 22278 26392 22284 26444
rect 22336 26392 22342 26444
rect 22465 26435 22523 26441
rect 22465 26401 22477 26435
rect 22511 26432 22523 26435
rect 22646 26432 22652 26444
rect 22511 26404 22652 26432
rect 22511 26401 22523 26404
rect 22465 26395 22523 26401
rect 22646 26392 22652 26404
rect 22704 26392 22710 26444
rect 23290 26392 23296 26444
rect 23348 26392 23354 26444
rect 23400 26441 23428 26472
rect 23385 26435 23443 26441
rect 23385 26401 23397 26435
rect 23431 26432 23443 26435
rect 25498 26432 25504 26444
rect 23431 26404 25504 26432
rect 23431 26401 23443 26404
rect 23385 26395 23443 26401
rect 25498 26392 25504 26404
rect 25556 26392 25562 26444
rect 25866 26392 25872 26444
rect 25924 26392 25930 26444
rect 26142 26392 26148 26444
rect 26200 26392 26206 26444
rect 28442 26392 28448 26444
rect 28500 26392 28506 26444
rect 28721 26435 28779 26441
rect 28721 26401 28733 26435
rect 28767 26432 28779 26435
rect 28994 26432 29000 26444
rect 28767 26404 29000 26432
rect 28767 26401 28779 26404
rect 28721 26395 28779 26401
rect 28994 26392 29000 26404
rect 29052 26432 29058 26444
rect 29733 26435 29791 26441
rect 29733 26432 29745 26435
rect 29052 26404 29745 26432
rect 29052 26392 29058 26404
rect 29733 26401 29745 26404
rect 29779 26432 29791 26435
rect 30098 26432 30104 26444
rect 29779 26404 30104 26432
rect 29779 26401 29791 26404
rect 29733 26395 29791 26401
rect 30098 26392 30104 26404
rect 30156 26392 30162 26444
rect 31018 26392 31024 26444
rect 31076 26432 31082 26444
rect 31076 26404 31248 26432
rect 31076 26392 31082 26404
rect 22186 26364 22192 26376
rect 22066 26336 22192 26364
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 22296 26364 22324 26392
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 22296 26336 23213 26364
rect 23201 26333 23213 26336
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 23842 26324 23848 26376
rect 23900 26364 23906 26376
rect 31220 26364 31248 26404
rect 33226 26392 33232 26444
rect 33284 26432 33290 26444
rect 33597 26435 33655 26441
rect 33597 26432 33609 26435
rect 33284 26404 33609 26432
rect 33284 26392 33290 26404
rect 33597 26401 33609 26404
rect 33643 26432 33655 26435
rect 33870 26432 33876 26444
rect 33643 26404 33876 26432
rect 33643 26401 33655 26404
rect 33597 26395 33655 26401
rect 33870 26392 33876 26404
rect 33928 26392 33934 26444
rect 31573 26367 31631 26373
rect 31573 26364 31585 26367
rect 23900 26336 24794 26364
rect 31220 26336 31585 26364
rect 23900 26324 23906 26336
rect 31573 26333 31585 26336
rect 31619 26333 31631 26367
rect 31573 26327 31631 26333
rect 33321 26367 33379 26373
rect 33321 26333 33333 26367
rect 33367 26364 33379 26367
rect 33686 26364 33692 26376
rect 33367 26336 33692 26364
rect 33367 26333 33379 26336
rect 33321 26327 33379 26333
rect 33686 26324 33692 26336
rect 33744 26324 33750 26376
rect 2317 26299 2375 26305
rect 2317 26265 2329 26299
rect 2363 26296 2375 26299
rect 2774 26296 2780 26308
rect 2363 26268 2780 26296
rect 2363 26265 2375 26268
rect 2317 26259 2375 26265
rect 2774 26256 2780 26268
rect 2832 26256 2838 26308
rect 4632 26268 4922 26296
rect 4632 26240 4660 26268
rect 5994 26256 6000 26308
rect 6052 26296 6058 26308
rect 6365 26299 6423 26305
rect 6365 26296 6377 26299
rect 6052 26268 6377 26296
rect 6052 26256 6058 26268
rect 6365 26265 6377 26268
rect 6411 26265 6423 26299
rect 6365 26259 6423 26265
rect 7009 26299 7067 26305
rect 7009 26265 7021 26299
rect 7055 26296 7067 26299
rect 7650 26296 7656 26308
rect 7055 26268 7656 26296
rect 7055 26265 7067 26268
rect 7009 26259 7067 26265
rect 7650 26256 7656 26268
rect 7708 26256 7714 26308
rect 9217 26299 9275 26305
rect 9217 26265 9229 26299
rect 9263 26296 9275 26299
rect 9309 26299 9367 26305
rect 9309 26296 9321 26299
rect 9263 26268 9321 26296
rect 9263 26265 9275 26268
rect 9217 26259 9275 26265
rect 9309 26265 9321 26268
rect 9355 26265 9367 26299
rect 9309 26259 9367 26265
rect 10597 26299 10655 26305
rect 10597 26265 10609 26299
rect 10643 26296 10655 26299
rect 10686 26296 10692 26308
rect 10643 26268 10692 26296
rect 10643 26265 10655 26268
rect 10597 26259 10655 26265
rect 10686 26256 10692 26268
rect 10744 26256 10750 26308
rect 11054 26296 11060 26308
rect 10980 26268 11060 26296
rect 2222 26188 2228 26240
rect 2280 26228 2286 26240
rect 2409 26231 2467 26237
rect 2409 26228 2421 26231
rect 2280 26200 2421 26228
rect 2280 26188 2286 26200
rect 2409 26197 2421 26200
rect 2455 26197 2467 26231
rect 2409 26191 2467 26197
rect 4614 26188 4620 26240
rect 4672 26188 4678 26240
rect 6822 26188 6828 26240
rect 6880 26188 6886 26240
rect 10410 26188 10416 26240
rect 10468 26228 10474 26240
rect 10870 26228 10876 26240
rect 10468 26200 10876 26228
rect 10468 26188 10474 26200
rect 10870 26188 10876 26200
rect 10928 26188 10934 26240
rect 10980 26228 11008 26268
rect 11054 26256 11060 26268
rect 11112 26256 11118 26308
rect 12342 26296 12348 26308
rect 11900 26268 12348 26296
rect 11900 26228 11928 26268
rect 12342 26256 12348 26268
rect 12400 26296 12406 26308
rect 13538 26296 13544 26308
rect 12400 26268 13544 26296
rect 12400 26256 12406 26268
rect 13538 26256 13544 26268
rect 13596 26256 13602 26308
rect 17402 26256 17408 26308
rect 17460 26256 17466 26308
rect 19242 26296 19248 26308
rect 18630 26268 19248 26296
rect 10980 26200 11928 26228
rect 12066 26188 12072 26240
rect 12124 26188 12130 26240
rect 14090 26188 14096 26240
rect 14148 26188 14154 26240
rect 14458 26188 14464 26240
rect 14516 26188 14522 26240
rect 18322 26188 18328 26240
rect 18380 26228 18386 26240
rect 18708 26228 18736 26268
rect 19242 26256 19248 26268
rect 19300 26296 19306 26308
rect 20714 26296 20720 26308
rect 19300 26268 20720 26296
rect 19300 26256 19306 26268
rect 20714 26256 20720 26268
rect 20772 26256 20778 26308
rect 26694 26256 26700 26308
rect 26752 26256 26758 26308
rect 27430 26256 27436 26308
rect 27488 26256 27494 26308
rect 30006 26256 30012 26308
rect 30064 26256 30070 26308
rect 30392 26268 30498 26296
rect 30392 26240 30420 26268
rect 32122 26256 32128 26308
rect 32180 26296 32186 26308
rect 32309 26299 32367 26305
rect 32309 26296 32321 26299
rect 32180 26268 32321 26296
rect 32180 26256 32186 26268
rect 32309 26265 32321 26268
rect 32355 26265 32367 26299
rect 32309 26259 32367 26265
rect 18380 26200 18736 26228
rect 18380 26188 18386 26200
rect 30374 26188 30380 26240
rect 30432 26188 30438 26240
rect 32398 26188 32404 26240
rect 32456 26228 32462 26240
rect 32953 26231 33011 26237
rect 32953 26228 32965 26231
rect 32456 26200 32965 26228
rect 32456 26188 32462 26200
rect 32953 26197 32965 26200
rect 32999 26197 33011 26231
rect 32953 26191 33011 26197
rect 33410 26188 33416 26240
rect 33468 26188 33474 26240
rect 1104 26138 37076 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 37076 26138
rect 1104 26064 37076 26086
rect 3694 25984 3700 26036
rect 3752 25984 3758 26036
rect 4706 25984 4712 26036
rect 4764 25984 4770 26036
rect 9674 25984 9680 26036
rect 9732 25984 9738 26036
rect 10134 25984 10140 26036
rect 10192 26024 10198 26036
rect 10965 26027 11023 26033
rect 10965 26024 10977 26027
rect 10192 25996 10977 26024
rect 10192 25984 10198 25996
rect 10965 25993 10977 25996
rect 11011 25993 11023 26027
rect 10965 25987 11023 25993
rect 14458 25984 14464 26036
rect 14516 26024 14522 26036
rect 14553 26027 14611 26033
rect 14553 26024 14565 26027
rect 14516 25996 14565 26024
rect 14516 25984 14522 25996
rect 14553 25993 14565 25996
rect 14599 25993 14611 26027
rect 14553 25987 14611 25993
rect 17034 25984 17040 26036
rect 17092 25984 17098 26036
rect 17402 25984 17408 26036
rect 17460 25984 17466 26036
rect 18874 26024 18880 26036
rect 17512 25996 18880 26024
rect 2682 25916 2688 25968
rect 2740 25956 2746 25968
rect 3513 25959 3571 25965
rect 3513 25956 3525 25959
rect 2740 25928 3525 25956
rect 2740 25916 2746 25928
rect 3513 25925 3525 25928
rect 3559 25925 3571 25959
rect 3513 25919 3571 25925
rect 3329 25891 3387 25897
rect 3329 25857 3341 25891
rect 3375 25857 3387 25891
rect 3329 25851 3387 25857
rect 2774 25780 2780 25832
rect 2832 25820 2838 25832
rect 3344 25820 3372 25851
rect 3786 25848 3792 25900
rect 3844 25888 3850 25900
rect 4249 25891 4307 25897
rect 4249 25888 4261 25891
rect 3844 25860 4261 25888
rect 3844 25848 3850 25860
rect 4249 25857 4261 25860
rect 4295 25888 4307 25891
rect 4724 25888 4752 25984
rect 6181 25959 6239 25965
rect 6181 25925 6193 25959
rect 6227 25956 6239 25959
rect 7650 25956 7656 25968
rect 6227 25928 7656 25956
rect 6227 25925 6239 25928
rect 6181 25919 6239 25925
rect 7650 25916 7656 25928
rect 7708 25916 7714 25968
rect 8202 25956 8208 25968
rect 7944 25928 8208 25956
rect 4295 25860 4752 25888
rect 4295 25857 4307 25860
rect 4249 25851 4307 25857
rect 6454 25848 6460 25900
rect 6512 25888 6518 25900
rect 6549 25891 6607 25897
rect 6549 25888 6561 25891
rect 6512 25860 6561 25888
rect 6512 25848 6518 25860
rect 6549 25857 6561 25860
rect 6595 25857 6607 25891
rect 6549 25851 6607 25857
rect 7006 25848 7012 25900
rect 7064 25888 7070 25900
rect 7944 25897 7972 25928
rect 8202 25916 8208 25928
rect 8260 25916 8266 25968
rect 8662 25916 8668 25968
rect 8720 25916 8726 25968
rect 7285 25891 7343 25897
rect 7285 25888 7297 25891
rect 7064 25860 7297 25888
rect 7064 25848 7070 25860
rect 7285 25857 7297 25860
rect 7331 25888 7343 25891
rect 7929 25891 7987 25897
rect 7929 25888 7941 25891
rect 7331 25860 7941 25888
rect 7331 25857 7343 25860
rect 7285 25851 7343 25857
rect 7929 25857 7941 25860
rect 7975 25857 7987 25891
rect 9692 25888 9720 25984
rect 10778 25916 10784 25968
rect 10836 25956 10842 25968
rect 10873 25959 10931 25965
rect 10873 25956 10885 25959
rect 10836 25928 10885 25956
rect 10836 25916 10842 25928
rect 10873 25925 10885 25928
rect 10919 25925 10931 25959
rect 10873 25919 10931 25925
rect 13538 25916 13544 25968
rect 13596 25916 13602 25968
rect 10137 25891 10195 25897
rect 10137 25888 10149 25891
rect 9692 25860 10149 25888
rect 7929 25851 7987 25857
rect 10137 25857 10149 25860
rect 10183 25888 10195 25891
rect 10597 25891 10655 25897
rect 10597 25888 10609 25891
rect 10183 25860 10609 25888
rect 10183 25857 10195 25860
rect 10137 25851 10195 25857
rect 10597 25857 10609 25860
rect 10643 25888 10655 25891
rect 11149 25891 11207 25897
rect 10643 25860 11008 25888
rect 10643 25857 10655 25860
rect 10597 25851 10655 25857
rect 4062 25820 4068 25832
rect 2832 25792 4068 25820
rect 2832 25780 2838 25792
rect 4062 25780 4068 25792
rect 4120 25780 4126 25832
rect 5718 25780 5724 25832
rect 5776 25820 5782 25832
rect 6641 25823 6699 25829
rect 6641 25820 6653 25823
rect 5776 25792 6653 25820
rect 5776 25780 5782 25792
rect 6641 25789 6653 25792
rect 6687 25789 6699 25823
rect 6641 25783 6699 25789
rect 6730 25780 6736 25832
rect 6788 25780 6794 25832
rect 6825 25823 6883 25829
rect 6825 25789 6837 25823
rect 6871 25789 6883 25823
rect 6825 25783 6883 25789
rect 8205 25823 8263 25829
rect 8205 25789 8217 25823
rect 8251 25820 8263 25823
rect 9214 25820 9220 25832
rect 8251 25792 9220 25820
rect 8251 25789 8263 25792
rect 8205 25783 8263 25789
rect 6454 25712 6460 25764
rect 6512 25752 6518 25764
rect 6840 25752 6868 25783
rect 9214 25780 9220 25792
rect 9272 25780 9278 25832
rect 9490 25780 9496 25832
rect 9548 25820 9554 25832
rect 9953 25823 10011 25829
rect 9953 25820 9965 25823
rect 9548 25792 9965 25820
rect 9548 25780 9554 25792
rect 9953 25789 9965 25792
rect 9999 25789 10011 25823
rect 9953 25783 10011 25789
rect 10042 25780 10048 25832
rect 10100 25780 10106 25832
rect 10229 25823 10287 25829
rect 10229 25789 10241 25823
rect 10275 25820 10287 25823
rect 10781 25823 10839 25829
rect 10275 25792 10732 25820
rect 10275 25789 10287 25792
rect 10229 25783 10287 25789
rect 6512 25724 6868 25752
rect 9769 25755 9827 25761
rect 6512 25712 6518 25724
rect 9769 25721 9781 25755
rect 9815 25752 9827 25755
rect 10502 25752 10508 25764
rect 9815 25724 10508 25752
rect 9815 25721 9827 25724
rect 9769 25715 9827 25721
rect 10502 25712 10508 25724
rect 10560 25712 10566 25764
rect 10704 25752 10732 25792
rect 10781 25789 10793 25823
rect 10827 25820 10839 25823
rect 10870 25820 10876 25832
rect 10827 25792 10876 25820
rect 10827 25789 10839 25792
rect 10781 25783 10839 25789
rect 10870 25780 10876 25792
rect 10928 25780 10934 25832
rect 10980 25820 11008 25860
rect 11149 25857 11161 25891
rect 11195 25888 11207 25891
rect 12066 25888 12072 25900
rect 11195 25860 12072 25888
rect 11195 25857 11207 25860
rect 11149 25851 11207 25857
rect 11333 25823 11391 25829
rect 11333 25820 11345 25823
rect 10980 25792 11345 25820
rect 11333 25789 11345 25792
rect 11379 25789 11391 25823
rect 11333 25783 11391 25789
rect 10704 25724 10916 25752
rect 5810 25644 5816 25696
rect 5868 25684 5874 25696
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 5868 25656 6377 25684
rect 5868 25644 5874 25656
rect 6365 25653 6377 25656
rect 6411 25653 6423 25687
rect 6365 25647 6423 25653
rect 10042 25644 10048 25696
rect 10100 25684 10106 25696
rect 10888 25693 10916 25724
rect 10413 25687 10471 25693
rect 10413 25684 10425 25687
rect 10100 25656 10425 25684
rect 10100 25644 10106 25656
rect 10413 25653 10425 25656
rect 10459 25653 10471 25687
rect 10413 25647 10471 25653
rect 10873 25687 10931 25693
rect 10873 25653 10885 25687
rect 10919 25684 10931 25687
rect 11440 25684 11468 25860
rect 12066 25848 12072 25860
rect 12124 25848 12130 25900
rect 12802 25848 12808 25900
rect 12860 25848 12866 25900
rect 17512 25888 17540 25996
rect 18874 25984 18880 25996
rect 18932 25984 18938 26036
rect 24946 26024 24952 26036
rect 24412 25996 24952 26024
rect 17954 25916 17960 25968
rect 18012 25916 18018 25968
rect 19242 25956 19248 25968
rect 19182 25928 19248 25956
rect 19242 25916 19248 25928
rect 19300 25916 19306 25968
rect 24412 25965 24440 25996
rect 24946 25984 24952 25996
rect 25004 26024 25010 26036
rect 26142 26024 26148 26036
rect 25004 25996 26148 26024
rect 25004 25984 25010 25996
rect 26142 25984 26148 25996
rect 26200 25984 26206 26036
rect 31478 26024 31484 26036
rect 29380 25996 31484 26024
rect 24397 25959 24455 25965
rect 24397 25925 24409 25959
rect 24443 25925 24455 25959
rect 24397 25919 24455 25925
rect 25774 25916 25780 25968
rect 25832 25916 25838 25968
rect 26510 25956 26516 25968
rect 26206 25928 26516 25956
rect 16868 25860 17540 25888
rect 16868 25832 16896 25860
rect 20346 25848 20352 25900
rect 20404 25888 20410 25900
rect 21453 25891 21511 25897
rect 21453 25888 21465 25891
rect 20404 25860 21465 25888
rect 20404 25848 20410 25860
rect 21453 25857 21465 25860
rect 21499 25857 21511 25891
rect 21453 25851 21511 25857
rect 25317 25891 25375 25897
rect 25317 25857 25329 25891
rect 25363 25857 25375 25891
rect 25317 25851 25375 25857
rect 25409 25891 25467 25897
rect 25409 25857 25421 25891
rect 25455 25888 25467 25891
rect 26206 25888 26234 25928
rect 26510 25916 26516 25928
rect 26568 25916 26574 25968
rect 25455 25860 26234 25888
rect 25455 25857 25467 25860
rect 25409 25851 25467 25857
rect 13081 25823 13139 25829
rect 13081 25789 13093 25823
rect 13127 25820 13139 25823
rect 14090 25820 14096 25832
rect 13127 25792 14096 25820
rect 13127 25789 13139 25792
rect 13081 25783 13139 25789
rect 14090 25780 14096 25792
rect 14148 25780 14154 25832
rect 16850 25780 16856 25832
rect 16908 25780 16914 25832
rect 16942 25780 16948 25832
rect 17000 25780 17006 25832
rect 17681 25823 17739 25829
rect 17681 25789 17693 25823
rect 17727 25820 17739 25823
rect 18506 25820 18512 25832
rect 17727 25792 18512 25820
rect 17727 25789 17739 25792
rect 17681 25783 17739 25789
rect 18506 25780 18512 25792
rect 18564 25780 18570 25832
rect 25332 25820 25360 25851
rect 28074 25848 28080 25900
rect 28132 25848 28138 25900
rect 28258 25848 28264 25900
rect 28316 25848 28322 25900
rect 29380 25897 29408 25996
rect 31478 25984 31484 25996
rect 31536 25984 31542 26036
rect 33686 25984 33692 26036
rect 33744 26024 33750 26036
rect 33873 26027 33931 26033
rect 33873 26024 33885 26027
rect 33744 25996 33885 26024
rect 33744 25984 33750 25996
rect 33873 25993 33885 25996
rect 33919 25993 33931 26027
rect 33873 25987 33931 25993
rect 30006 25916 30012 25968
rect 30064 25956 30070 25968
rect 30101 25959 30159 25965
rect 30101 25956 30113 25959
rect 30064 25928 30113 25956
rect 30064 25916 30070 25928
rect 30101 25925 30113 25928
rect 30147 25925 30159 25959
rect 30101 25919 30159 25925
rect 30374 25916 30380 25968
rect 30432 25956 30438 25968
rect 30432 25928 30958 25956
rect 30432 25916 30438 25928
rect 32398 25916 32404 25968
rect 32456 25916 32462 25968
rect 29365 25891 29423 25897
rect 29365 25857 29377 25891
rect 29411 25857 29423 25891
rect 29365 25851 29423 25857
rect 29457 25891 29515 25897
rect 29457 25857 29469 25891
rect 29503 25857 29515 25891
rect 29457 25851 29515 25857
rect 25332 25792 25452 25820
rect 24949 25755 25007 25761
rect 24949 25721 24961 25755
rect 24995 25752 25007 25755
rect 25130 25752 25136 25764
rect 24995 25724 25136 25752
rect 24995 25721 25007 25724
rect 24949 25715 25007 25721
rect 25130 25712 25136 25724
rect 25188 25712 25194 25764
rect 25424 25752 25452 25792
rect 25498 25780 25504 25832
rect 25556 25780 25562 25832
rect 26234 25780 26240 25832
rect 26292 25820 26298 25832
rect 26513 25823 26571 25829
rect 26513 25820 26525 25823
rect 26292 25792 26525 25820
rect 26292 25780 26298 25792
rect 26513 25789 26525 25792
rect 26559 25820 26571 25823
rect 26694 25820 26700 25832
rect 26559 25792 26700 25820
rect 26559 25789 26571 25792
rect 26513 25783 26571 25789
rect 26694 25780 26700 25792
rect 26752 25780 26758 25832
rect 27617 25823 27675 25829
rect 27617 25789 27629 25823
rect 27663 25820 27675 25823
rect 27798 25820 27804 25832
rect 27663 25792 27804 25820
rect 27663 25789 27675 25792
rect 27617 25783 27675 25789
rect 27798 25780 27804 25792
rect 27856 25780 27862 25832
rect 28350 25780 28356 25832
rect 28408 25780 28414 25832
rect 25958 25752 25964 25764
rect 25424 25724 25964 25752
rect 25958 25712 25964 25724
rect 26016 25712 26022 25764
rect 10919 25656 11468 25684
rect 10919 25653 10931 25656
rect 10873 25647 10931 25653
rect 19426 25644 19432 25696
rect 19484 25684 19490 25696
rect 20990 25684 20996 25696
rect 19484 25656 20996 25684
rect 19484 25644 19490 25656
rect 20990 25644 20996 25656
rect 21048 25644 21054 25696
rect 29472 25684 29500 25851
rect 29638 25848 29644 25900
rect 29696 25848 29702 25900
rect 33502 25848 33508 25900
rect 33560 25888 33566 25900
rect 34054 25888 34060 25900
rect 33560 25860 34060 25888
rect 33560 25848 33566 25860
rect 34054 25848 34060 25860
rect 34112 25848 34118 25900
rect 29546 25780 29552 25832
rect 29604 25820 29610 25832
rect 30190 25820 30196 25832
rect 29604 25792 30196 25820
rect 29604 25780 29610 25792
rect 30190 25780 30196 25792
rect 30248 25780 30254 25832
rect 30469 25823 30527 25829
rect 30469 25789 30481 25823
rect 30515 25820 30527 25823
rect 31110 25820 31116 25832
rect 30515 25792 31116 25820
rect 30515 25789 30527 25792
rect 30469 25783 30527 25789
rect 31110 25780 31116 25792
rect 31168 25780 31174 25832
rect 32122 25780 32128 25832
rect 32180 25780 32186 25832
rect 30650 25684 30656 25696
rect 29472 25656 30656 25684
rect 30650 25644 30656 25656
rect 30708 25644 30714 25696
rect 31754 25644 31760 25696
rect 31812 25684 31818 25696
rect 31941 25687 31999 25693
rect 31941 25684 31953 25687
rect 31812 25656 31953 25684
rect 31812 25644 31818 25656
rect 31941 25653 31953 25656
rect 31987 25653 31999 25687
rect 31941 25647 31999 25653
rect 1104 25594 37076 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 37076 25594
rect 1104 25520 37076 25542
rect 2774 25480 2780 25492
rect 2332 25452 2780 25480
rect 842 25372 848 25424
rect 900 25412 906 25424
rect 1397 25415 1455 25421
rect 1397 25412 1409 25415
rect 900 25384 1409 25412
rect 900 25372 906 25384
rect 1397 25381 1409 25384
rect 1443 25381 1455 25415
rect 1397 25375 1455 25381
rect 2222 25344 2228 25356
rect 1872 25316 2228 25344
rect 1578 25236 1584 25288
rect 1636 25236 1642 25288
rect 1872 25285 1900 25316
rect 2222 25304 2228 25316
rect 2280 25304 2286 25356
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25245 1915 25279
rect 1857 25239 1915 25245
rect 2041 25279 2099 25285
rect 2041 25245 2053 25279
rect 2087 25245 2099 25279
rect 2041 25239 2099 25245
rect 2056 25208 2084 25239
rect 2130 25236 2136 25288
rect 2188 25236 2194 25288
rect 2332 25285 2360 25452
rect 2774 25440 2780 25452
rect 2832 25440 2838 25492
rect 3237 25483 3295 25489
rect 3237 25449 3249 25483
rect 3283 25480 3295 25483
rect 3510 25480 3516 25492
rect 3283 25452 3516 25480
rect 3283 25449 3295 25452
rect 3237 25443 3295 25449
rect 3510 25440 3516 25452
rect 3568 25480 3574 25492
rect 5350 25480 5356 25492
rect 3568 25452 5356 25480
rect 3568 25440 3574 25452
rect 5350 25440 5356 25452
rect 5408 25440 5414 25492
rect 5902 25440 5908 25492
rect 5960 25440 5966 25492
rect 6089 25483 6147 25489
rect 6089 25449 6101 25483
rect 6135 25480 6147 25483
rect 6362 25480 6368 25492
rect 6135 25452 6368 25480
rect 6135 25449 6147 25452
rect 6089 25443 6147 25449
rect 6362 25440 6368 25452
rect 6420 25440 6426 25492
rect 6730 25480 6736 25492
rect 6472 25452 6736 25480
rect 2682 25372 2688 25424
rect 2740 25412 2746 25424
rect 3053 25415 3111 25421
rect 3053 25412 3065 25415
rect 2740 25384 3065 25412
rect 2740 25372 2746 25384
rect 3053 25381 3065 25384
rect 3099 25381 3111 25415
rect 3053 25375 3111 25381
rect 5920 25412 5948 25440
rect 6472 25412 6500 25452
rect 6730 25440 6736 25452
rect 6788 25480 6794 25492
rect 7009 25483 7067 25489
rect 7009 25480 7021 25483
rect 6788 25452 7021 25480
rect 6788 25440 6794 25452
rect 7009 25449 7021 25452
rect 7055 25449 7067 25483
rect 7009 25443 7067 25449
rect 10134 25440 10140 25492
rect 10192 25440 10198 25492
rect 10502 25440 10508 25492
rect 10560 25480 10566 25492
rect 10597 25483 10655 25489
rect 10597 25480 10609 25483
rect 10560 25452 10609 25480
rect 10560 25440 10566 25452
rect 10597 25449 10609 25452
rect 10643 25449 10655 25483
rect 10597 25443 10655 25449
rect 10686 25440 10692 25492
rect 10744 25480 10750 25492
rect 10781 25483 10839 25489
rect 10781 25480 10793 25483
rect 10744 25452 10793 25480
rect 10744 25440 10750 25452
rect 10781 25449 10793 25452
rect 10827 25449 10839 25483
rect 10781 25443 10839 25449
rect 12056 25483 12114 25489
rect 12056 25449 12068 25483
rect 12102 25480 12114 25483
rect 14093 25483 14151 25489
rect 14093 25480 14105 25483
rect 12102 25452 14105 25480
rect 12102 25449 12114 25452
rect 12056 25443 12114 25449
rect 14093 25449 14105 25452
rect 14139 25449 14151 25483
rect 14093 25443 14151 25449
rect 16669 25483 16727 25489
rect 16669 25449 16681 25483
rect 16715 25480 16727 25483
rect 16942 25480 16948 25492
rect 16715 25452 16948 25480
rect 16715 25449 16727 25452
rect 16669 25443 16727 25449
rect 16942 25440 16948 25452
rect 17000 25440 17006 25492
rect 18693 25483 18751 25489
rect 18693 25449 18705 25483
rect 18739 25480 18751 25483
rect 18782 25480 18788 25492
rect 18739 25452 18788 25480
rect 18739 25449 18751 25452
rect 18693 25443 18751 25449
rect 18782 25440 18788 25452
rect 18840 25440 18846 25492
rect 21652 25452 28948 25480
rect 5920 25384 6500 25412
rect 6549 25415 6607 25421
rect 2774 25304 2780 25356
rect 2832 25304 2838 25356
rect 3142 25304 3148 25356
rect 3200 25344 3206 25356
rect 3786 25344 3792 25356
rect 3200 25316 3792 25344
rect 3200 25304 3206 25316
rect 3786 25304 3792 25316
rect 3844 25304 3850 25356
rect 5537 25347 5595 25353
rect 5537 25313 5549 25347
rect 5583 25313 5595 25347
rect 5920 25344 5948 25384
rect 6549 25381 6561 25415
rect 6595 25412 6607 25415
rect 6822 25412 6828 25424
rect 6595 25384 6828 25412
rect 6595 25381 6607 25384
rect 6549 25375 6607 25381
rect 6822 25372 6828 25384
rect 6880 25372 6886 25424
rect 9861 25415 9919 25421
rect 9861 25381 9873 25415
rect 9907 25381 9919 25415
rect 9861 25375 9919 25381
rect 6086 25344 6092 25356
rect 5920 25316 6092 25344
rect 5537 25307 5595 25313
rect 2317 25279 2375 25285
rect 2317 25245 2329 25279
rect 2363 25245 2375 25279
rect 5552 25276 5580 25307
rect 6086 25304 6092 25316
rect 6144 25304 6150 25356
rect 6457 25347 6515 25353
rect 6457 25313 6469 25347
rect 6503 25344 6515 25347
rect 9876 25344 9904 25375
rect 14458 25372 14464 25424
rect 14516 25412 14522 25424
rect 14516 25384 14596 25412
rect 14516 25372 14522 25384
rect 6503 25316 9904 25344
rect 6503 25313 6515 25316
rect 6457 25307 6515 25313
rect 10226 25304 10232 25356
rect 10284 25304 10290 25356
rect 14568 25353 14596 25384
rect 14553 25347 14611 25353
rect 14553 25313 14565 25347
rect 14599 25313 14611 25347
rect 14553 25307 14611 25313
rect 14734 25304 14740 25356
rect 14792 25304 14798 25356
rect 16945 25347 17003 25353
rect 16945 25344 16957 25347
rect 14936 25316 16957 25344
rect 14936 25288 14964 25316
rect 16945 25313 16957 25316
rect 16991 25313 17003 25347
rect 16945 25307 17003 25313
rect 17218 25304 17224 25356
rect 17276 25304 17282 25356
rect 5718 25276 5724 25288
rect 2317 25239 2375 25245
rect 2746 25248 3372 25276
rect 5552 25248 5724 25276
rect 2746 25208 2774 25248
rect 2056 25180 2774 25208
rect 3344 25152 3372 25248
rect 5718 25236 5724 25248
rect 5776 25236 5782 25288
rect 5902 25236 5908 25288
rect 5960 25236 5966 25288
rect 6362 25236 6368 25288
rect 6420 25236 6426 25288
rect 6546 25236 6552 25288
rect 6604 25276 6610 25288
rect 6641 25279 6699 25285
rect 6641 25276 6653 25279
rect 6604 25248 6653 25276
rect 6604 25236 6610 25248
rect 6641 25245 6653 25248
rect 6687 25245 6699 25279
rect 6641 25239 6699 25245
rect 6730 25236 6736 25288
rect 6788 25276 6794 25288
rect 6788 25248 7236 25276
rect 6788 25236 6794 25248
rect 4065 25211 4123 25217
rect 4065 25177 4077 25211
rect 4111 25208 4123 25211
rect 4338 25208 4344 25220
rect 4111 25180 4344 25208
rect 4111 25177 4123 25180
rect 4065 25171 4123 25177
rect 4338 25168 4344 25180
rect 4396 25168 4402 25220
rect 4522 25168 4528 25220
rect 4580 25168 4586 25220
rect 5442 25168 5448 25220
rect 5500 25208 5506 25220
rect 5500 25180 6868 25208
rect 5500 25168 5506 25180
rect 1854 25100 1860 25152
rect 1912 25140 1918 25152
rect 1949 25143 2007 25149
rect 1949 25140 1961 25143
rect 1912 25112 1961 25140
rect 1912 25100 1918 25112
rect 1949 25109 1961 25112
rect 1995 25109 2007 25143
rect 1949 25103 2007 25109
rect 3326 25100 3332 25152
rect 3384 25140 3390 25152
rect 6840 25149 6868 25180
rect 6914 25168 6920 25220
rect 6972 25217 6978 25220
rect 7208 25217 7236 25248
rect 10042 25236 10048 25288
rect 10100 25236 10106 25288
rect 11790 25236 11796 25288
rect 11848 25236 11854 25288
rect 14458 25236 14464 25288
rect 14516 25276 14522 25288
rect 14918 25276 14924 25288
rect 14516 25248 14924 25276
rect 14516 25236 14522 25248
rect 14918 25236 14924 25248
rect 14976 25236 14982 25288
rect 19242 25276 19248 25288
rect 18354 25248 19248 25276
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 20438 25236 20444 25288
rect 20496 25276 20502 25288
rect 21652 25285 21680 25452
rect 21913 25347 21971 25353
rect 21913 25313 21925 25347
rect 21959 25344 21971 25347
rect 22278 25344 22284 25356
rect 21959 25316 22284 25344
rect 21959 25313 21971 25316
rect 21913 25307 21971 25313
rect 22278 25304 22284 25316
rect 22336 25344 22342 25356
rect 22336 25316 22968 25344
rect 22336 25304 22342 25316
rect 20533 25279 20591 25285
rect 20533 25276 20545 25279
rect 20496 25248 20545 25276
rect 20496 25236 20502 25248
rect 20533 25245 20545 25248
rect 20579 25245 20591 25279
rect 20533 25239 20591 25245
rect 21637 25279 21695 25285
rect 21637 25245 21649 25279
rect 21683 25245 21695 25279
rect 21637 25239 21695 25245
rect 21818 25236 21824 25288
rect 21876 25236 21882 25288
rect 22741 25279 22799 25285
rect 22741 25245 22753 25279
rect 22787 25276 22799 25279
rect 22830 25276 22836 25288
rect 22787 25248 22836 25276
rect 22787 25245 22799 25248
rect 22741 25239 22799 25245
rect 22830 25236 22836 25248
rect 22888 25236 22894 25288
rect 22940 25285 22968 25316
rect 24946 25304 24952 25356
rect 25004 25304 25010 25356
rect 28920 25353 28948 25452
rect 28905 25347 28963 25353
rect 28905 25313 28917 25347
rect 28951 25344 28963 25347
rect 29638 25344 29644 25356
rect 28951 25316 29644 25344
rect 28951 25313 28963 25316
rect 28905 25307 28963 25313
rect 29638 25304 29644 25316
rect 29696 25344 29702 25356
rect 30558 25344 30564 25356
rect 29696 25316 30564 25344
rect 29696 25304 29702 25316
rect 30558 25304 30564 25316
rect 30616 25344 30622 25356
rect 30616 25316 32260 25344
rect 30616 25304 30622 25316
rect 22925 25279 22983 25285
rect 22925 25245 22937 25279
rect 22971 25245 22983 25279
rect 22925 25239 22983 25245
rect 23017 25279 23075 25285
rect 23017 25245 23029 25279
rect 23063 25276 23075 25279
rect 23382 25276 23388 25288
rect 23063 25248 23388 25276
rect 23063 25245 23075 25248
rect 23017 25239 23075 25245
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 27430 25276 27436 25288
rect 26358 25248 27436 25276
rect 27430 25236 27436 25248
rect 27488 25236 27494 25288
rect 30009 25279 30067 25285
rect 30009 25245 30021 25279
rect 30055 25276 30067 25279
rect 30055 25248 30144 25276
rect 30055 25245 30067 25248
rect 30009 25239 30067 25245
rect 6972 25211 7035 25217
rect 6972 25177 6989 25211
rect 7023 25177 7035 25211
rect 6972 25171 7035 25177
rect 7193 25211 7251 25217
rect 7193 25177 7205 25211
rect 7239 25177 7251 25211
rect 7193 25171 7251 25177
rect 6972 25168 6978 25171
rect 9950 25168 9956 25220
rect 10008 25208 10014 25220
rect 10321 25211 10379 25217
rect 10321 25208 10333 25211
rect 10008 25180 10333 25208
rect 10008 25168 10014 25180
rect 10321 25177 10333 25180
rect 10367 25177 10379 25211
rect 10321 25171 10379 25177
rect 10413 25211 10471 25217
rect 10413 25177 10425 25211
rect 10459 25177 10471 25211
rect 10413 25171 10471 25177
rect 6181 25143 6239 25149
rect 6181 25140 6193 25143
rect 3384 25112 6193 25140
rect 3384 25100 3390 25112
rect 6181 25109 6193 25112
rect 6227 25109 6239 25143
rect 6181 25103 6239 25109
rect 6825 25143 6883 25149
rect 6825 25109 6837 25143
rect 6871 25109 6883 25143
rect 6825 25103 6883 25109
rect 10226 25100 10232 25152
rect 10284 25140 10290 25152
rect 10428 25140 10456 25171
rect 10594 25168 10600 25220
rect 10652 25217 10658 25220
rect 10652 25211 10671 25217
rect 10659 25177 10671 25211
rect 13814 25208 13820 25220
rect 13294 25180 13820 25208
rect 10652 25171 10671 25177
rect 10652 25168 10658 25171
rect 13814 25168 13820 25180
rect 13872 25168 13878 25220
rect 15194 25168 15200 25220
rect 15252 25168 15258 25220
rect 15838 25168 15844 25220
rect 15896 25168 15902 25220
rect 18506 25168 18512 25220
rect 18564 25208 18570 25220
rect 19705 25211 19763 25217
rect 19705 25208 19717 25211
rect 18564 25180 19717 25208
rect 18564 25168 18570 25180
rect 19705 25177 19717 25180
rect 19751 25208 19763 25211
rect 20346 25208 20352 25220
rect 19751 25180 20352 25208
rect 19751 25177 19763 25180
rect 19705 25171 19763 25177
rect 20346 25168 20352 25180
rect 20404 25168 20410 25220
rect 20806 25168 20812 25220
rect 20864 25208 20870 25220
rect 21177 25211 21235 25217
rect 21177 25208 21189 25211
rect 20864 25180 21189 25208
rect 20864 25168 20870 25180
rect 21177 25177 21189 25180
rect 21223 25177 21235 25211
rect 21177 25171 21235 25177
rect 22094 25168 22100 25220
rect 22152 25208 22158 25220
rect 22281 25211 22339 25217
rect 22281 25208 22293 25211
rect 22152 25180 22293 25208
rect 22152 25168 22158 25180
rect 22281 25177 22293 25180
rect 22327 25177 22339 25211
rect 22281 25171 22339 25177
rect 25222 25168 25228 25220
rect 25280 25168 25286 25220
rect 26602 25168 26608 25220
rect 26660 25208 26666 25220
rect 27157 25211 27215 25217
rect 27157 25208 27169 25211
rect 26660 25180 27169 25208
rect 26660 25168 26666 25180
rect 27157 25177 27169 25180
rect 27203 25208 27215 25211
rect 30116 25208 30144 25248
rect 30190 25236 30196 25288
rect 30248 25276 30254 25288
rect 31113 25279 31171 25285
rect 31113 25276 31125 25279
rect 30248 25248 31125 25276
rect 30248 25236 30254 25248
rect 31113 25245 31125 25248
rect 31159 25276 31171 25279
rect 32122 25276 32128 25288
rect 31159 25248 32128 25276
rect 31159 25245 31171 25248
rect 31113 25239 31171 25245
rect 32122 25236 32128 25248
rect 32180 25236 32186 25288
rect 32232 25276 32260 25316
rect 33410 25304 33416 25356
rect 33468 25344 33474 25356
rect 34057 25347 34115 25353
rect 34057 25344 34069 25347
rect 33468 25316 34069 25344
rect 33468 25304 33474 25316
rect 34057 25313 34069 25316
rect 34103 25344 34115 25347
rect 34422 25344 34428 25356
rect 34103 25316 34428 25344
rect 34103 25313 34115 25316
rect 34057 25307 34115 25313
rect 34422 25304 34428 25316
rect 34480 25304 34486 25356
rect 33778 25276 33784 25288
rect 32232 25248 33784 25276
rect 33778 25236 33784 25248
rect 33836 25236 33842 25288
rect 33965 25279 34023 25285
rect 33965 25245 33977 25279
rect 34011 25245 34023 25279
rect 33965 25239 34023 25245
rect 27203 25180 30144 25208
rect 27203 25177 27215 25180
rect 27157 25171 27215 25177
rect 10284 25112 10456 25140
rect 13541 25143 13599 25149
rect 10284 25100 10290 25112
rect 13541 25109 13553 25143
rect 13587 25140 13599 25143
rect 13998 25140 14004 25152
rect 13587 25112 14004 25140
rect 13587 25109 13599 25112
rect 13541 25103 13599 25109
rect 13998 25100 14004 25112
rect 14056 25140 14062 25152
rect 14461 25143 14519 25149
rect 14461 25140 14473 25143
rect 14056 25112 14473 25140
rect 14056 25100 14062 25112
rect 14461 25109 14473 25112
rect 14507 25109 14519 25143
rect 14461 25103 14519 25109
rect 26697 25143 26755 25149
rect 26697 25109 26709 25143
rect 26743 25140 26755 25143
rect 27430 25140 27436 25152
rect 26743 25112 27436 25140
rect 26743 25109 26755 25112
rect 26697 25103 26755 25109
rect 27430 25100 27436 25112
rect 27488 25100 27494 25152
rect 30116 25140 30144 25180
rect 30466 25168 30472 25220
rect 30524 25208 30530 25220
rect 30653 25211 30711 25217
rect 30653 25208 30665 25211
rect 30524 25180 30665 25208
rect 30524 25168 30530 25180
rect 30653 25177 30665 25180
rect 30699 25208 30711 25211
rect 31386 25208 31392 25220
rect 30699 25180 31392 25208
rect 30699 25177 30711 25180
rect 30653 25171 30711 25177
rect 31386 25168 31392 25180
rect 31444 25168 31450 25220
rect 33318 25168 33324 25220
rect 33376 25168 33382 25220
rect 33980 25208 34008 25239
rect 34514 25208 34520 25220
rect 33980 25180 34520 25208
rect 34514 25168 34520 25180
rect 34572 25168 34578 25220
rect 35434 25140 35440 25152
rect 30116 25112 35440 25140
rect 35434 25100 35440 25112
rect 35492 25100 35498 25152
rect 1104 25050 37076 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 37076 25050
rect 1104 24976 37076 24998
rect 1397 24939 1455 24945
rect 1397 24905 1409 24939
rect 1443 24936 1455 24939
rect 1578 24936 1584 24948
rect 1443 24908 1584 24936
rect 1443 24905 1455 24908
rect 1397 24899 1455 24905
rect 1578 24896 1584 24908
rect 1636 24896 1642 24948
rect 2130 24896 2136 24948
rect 2188 24936 2194 24948
rect 2682 24936 2688 24948
rect 2188 24908 2688 24936
rect 2188 24896 2194 24908
rect 2682 24896 2688 24908
rect 2740 24936 2746 24948
rect 2740 24908 3280 24936
rect 2740 24896 2746 24908
rect 2958 24868 2964 24880
rect 2438 24840 2964 24868
rect 2958 24828 2964 24840
rect 3016 24828 3022 24880
rect 3142 24760 3148 24812
rect 3200 24760 3206 24812
rect 3252 24809 3280 24908
rect 4338 24896 4344 24948
rect 4396 24896 4402 24948
rect 5718 24896 5724 24948
rect 5776 24936 5782 24948
rect 5905 24939 5963 24945
rect 5905 24936 5917 24939
rect 5776 24908 5917 24936
rect 5776 24896 5782 24908
rect 5905 24905 5917 24908
rect 5951 24905 5963 24939
rect 5905 24899 5963 24905
rect 5997 24939 6055 24945
rect 5997 24905 6009 24939
rect 6043 24936 6055 24939
rect 6086 24936 6092 24948
rect 6043 24908 6092 24936
rect 6043 24905 6055 24908
rect 5997 24899 6055 24905
rect 6086 24896 6092 24908
rect 6144 24896 6150 24948
rect 13998 24896 14004 24948
rect 14056 24896 14062 24948
rect 15194 24896 15200 24948
rect 15252 24936 15258 24948
rect 15657 24939 15715 24945
rect 15657 24936 15669 24939
rect 15252 24908 15669 24936
rect 15252 24896 15258 24908
rect 15657 24905 15669 24908
rect 15703 24905 15715 24939
rect 15657 24899 15715 24905
rect 16025 24939 16083 24945
rect 16025 24905 16037 24939
rect 16071 24936 16083 24939
rect 16942 24936 16948 24948
rect 16071 24908 16948 24936
rect 16071 24905 16083 24908
rect 16025 24899 16083 24905
rect 16942 24896 16948 24908
rect 17000 24896 17006 24948
rect 22922 24936 22928 24948
rect 20824 24908 22928 24936
rect 4522 24868 4528 24880
rect 4080 24840 4528 24868
rect 3237 24803 3295 24809
rect 3237 24769 3249 24803
rect 3283 24769 3295 24803
rect 3237 24763 3295 24769
rect 2869 24735 2927 24741
rect 2869 24701 2881 24735
rect 2915 24732 2927 24735
rect 3326 24732 3332 24744
rect 2915 24704 3332 24732
rect 2915 24701 2927 24704
rect 2869 24695 2927 24701
rect 3326 24692 3332 24704
rect 3384 24692 3390 24744
rect 4080 24664 4108 24840
rect 4522 24828 4528 24840
rect 4580 24828 4586 24880
rect 4709 24871 4767 24877
rect 4709 24837 4721 24871
rect 4755 24868 4767 24871
rect 5442 24868 5448 24880
rect 4755 24840 5448 24868
rect 4755 24837 4767 24840
rect 4709 24831 4767 24837
rect 4154 24760 4160 24812
rect 4212 24760 4218 24812
rect 4798 24760 4804 24812
rect 4856 24800 4862 24812
rect 5184 24809 5212 24840
rect 5442 24828 5448 24840
rect 5500 24828 5506 24880
rect 5813 24871 5871 24877
rect 5813 24837 5825 24871
rect 5859 24868 5871 24871
rect 6362 24868 6368 24880
rect 5859 24840 6368 24868
rect 5859 24837 5871 24840
rect 5813 24831 5871 24837
rect 6362 24828 6368 24840
rect 6420 24828 6426 24880
rect 7006 24868 7012 24880
rect 6840 24840 7012 24868
rect 5169 24803 5227 24809
rect 4856 24772 5028 24800
rect 4856 24760 4862 24772
rect 4893 24735 4951 24741
rect 4893 24701 4905 24735
rect 4939 24701 4951 24735
rect 5000 24732 5028 24772
rect 5169 24769 5181 24803
rect 5215 24769 5227 24803
rect 5169 24763 5227 24769
rect 5350 24760 5356 24812
rect 5408 24760 5414 24812
rect 5902 24760 5908 24812
rect 5960 24800 5966 24812
rect 6181 24803 6239 24809
rect 6181 24800 6193 24803
rect 5960 24772 6193 24800
rect 5960 24760 5966 24772
rect 6181 24769 6193 24772
rect 6227 24800 6239 24803
rect 6730 24800 6736 24812
rect 6227 24772 6736 24800
rect 6227 24769 6239 24772
rect 6181 24763 6239 24769
rect 6730 24760 6736 24772
rect 6788 24760 6794 24812
rect 6840 24809 6868 24840
rect 7006 24828 7012 24840
rect 7064 24828 7070 24880
rect 8662 24868 8668 24880
rect 8326 24854 8668 24868
rect 8312 24840 8668 24854
rect 6825 24803 6883 24809
rect 6825 24769 6837 24803
rect 6871 24769 6883 24803
rect 6825 24763 6883 24769
rect 8312 24744 8340 24840
rect 8662 24828 8668 24840
rect 8720 24828 8726 24880
rect 19242 24828 19248 24880
rect 19300 24828 19306 24880
rect 11054 24760 11060 24812
rect 11112 24800 11118 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11112 24772 11713 24800
rect 11112 24760 11118 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 13906 24760 13912 24812
rect 13964 24760 13970 24812
rect 18506 24760 18512 24812
rect 18564 24760 18570 24812
rect 20438 24760 20444 24812
rect 20496 24800 20502 24812
rect 20824 24809 20852 24908
rect 22922 24896 22928 24908
rect 22980 24896 22986 24948
rect 28350 24896 28356 24948
rect 28408 24936 28414 24948
rect 28718 24936 28724 24948
rect 28408 24908 28724 24936
rect 28408 24896 28414 24908
rect 28718 24896 28724 24908
rect 28776 24936 28782 24948
rect 28905 24939 28963 24945
rect 28905 24936 28917 24939
rect 28776 24908 28917 24936
rect 28776 24896 28782 24908
rect 28905 24905 28917 24908
rect 28951 24905 28963 24939
rect 28905 24899 28963 24905
rect 34422 24896 34428 24948
rect 34480 24896 34486 24948
rect 22094 24828 22100 24880
rect 22152 24828 22158 24880
rect 22554 24828 22560 24880
rect 22612 24828 22618 24880
rect 23676 24840 24426 24868
rect 20809 24803 20867 24809
rect 20809 24800 20821 24803
rect 20496 24772 20821 24800
rect 20496 24760 20502 24772
rect 20809 24769 20821 24772
rect 20855 24769 20867 24803
rect 20809 24763 20867 24769
rect 20990 24760 20996 24812
rect 21048 24760 21054 24812
rect 23676 24800 23704 24840
rect 25498 24828 25504 24880
rect 25556 24868 25562 24880
rect 25556 24840 26004 24868
rect 25556 24828 25562 24840
rect 23308 24772 23704 24800
rect 5261 24735 5319 24741
rect 5261 24732 5273 24735
rect 5000 24704 5273 24732
rect 4893 24695 4951 24701
rect 5261 24701 5273 24704
rect 5307 24701 5319 24735
rect 5261 24695 5319 24701
rect 3068 24636 4108 24664
rect 4908 24664 4936 24695
rect 7098 24692 7104 24744
rect 7156 24692 7162 24744
rect 8294 24692 8300 24744
rect 8352 24692 8358 24744
rect 13449 24735 13507 24741
rect 13449 24701 13461 24735
rect 13495 24732 13507 24735
rect 13814 24732 13820 24744
rect 13495 24704 13820 24732
rect 13495 24701 13507 24704
rect 13449 24695 13507 24701
rect 13814 24692 13820 24704
rect 13872 24692 13878 24744
rect 14185 24735 14243 24741
rect 14185 24701 14197 24735
rect 14231 24732 14243 24735
rect 14734 24732 14740 24744
rect 14231 24704 14740 24732
rect 14231 24701 14243 24704
rect 14185 24695 14243 24701
rect 14734 24692 14740 24704
rect 14792 24692 14798 24744
rect 16114 24692 16120 24744
rect 16172 24692 16178 24744
rect 16298 24692 16304 24744
rect 16356 24732 16362 24744
rect 16850 24732 16856 24744
rect 16356 24704 16856 24732
rect 16356 24692 16362 24704
rect 16850 24692 16856 24704
rect 16908 24692 16914 24744
rect 18785 24735 18843 24741
rect 18785 24701 18797 24735
rect 18831 24732 18843 24735
rect 20349 24735 20407 24741
rect 20349 24732 20361 24735
rect 18831 24704 20361 24732
rect 18831 24701 18843 24704
rect 18785 24695 18843 24701
rect 20349 24701 20361 24704
rect 20395 24701 20407 24735
rect 21085 24735 21143 24741
rect 21085 24732 21097 24735
rect 20349 24695 20407 24701
rect 20456 24704 21097 24732
rect 5718 24664 5724 24676
rect 4908 24636 5724 24664
rect 3068 24608 3096 24636
rect 5718 24624 5724 24636
rect 5776 24624 5782 24676
rect 19886 24624 19892 24676
rect 19944 24664 19950 24676
rect 20257 24667 20315 24673
rect 20257 24664 20269 24667
rect 19944 24636 20269 24664
rect 19944 24624 19950 24636
rect 20257 24633 20269 24636
rect 20303 24664 20315 24667
rect 20456 24664 20484 24704
rect 21085 24701 21097 24704
rect 21131 24701 21143 24735
rect 21085 24695 21143 24701
rect 21821 24735 21879 24741
rect 21821 24701 21833 24735
rect 21867 24701 21879 24735
rect 21821 24695 21879 24701
rect 20303 24636 20484 24664
rect 20303 24633 20315 24636
rect 20257 24627 20315 24633
rect 3050 24556 3056 24608
rect 3108 24556 3114 24608
rect 3694 24556 3700 24608
rect 3752 24556 3758 24608
rect 5629 24599 5687 24605
rect 5629 24565 5641 24599
rect 5675 24596 5687 24599
rect 6546 24596 6552 24608
rect 5675 24568 6552 24596
rect 5675 24565 5687 24568
rect 5629 24559 5687 24565
rect 6546 24556 6552 24568
rect 6604 24556 6610 24608
rect 6730 24556 6736 24608
rect 6788 24596 6794 24608
rect 8573 24599 8631 24605
rect 8573 24596 8585 24599
rect 6788 24568 8585 24596
rect 6788 24556 6794 24568
rect 8573 24565 8585 24568
rect 8619 24565 8631 24599
rect 8573 24559 8631 24565
rect 13078 24556 13084 24608
rect 13136 24596 13142 24608
rect 13541 24599 13599 24605
rect 13541 24596 13553 24599
rect 13136 24568 13553 24596
rect 13136 24556 13142 24568
rect 13541 24565 13553 24568
rect 13587 24565 13599 24599
rect 13541 24559 13599 24565
rect 20346 24556 20352 24608
rect 20404 24596 20410 24608
rect 21836 24596 21864 24695
rect 22554 24692 22560 24744
rect 22612 24732 22618 24744
rect 23308 24732 23336 24772
rect 25866 24760 25872 24812
rect 25924 24760 25930 24812
rect 25976 24800 26004 24840
rect 27522 24828 27528 24880
rect 27580 24868 27586 24880
rect 29546 24868 29552 24880
rect 27580 24840 27922 24868
rect 29012 24840 29552 24868
rect 27580 24828 27586 24840
rect 29012 24809 29040 24840
rect 29546 24828 29552 24840
rect 29604 24828 29610 24880
rect 33502 24828 33508 24880
rect 33560 24828 33566 24880
rect 28997 24803 29055 24809
rect 25976 24772 26096 24800
rect 26068 24744 26096 24772
rect 28997 24769 29009 24803
rect 29043 24769 29055 24803
rect 28997 24763 29055 24769
rect 30374 24760 30380 24812
rect 30432 24760 30438 24812
rect 31202 24760 31208 24812
rect 31260 24760 31266 24812
rect 22612 24704 23336 24732
rect 22612 24692 22618 24704
rect 23382 24692 23388 24744
rect 23440 24732 23446 24744
rect 23569 24735 23627 24741
rect 23569 24732 23581 24735
rect 23440 24704 23581 24732
rect 23440 24692 23446 24704
rect 23569 24701 23581 24704
rect 23615 24701 23627 24735
rect 23569 24695 23627 24701
rect 23658 24692 23664 24744
rect 23716 24692 23722 24744
rect 23934 24692 23940 24744
rect 23992 24692 23998 24744
rect 25961 24735 26019 24741
rect 25961 24701 25973 24735
rect 26007 24701 26019 24735
rect 25961 24695 26019 24701
rect 25038 24624 25044 24676
rect 25096 24664 25102 24676
rect 25501 24667 25559 24673
rect 25501 24664 25513 24667
rect 25096 24636 25513 24664
rect 25096 24624 25102 24636
rect 25501 24633 25513 24636
rect 25547 24633 25559 24667
rect 25501 24627 25559 24633
rect 20404 24568 21864 24596
rect 20404 24556 20410 24568
rect 23198 24556 23204 24608
rect 23256 24596 23262 24608
rect 25409 24599 25467 24605
rect 25409 24596 25421 24599
rect 23256 24568 25421 24596
rect 23256 24556 23262 24568
rect 25409 24565 25421 24568
rect 25455 24596 25467 24599
rect 25976 24596 26004 24695
rect 26050 24692 26056 24744
rect 26108 24692 26114 24744
rect 26234 24692 26240 24744
rect 26292 24732 26298 24744
rect 27157 24735 27215 24741
rect 27157 24732 27169 24735
rect 26292 24704 27169 24732
rect 26292 24692 26298 24704
rect 27157 24701 27169 24704
rect 27203 24701 27215 24735
rect 27157 24695 27215 24701
rect 27433 24735 27491 24741
rect 27433 24701 27445 24735
rect 27479 24732 27491 24735
rect 27798 24732 27804 24744
rect 27479 24704 27804 24732
rect 27479 24701 27491 24704
rect 27433 24695 27491 24701
rect 27798 24692 27804 24704
rect 27856 24692 27862 24744
rect 29273 24735 29331 24741
rect 29273 24701 29285 24735
rect 29319 24732 29331 24735
rect 29362 24732 29368 24744
rect 29319 24704 29368 24732
rect 29319 24701 29331 24704
rect 29273 24695 29331 24701
rect 29362 24692 29368 24704
rect 29420 24692 29426 24744
rect 31297 24735 31355 24741
rect 31297 24732 31309 24735
rect 30760 24704 31309 24732
rect 25455 24568 26004 24596
rect 25455 24565 25467 24568
rect 25409 24559 25467 24565
rect 28626 24556 28632 24608
rect 28684 24596 28690 24608
rect 30760 24605 30788 24704
rect 31297 24701 31309 24704
rect 31343 24701 31355 24735
rect 31297 24695 31355 24701
rect 31481 24735 31539 24741
rect 31481 24701 31493 24735
rect 31527 24732 31539 24735
rect 32030 24732 32036 24744
rect 31527 24704 32036 24732
rect 31527 24701 31539 24704
rect 31481 24695 31539 24701
rect 32030 24692 32036 24704
rect 32088 24692 32094 24744
rect 32122 24692 32128 24744
rect 32180 24732 32186 24744
rect 32677 24735 32735 24741
rect 32677 24732 32689 24735
rect 32180 24704 32689 24732
rect 32180 24692 32186 24704
rect 32677 24701 32689 24704
rect 32723 24701 32735 24735
rect 32677 24695 32735 24701
rect 32953 24735 33011 24741
rect 32953 24701 32965 24735
rect 32999 24732 33011 24735
rect 33318 24732 33324 24744
rect 32999 24704 33324 24732
rect 32999 24701 33011 24704
rect 32953 24695 33011 24701
rect 33318 24692 33324 24704
rect 33376 24692 33382 24744
rect 30745 24599 30803 24605
rect 30745 24596 30757 24599
rect 28684 24568 30757 24596
rect 28684 24556 28690 24568
rect 30745 24565 30757 24568
rect 30791 24565 30803 24599
rect 30745 24559 30803 24565
rect 30834 24556 30840 24608
rect 30892 24556 30898 24608
rect 1104 24506 37076 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 37076 24506
rect 1104 24432 37076 24454
rect 7098 24352 7104 24404
rect 7156 24392 7162 24404
rect 7377 24395 7435 24401
rect 7377 24392 7389 24395
rect 7156 24364 7389 24392
rect 7156 24352 7162 24364
rect 7377 24361 7389 24364
rect 7423 24361 7435 24395
rect 7377 24355 7435 24361
rect 13906 24352 13912 24404
rect 13964 24352 13970 24404
rect 16114 24352 16120 24404
rect 16172 24392 16178 24404
rect 16209 24395 16267 24401
rect 16209 24392 16221 24395
rect 16172 24364 16221 24392
rect 16172 24352 16178 24364
rect 16209 24361 16221 24364
rect 16255 24361 16267 24395
rect 16209 24355 16267 24361
rect 22278 24352 22284 24404
rect 22336 24352 22342 24404
rect 25866 24352 25872 24404
rect 25924 24392 25930 24404
rect 26145 24395 26203 24401
rect 26145 24392 26157 24395
rect 25924 24364 26157 24392
rect 25924 24352 25930 24364
rect 26145 24361 26157 24364
rect 26191 24361 26203 24395
rect 26145 24355 26203 24361
rect 27985 24395 28043 24401
rect 27985 24361 27997 24395
rect 28031 24392 28043 24395
rect 28258 24392 28264 24404
rect 28031 24364 28264 24392
rect 28031 24361 28043 24364
rect 27985 24355 28043 24361
rect 28258 24352 28264 24364
rect 28316 24352 28322 24404
rect 31202 24352 31208 24404
rect 31260 24392 31266 24404
rect 31297 24395 31355 24401
rect 31297 24392 31309 24395
rect 31260 24364 31309 24392
rect 31260 24352 31266 24364
rect 31297 24361 31309 24364
rect 31343 24392 31355 24395
rect 31343 24364 31892 24392
rect 31343 24361 31355 24364
rect 31297 24355 31355 24361
rect 7469 24327 7527 24333
rect 7469 24293 7481 24327
rect 7515 24293 7527 24327
rect 20438 24324 20444 24336
rect 7469 24287 7527 24293
rect 19720 24296 20444 24324
rect 1581 24259 1639 24265
rect 1581 24225 1593 24259
rect 1627 24256 1639 24259
rect 3142 24256 3148 24268
rect 1627 24228 3148 24256
rect 1627 24225 1639 24228
rect 1581 24219 1639 24225
rect 3142 24216 3148 24228
rect 3200 24216 3206 24268
rect 3605 24259 3663 24265
rect 3605 24225 3617 24259
rect 3651 24256 3663 24259
rect 4062 24256 4068 24268
rect 3651 24228 4068 24256
rect 3651 24225 3663 24228
rect 3605 24219 3663 24225
rect 4062 24216 4068 24228
rect 4120 24216 4126 24268
rect 2958 24148 2964 24200
rect 3016 24148 3022 24200
rect 6914 24148 6920 24200
rect 6972 24188 6978 24200
rect 7101 24191 7159 24197
rect 7101 24188 7113 24191
rect 6972 24160 7113 24188
rect 6972 24148 6978 24160
rect 7101 24157 7113 24160
rect 7147 24188 7159 24191
rect 7377 24191 7435 24197
rect 7147 24160 7328 24188
rect 7147 24157 7159 24160
rect 7101 24151 7159 24157
rect 1854 24080 1860 24132
rect 1912 24080 1918 24132
rect 6730 24080 6736 24132
rect 6788 24120 6794 24132
rect 7193 24123 7251 24129
rect 7193 24120 7205 24123
rect 6788 24092 7205 24120
rect 6788 24080 6794 24092
rect 7193 24089 7205 24092
rect 7239 24089 7251 24123
rect 7300 24120 7328 24160
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 7484 24188 7512 24287
rect 11790 24216 11796 24268
rect 11848 24256 11854 24268
rect 12158 24256 12164 24268
rect 11848 24228 12164 24256
rect 11848 24216 11854 24228
rect 12158 24216 12164 24228
rect 12216 24216 12222 24268
rect 12437 24259 12495 24265
rect 12437 24225 12449 24259
rect 12483 24256 12495 24259
rect 13078 24256 13084 24268
rect 12483 24228 13084 24256
rect 12483 24225 12495 24228
rect 12437 24219 12495 24225
rect 13078 24216 13084 24228
rect 13136 24216 13142 24268
rect 18141 24259 18199 24265
rect 18141 24225 18153 24259
rect 18187 24256 18199 24259
rect 18506 24256 18512 24268
rect 18187 24228 18512 24256
rect 18187 24225 18199 24228
rect 18141 24219 18199 24225
rect 18506 24216 18512 24228
rect 18564 24216 18570 24268
rect 7423 24160 7512 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 7742 24148 7748 24200
rect 7800 24148 7806 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 15838 24148 15844 24200
rect 15896 24188 15902 24200
rect 19720 24197 19748 24296
rect 20438 24284 20444 24296
rect 20496 24284 20502 24336
rect 31110 24284 31116 24336
rect 31168 24324 31174 24336
rect 31389 24327 31447 24333
rect 31389 24324 31401 24327
rect 31168 24296 31401 24324
rect 31168 24284 31174 24296
rect 31389 24293 31401 24296
rect 31435 24293 31447 24327
rect 31389 24287 31447 24293
rect 20346 24216 20352 24268
rect 20404 24256 20410 24268
rect 20533 24259 20591 24265
rect 20533 24256 20545 24259
rect 20404 24228 20545 24256
rect 20404 24216 20410 24228
rect 20533 24225 20545 24228
rect 20579 24225 20591 24259
rect 20533 24219 20591 24225
rect 20806 24216 20812 24268
rect 20864 24216 20870 24268
rect 23658 24216 23664 24268
rect 23716 24256 23722 24268
rect 24397 24259 24455 24265
rect 24397 24256 24409 24259
rect 23716 24228 24409 24256
rect 23716 24216 23722 24228
rect 24397 24225 24409 24228
rect 24443 24225 24455 24259
rect 24397 24219 24455 24225
rect 24673 24259 24731 24265
rect 24673 24225 24685 24259
rect 24719 24256 24731 24259
rect 25038 24256 25044 24268
rect 24719 24228 25044 24256
rect 24719 24225 24731 24228
rect 24673 24219 24731 24225
rect 25038 24216 25044 24228
rect 25096 24216 25102 24268
rect 28626 24216 28632 24268
rect 28684 24216 28690 24268
rect 29362 24216 29368 24268
rect 29420 24216 29426 24268
rect 29825 24259 29883 24265
rect 29825 24225 29837 24259
rect 29871 24256 29883 24259
rect 30834 24256 30840 24268
rect 29871 24228 30840 24256
rect 29871 24225 29883 24228
rect 29825 24219 29883 24225
rect 30834 24216 30840 24228
rect 30892 24216 30898 24268
rect 31864 24265 31892 24364
rect 34514 24352 34520 24404
rect 34572 24352 34578 24404
rect 31849 24259 31907 24265
rect 31849 24225 31861 24259
rect 31895 24225 31907 24259
rect 31849 24219 31907 24225
rect 32030 24216 32036 24268
rect 32088 24216 32094 24268
rect 32122 24216 32128 24268
rect 32180 24256 32186 24268
rect 32769 24259 32827 24265
rect 32769 24256 32781 24259
rect 32180 24228 32781 24256
rect 32180 24216 32186 24228
rect 32769 24225 32781 24228
rect 32815 24225 32827 24259
rect 32769 24219 32827 24225
rect 19705 24191 19763 24197
rect 15896 24160 16790 24188
rect 15896 24148 15902 24160
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 19886 24148 19892 24200
rect 19944 24148 19950 24200
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24188 20039 24191
rect 20070 24188 20076 24200
rect 20027 24160 20076 24188
rect 20027 24157 20039 24160
rect 19981 24151 20039 24157
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 22554 24188 22560 24200
rect 21942 24160 22560 24188
rect 22554 24148 22560 24160
rect 22612 24188 22618 24200
rect 22612 24160 24256 24188
rect 22612 24148 22618 24160
rect 7469 24123 7527 24129
rect 7469 24120 7481 24123
rect 7300 24092 7481 24120
rect 7193 24083 7251 24089
rect 7469 24089 7481 24092
rect 7515 24089 7527 24123
rect 13814 24120 13820 24132
rect 13662 24092 13820 24120
rect 7469 24083 7527 24089
rect 7208 24052 7236 24083
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 14734 24080 14740 24132
rect 14792 24080 14798 24132
rect 17770 24080 17776 24132
rect 17828 24120 17834 24132
rect 17865 24123 17923 24129
rect 17865 24120 17877 24123
rect 17828 24092 17877 24120
rect 17828 24080 17834 24092
rect 17865 24089 17877 24092
rect 17911 24089 17923 24123
rect 17865 24083 17923 24089
rect 19245 24123 19303 24129
rect 19245 24089 19257 24123
rect 19291 24120 19303 24123
rect 19291 24092 20024 24120
rect 19291 24089 19303 24092
rect 19245 24083 19303 24089
rect 19996 24064 20024 24092
rect 24118 24080 24124 24132
rect 24176 24080 24182 24132
rect 24228 24120 24256 24160
rect 26234 24148 26240 24200
rect 26292 24148 26298 24200
rect 27522 24148 27528 24200
rect 27580 24188 27586 24200
rect 27580 24174 27646 24188
rect 27580 24160 27660 24174
rect 27580 24148 27586 24160
rect 24228 24092 25162 24120
rect 7653 24055 7711 24061
rect 7653 24052 7665 24055
rect 7208 24024 7665 24052
rect 7653 24021 7665 24024
rect 7699 24021 7711 24055
rect 7653 24015 7711 24021
rect 16390 24012 16396 24064
rect 16448 24012 16454 24064
rect 19978 24012 19984 24064
rect 20036 24012 20042 24064
rect 22833 24055 22891 24061
rect 22833 24021 22845 24055
rect 22879 24052 22891 24055
rect 22922 24052 22928 24064
rect 22879 24024 22928 24052
rect 22879 24021 22891 24024
rect 22833 24015 22891 24021
rect 22922 24012 22928 24024
rect 22980 24012 22986 24064
rect 25056 24052 25084 24092
rect 26510 24080 26516 24132
rect 26568 24080 26574 24132
rect 27632 24052 27660 24160
rect 28718 24148 28724 24200
rect 28776 24148 28782 24200
rect 28902 24148 28908 24200
rect 28960 24148 28966 24200
rect 29546 24148 29552 24200
rect 29604 24148 29610 24200
rect 31754 24148 31760 24200
rect 31812 24148 31818 24200
rect 32048 24188 32076 24216
rect 32048 24160 32168 24188
rect 30374 24080 30380 24132
rect 30432 24080 30438 24132
rect 25056 24024 27660 24052
rect 32140 24052 32168 24160
rect 33042 24080 33048 24132
rect 33100 24080 33106 24132
rect 33502 24080 33508 24132
rect 33560 24080 33566 24132
rect 33226 24052 33232 24064
rect 32140 24024 33232 24052
rect 33226 24012 33232 24024
rect 33284 24052 33290 24064
rect 34054 24052 34060 24064
rect 33284 24024 34060 24052
rect 33284 24012 33290 24024
rect 34054 24012 34060 24024
rect 34112 24012 34118 24064
rect 1104 23962 37076 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 37076 23962
rect 1104 23888 37076 23910
rect 5626 23848 5632 23860
rect 5000 23820 5632 23848
rect 3694 23740 3700 23792
rect 3752 23780 3758 23792
rect 5000 23789 5028 23820
rect 5626 23808 5632 23820
rect 5684 23848 5690 23860
rect 7742 23848 7748 23860
rect 5684 23820 7748 23848
rect 5684 23808 5690 23820
rect 7742 23808 7748 23820
rect 7800 23848 7806 23860
rect 7800 23820 9444 23848
rect 7800 23808 7806 23820
rect 4985 23783 5043 23789
rect 4985 23780 4997 23783
rect 3752 23752 4997 23780
rect 3752 23740 3758 23752
rect 4985 23749 4997 23752
rect 5031 23749 5043 23783
rect 4985 23743 5043 23749
rect 5074 23740 5080 23792
rect 5132 23780 5138 23792
rect 5185 23783 5243 23789
rect 5185 23780 5197 23783
rect 5132 23752 5197 23780
rect 5132 23740 5138 23752
rect 5185 23749 5197 23752
rect 5231 23749 5243 23783
rect 5185 23743 5243 23749
rect 5350 23740 5356 23792
rect 5408 23780 5414 23792
rect 9125 23783 9183 23789
rect 5408 23752 8064 23780
rect 5408 23740 5414 23752
rect 8036 23724 8064 23752
rect 9125 23749 9137 23783
rect 9171 23749 9183 23783
rect 9125 23743 9183 23749
rect 842 23672 848 23724
rect 900 23712 906 23724
rect 1397 23715 1455 23721
rect 1397 23712 1409 23715
rect 900 23684 1409 23712
rect 900 23672 906 23684
rect 1397 23681 1409 23684
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 2130 23712 2136 23724
rect 1719 23684 2136 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 2130 23672 2136 23684
rect 2188 23672 2194 23724
rect 6546 23672 6552 23724
rect 6604 23672 6610 23724
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23712 6791 23715
rect 6914 23712 6920 23724
rect 6779 23684 6920 23712
rect 6779 23681 6791 23684
rect 6733 23675 6791 23681
rect 6914 23672 6920 23684
rect 6972 23672 6978 23724
rect 8018 23672 8024 23724
rect 8076 23712 8082 23724
rect 8205 23715 8263 23721
rect 8205 23712 8217 23715
rect 8076 23684 8217 23712
rect 8076 23672 8082 23684
rect 8205 23681 8217 23684
rect 8251 23681 8263 23715
rect 8205 23675 8263 23681
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23712 8447 23715
rect 8570 23712 8576 23724
rect 8435 23684 8576 23712
rect 8435 23681 8447 23684
rect 8389 23675 8447 23681
rect 8570 23672 8576 23684
rect 8628 23712 8634 23724
rect 8665 23715 8723 23721
rect 8665 23712 8677 23715
rect 8628 23684 8677 23712
rect 8628 23672 8634 23684
rect 8665 23681 8677 23684
rect 8711 23681 8723 23715
rect 8665 23675 8723 23681
rect 8754 23672 8760 23724
rect 8812 23712 8818 23724
rect 9140 23712 9168 23743
rect 9214 23740 9220 23792
rect 9272 23780 9278 23792
rect 9325 23783 9383 23789
rect 9325 23780 9337 23783
rect 9272 23752 9337 23780
rect 9272 23740 9278 23752
rect 9325 23749 9337 23752
rect 9371 23749 9383 23783
rect 9416 23780 9444 23820
rect 9490 23808 9496 23860
rect 9548 23808 9554 23860
rect 10134 23808 10140 23860
rect 10192 23808 10198 23860
rect 10686 23848 10692 23860
rect 10244 23820 10692 23848
rect 10244 23792 10272 23820
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 13541 23851 13599 23857
rect 13541 23817 13553 23851
rect 13587 23848 13599 23851
rect 13906 23848 13912 23860
rect 13587 23820 13912 23848
rect 13587 23817 13599 23820
rect 13541 23811 13599 23817
rect 13906 23808 13912 23820
rect 13964 23808 13970 23860
rect 14734 23808 14740 23860
rect 14792 23848 14798 23860
rect 15473 23851 15531 23857
rect 15473 23848 15485 23851
rect 14792 23820 15485 23848
rect 14792 23808 14798 23820
rect 15473 23817 15485 23820
rect 15519 23817 15531 23851
rect 15473 23811 15531 23817
rect 15841 23851 15899 23857
rect 15841 23817 15853 23851
rect 15887 23848 15899 23851
rect 16114 23848 16120 23860
rect 15887 23820 16120 23848
rect 15887 23817 15899 23820
rect 15841 23811 15899 23817
rect 16114 23808 16120 23820
rect 16172 23808 16178 23860
rect 17770 23808 17776 23860
rect 17828 23808 17834 23860
rect 18509 23851 18567 23857
rect 18509 23817 18521 23851
rect 18555 23848 18567 23851
rect 18690 23848 18696 23860
rect 18555 23820 18696 23848
rect 18555 23817 18567 23820
rect 18509 23811 18567 23817
rect 18690 23808 18696 23820
rect 18748 23848 18754 23860
rect 20070 23848 20076 23860
rect 18748 23820 20076 23848
rect 18748 23808 18754 23820
rect 20070 23808 20076 23820
rect 20128 23808 20134 23860
rect 25222 23808 25228 23860
rect 25280 23848 25286 23860
rect 25317 23851 25375 23857
rect 25317 23848 25329 23851
rect 25280 23820 25329 23848
rect 25280 23808 25286 23820
rect 25317 23817 25329 23820
rect 25363 23817 25375 23851
rect 25317 23811 25375 23817
rect 25777 23851 25835 23857
rect 25777 23817 25789 23851
rect 25823 23848 25835 23851
rect 25866 23848 25872 23860
rect 25823 23820 25872 23848
rect 25823 23817 25835 23820
rect 25777 23811 25835 23817
rect 25866 23808 25872 23820
rect 25924 23808 25930 23860
rect 26510 23808 26516 23860
rect 26568 23848 26574 23860
rect 26973 23851 27031 23857
rect 26973 23848 26985 23851
rect 26568 23820 26985 23848
rect 26568 23808 26574 23820
rect 26973 23817 26985 23820
rect 27019 23817 27031 23851
rect 26973 23811 27031 23817
rect 27341 23851 27399 23857
rect 27341 23817 27353 23851
rect 27387 23848 27399 23851
rect 28258 23848 28264 23860
rect 27387 23820 28264 23848
rect 27387 23817 27399 23820
rect 27341 23811 27399 23817
rect 28258 23808 28264 23820
rect 28316 23808 28322 23860
rect 33042 23808 33048 23860
rect 33100 23848 33106 23860
rect 34333 23851 34391 23857
rect 34333 23848 34345 23851
rect 33100 23820 34345 23848
rect 33100 23808 33106 23820
rect 34333 23817 34345 23820
rect 34379 23817 34391 23851
rect 34333 23811 34391 23817
rect 34514 23808 34520 23860
rect 34572 23848 34578 23860
rect 34701 23851 34759 23857
rect 34701 23848 34713 23851
rect 34572 23820 34713 23848
rect 34572 23808 34578 23820
rect 34701 23817 34713 23820
rect 34747 23817 34759 23851
rect 34701 23811 34759 23817
rect 10226 23780 10232 23792
rect 9416 23752 10232 23780
rect 9325 23743 9383 23749
rect 10226 23740 10232 23752
rect 10284 23740 10290 23792
rect 15933 23783 15991 23789
rect 10459 23749 10517 23755
rect 10459 23746 10471 23749
rect 9677 23715 9735 23721
rect 9677 23712 9689 23715
rect 8812 23684 9689 23712
rect 8812 23672 8818 23684
rect 9677 23681 9689 23684
rect 9723 23681 9735 23715
rect 9677 23675 9735 23681
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 9953 23715 10011 23721
rect 9953 23712 9965 23715
rect 9824 23684 9965 23712
rect 9824 23672 9830 23684
rect 9953 23681 9965 23684
rect 9999 23681 10011 23715
rect 10444 23715 10471 23746
rect 10505 23724 10517 23749
rect 15933 23749 15945 23783
rect 15979 23780 15991 23783
rect 16390 23780 16396 23792
rect 15979 23752 16396 23780
rect 15979 23749 15991 23752
rect 15933 23743 15991 23749
rect 16390 23740 16396 23752
rect 16448 23780 16454 23792
rect 17405 23783 17463 23789
rect 17405 23780 17417 23783
rect 16448 23752 17417 23780
rect 16448 23740 16454 23752
rect 17405 23749 17417 23752
rect 17451 23749 17463 23783
rect 17405 23743 17463 23749
rect 19242 23740 19248 23792
rect 19300 23740 19306 23792
rect 19978 23740 19984 23792
rect 20036 23740 20042 23792
rect 23934 23740 23940 23792
rect 23992 23740 23998 23792
rect 25685 23783 25743 23789
rect 25685 23749 25697 23783
rect 25731 23780 25743 23783
rect 27430 23780 27436 23792
rect 25731 23752 27436 23780
rect 25731 23749 25743 23752
rect 25685 23743 25743 23749
rect 27430 23740 27436 23752
rect 27488 23740 27494 23792
rect 30466 23740 30472 23792
rect 30524 23780 30530 23792
rect 30524 23752 30880 23780
rect 30524 23740 30530 23752
rect 10505 23715 10508 23724
rect 10444 23684 10508 23715
rect 9953 23675 10011 23681
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 13906 23712 13912 23724
rect 13495 23684 13912 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 20257 23715 20315 23721
rect 20257 23681 20269 23715
rect 20303 23712 20315 23715
rect 20346 23712 20352 23724
rect 20303 23684 20352 23712
rect 20303 23681 20315 23684
rect 20257 23675 20315 23681
rect 9861 23647 9919 23653
rect 9861 23613 9873 23647
rect 9907 23644 9919 23647
rect 10870 23644 10876 23656
rect 9907 23616 10876 23644
rect 9907 23613 9919 23616
rect 9861 23607 9919 23613
rect 10870 23604 10876 23616
rect 10928 23604 10934 23656
rect 13725 23647 13783 23653
rect 13725 23613 13737 23647
rect 13771 23644 13783 23647
rect 15378 23644 15384 23656
rect 13771 23616 15384 23644
rect 13771 23613 13783 23616
rect 13725 23607 13783 23613
rect 15378 23604 15384 23616
rect 15436 23644 15442 23656
rect 16117 23647 16175 23653
rect 16117 23644 16129 23647
rect 15436 23616 16129 23644
rect 15436 23604 15442 23616
rect 16117 23613 16129 23616
rect 16163 23644 16175 23647
rect 16298 23644 16304 23656
rect 16163 23616 16304 23644
rect 16163 23613 16175 23616
rect 16117 23607 16175 23613
rect 16298 23604 16304 23616
rect 16356 23644 16362 23656
rect 17126 23644 17132 23656
rect 16356 23616 17132 23644
rect 16356 23604 16362 23616
rect 17126 23604 17132 23616
rect 17184 23604 17190 23656
rect 17310 23604 17316 23656
rect 17368 23604 17374 23656
rect 19610 23604 19616 23656
rect 19668 23644 19674 23656
rect 20272 23644 20300 23675
rect 20346 23672 20352 23684
rect 20404 23672 20410 23724
rect 23198 23672 23204 23724
rect 23256 23672 23262 23724
rect 23293 23715 23351 23721
rect 23293 23681 23305 23715
rect 23339 23712 23351 23715
rect 23382 23712 23388 23724
rect 23339 23684 23388 23712
rect 23339 23681 23351 23684
rect 23293 23675 23351 23681
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 23474 23672 23480 23724
rect 23532 23672 23538 23724
rect 24118 23672 24124 23724
rect 24176 23712 24182 23724
rect 25041 23715 25099 23721
rect 25041 23712 25053 23715
rect 24176 23684 25053 23712
rect 24176 23672 24182 23684
rect 25041 23681 25053 23684
rect 25087 23712 25099 23715
rect 26510 23712 26516 23724
rect 25087 23684 26516 23712
rect 25087 23681 25099 23684
rect 25041 23675 25099 23681
rect 26510 23672 26516 23684
rect 26568 23672 26574 23724
rect 30558 23672 30564 23724
rect 30616 23672 30622 23724
rect 30742 23672 30748 23724
rect 30800 23672 30806 23724
rect 30852 23712 30880 23752
rect 31754 23740 31760 23792
rect 31812 23780 31818 23792
rect 31812 23752 32812 23780
rect 31812 23740 31818 23752
rect 32784 23721 32812 23752
rect 32876 23752 33916 23780
rect 32876 23721 32904 23752
rect 33888 23724 33916 23752
rect 32585 23715 32643 23721
rect 32585 23712 32597 23715
rect 30852 23684 32597 23712
rect 32585 23681 32597 23684
rect 32631 23681 32643 23715
rect 32585 23675 32643 23681
rect 32769 23715 32827 23721
rect 32769 23681 32781 23715
rect 32815 23681 32827 23715
rect 32769 23675 32827 23681
rect 32861 23715 32919 23721
rect 32861 23681 32873 23715
rect 32907 23681 32919 23715
rect 33689 23715 33747 23721
rect 33689 23712 33701 23715
rect 32861 23675 32919 23681
rect 32968 23684 33701 23712
rect 19668 23616 20300 23644
rect 23492 23644 23520 23672
rect 23750 23644 23756 23656
rect 23492 23616 23756 23644
rect 19668 23604 19674 23616
rect 23750 23604 23756 23616
rect 23808 23644 23814 23656
rect 24213 23647 24271 23653
rect 24213 23644 24225 23647
rect 23808 23616 24225 23644
rect 23808 23604 23814 23616
rect 24213 23613 24225 23616
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 25961 23647 26019 23653
rect 25961 23613 25973 23647
rect 26007 23644 26019 23647
rect 26050 23644 26056 23656
rect 26007 23616 26056 23644
rect 26007 23613 26019 23616
rect 25961 23607 26019 23613
rect 5810 23576 5816 23588
rect 5184 23548 5816 23576
rect 5184 23517 5212 23548
rect 5810 23536 5816 23548
rect 5868 23536 5874 23588
rect 24228 23576 24256 23607
rect 26050 23604 26056 23616
rect 26108 23644 26114 23656
rect 27522 23644 27528 23656
rect 26108 23616 27528 23644
rect 26108 23604 26114 23616
rect 27522 23604 27528 23616
rect 27580 23604 27586 23656
rect 30101 23647 30159 23653
rect 30101 23613 30113 23647
rect 30147 23644 30159 23647
rect 30190 23644 30196 23656
rect 30147 23616 30196 23644
rect 30147 23613 30159 23616
rect 30101 23607 30159 23613
rect 30190 23604 30196 23616
rect 30248 23604 30254 23656
rect 30650 23604 30656 23656
rect 30708 23644 30714 23656
rect 30837 23647 30895 23653
rect 30837 23644 30849 23647
rect 30708 23616 30849 23644
rect 30708 23604 30714 23616
rect 30837 23613 30849 23616
rect 30883 23613 30895 23647
rect 30837 23607 30895 23613
rect 32125 23647 32183 23653
rect 32125 23613 32137 23647
rect 32171 23644 32183 23647
rect 32398 23644 32404 23656
rect 32171 23616 32404 23644
rect 32171 23613 32183 23616
rect 32125 23607 32183 23613
rect 32398 23604 32404 23616
rect 32456 23604 32462 23656
rect 32600 23644 32628 23675
rect 32968 23644 32996 23684
rect 33689 23681 33701 23684
rect 33735 23681 33747 23715
rect 33689 23675 33747 23681
rect 33870 23672 33876 23724
rect 33928 23672 33934 23724
rect 34054 23672 34060 23724
rect 34112 23712 34118 23724
rect 34112 23684 34928 23712
rect 34112 23672 34118 23684
rect 32600 23616 32996 23644
rect 33226 23604 33232 23656
rect 33284 23604 33290 23656
rect 33965 23647 34023 23653
rect 33965 23613 33977 23647
rect 34011 23644 34023 23647
rect 34422 23644 34428 23656
rect 34011 23616 34428 23644
rect 34011 23613 34023 23616
rect 33965 23607 34023 23613
rect 34422 23604 34428 23616
rect 34480 23644 34486 23656
rect 34900 23653 34928 23684
rect 34793 23647 34851 23653
rect 34793 23644 34805 23647
rect 34480 23616 34805 23644
rect 34480 23604 34486 23616
rect 34793 23613 34805 23616
rect 34839 23613 34851 23647
rect 34793 23607 34851 23613
rect 34885 23647 34943 23653
rect 34885 23613 34897 23647
rect 34931 23613 34943 23647
rect 34885 23607 34943 23613
rect 27614 23576 27620 23588
rect 24228 23548 27620 23576
rect 27614 23536 27620 23548
rect 27672 23576 27678 23588
rect 28074 23576 28080 23588
rect 27672 23548 28080 23576
rect 27672 23536 27678 23548
rect 28074 23536 28080 23548
rect 28132 23576 28138 23588
rect 28902 23576 28908 23588
rect 28132 23548 28908 23576
rect 28132 23536 28138 23548
rect 28902 23536 28908 23548
rect 28960 23536 28966 23588
rect 5169 23511 5227 23517
rect 5169 23477 5181 23511
rect 5215 23477 5227 23511
rect 5169 23471 5227 23477
rect 5258 23468 5264 23520
rect 5316 23508 5322 23520
rect 5353 23511 5411 23517
rect 5353 23508 5365 23511
rect 5316 23480 5365 23508
rect 5316 23468 5322 23480
rect 5353 23477 5365 23480
rect 5399 23477 5411 23511
rect 5353 23471 5411 23477
rect 5534 23468 5540 23520
rect 5592 23508 5598 23520
rect 6178 23508 6184 23520
rect 5592 23480 6184 23508
rect 5592 23468 5598 23480
rect 6178 23468 6184 23480
rect 6236 23508 6242 23520
rect 6365 23511 6423 23517
rect 6365 23508 6377 23511
rect 6236 23480 6377 23508
rect 6236 23468 6242 23480
rect 6365 23477 6377 23480
rect 6411 23477 6423 23511
rect 6365 23471 6423 23477
rect 8205 23511 8263 23517
rect 8205 23477 8217 23511
rect 8251 23508 8263 23511
rect 8662 23508 8668 23520
rect 8251 23480 8668 23508
rect 8251 23477 8263 23480
rect 8205 23471 8263 23477
rect 8662 23468 8668 23480
rect 8720 23468 8726 23520
rect 9122 23468 9128 23520
rect 9180 23508 9186 23520
rect 9309 23511 9367 23517
rect 9309 23508 9321 23511
rect 9180 23480 9321 23508
rect 9180 23468 9186 23480
rect 9309 23477 9321 23480
rect 9355 23477 9367 23511
rect 9309 23471 9367 23477
rect 9674 23468 9680 23520
rect 9732 23468 9738 23520
rect 10410 23468 10416 23520
rect 10468 23468 10474 23520
rect 10594 23468 10600 23520
rect 10652 23468 10658 23520
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 13081 23511 13139 23517
rect 13081 23508 13093 23511
rect 12492 23480 13093 23508
rect 12492 23468 12498 23480
rect 13081 23477 13093 23480
rect 13127 23477 13139 23511
rect 13081 23471 13139 23477
rect 1104 23418 37076 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 37076 23418
rect 1104 23344 37076 23366
rect 4801 23307 4859 23313
rect 4801 23273 4813 23307
rect 4847 23304 4859 23307
rect 5074 23304 5080 23316
rect 4847 23276 5080 23304
rect 4847 23273 4859 23276
rect 4801 23267 4859 23273
rect 5074 23264 5080 23276
rect 5132 23264 5138 23316
rect 6362 23264 6368 23316
rect 6420 23304 6426 23316
rect 6733 23307 6791 23313
rect 6733 23304 6745 23307
rect 6420 23276 6745 23304
rect 6420 23264 6426 23276
rect 6733 23273 6745 23276
rect 6779 23273 6791 23307
rect 6733 23267 6791 23273
rect 8754 23264 8760 23316
rect 8812 23264 8818 23316
rect 9125 23307 9183 23313
rect 9125 23273 9137 23307
rect 9171 23304 9183 23307
rect 9214 23304 9220 23316
rect 9171 23276 9220 23304
rect 9171 23273 9183 23276
rect 9125 23267 9183 23273
rect 9214 23264 9220 23276
rect 9272 23264 9278 23316
rect 9309 23307 9367 23313
rect 9309 23273 9321 23307
rect 9355 23304 9367 23307
rect 9674 23304 9680 23316
rect 9355 23276 9680 23304
rect 9355 23273 9367 23276
rect 9309 23267 9367 23273
rect 9674 23264 9680 23276
rect 9732 23264 9738 23316
rect 10137 23307 10195 23313
rect 10137 23273 10149 23307
rect 10183 23304 10195 23307
rect 10410 23304 10416 23316
rect 10183 23276 10416 23304
rect 10183 23273 10195 23276
rect 10137 23267 10195 23273
rect 10410 23264 10416 23276
rect 10468 23264 10474 23316
rect 13906 23264 13912 23316
rect 13964 23304 13970 23316
rect 23474 23304 23480 23316
rect 13964 23276 14596 23304
rect 13964 23264 13970 23276
rect 9490 23196 9496 23248
rect 9548 23236 9554 23248
rect 9766 23236 9772 23248
rect 9548 23208 9772 23236
rect 9548 23196 9554 23208
rect 9766 23196 9772 23208
rect 9824 23196 9830 23248
rect 3142 23128 3148 23180
rect 3200 23168 3206 23180
rect 4985 23171 5043 23177
rect 4985 23168 4997 23171
rect 3200 23140 4997 23168
rect 3200 23128 3206 23140
rect 4985 23137 4997 23140
rect 5031 23137 5043 23171
rect 4985 23131 5043 23137
rect 5258 23128 5264 23180
rect 5316 23128 5322 23180
rect 7009 23171 7067 23177
rect 7009 23137 7021 23171
rect 7055 23168 7067 23171
rect 10318 23168 10324 23180
rect 7055 23140 10324 23168
rect 7055 23137 7067 23140
rect 7009 23131 7067 23137
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 12158 23128 12164 23180
rect 12216 23128 12222 23180
rect 12434 23128 12440 23180
rect 12492 23128 12498 23180
rect 14568 23177 14596 23276
rect 18524 23276 23480 23304
rect 14553 23171 14611 23177
rect 14553 23137 14565 23171
rect 14599 23137 14611 23171
rect 14553 23131 14611 23137
rect 14642 23128 14648 23180
rect 14700 23128 14706 23180
rect 2774 23060 2780 23112
rect 2832 23060 2838 23112
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23100 3019 23103
rect 3694 23100 3700 23112
rect 3007 23072 3700 23100
rect 3007 23069 3019 23072
rect 2961 23063 3019 23069
rect 3694 23060 3700 23072
rect 3752 23060 3758 23112
rect 3789 23103 3847 23109
rect 3789 23069 3801 23103
rect 3835 23069 3847 23103
rect 3789 23063 3847 23069
rect 3804 23032 3832 23063
rect 3970 23060 3976 23112
rect 4028 23060 4034 23112
rect 4062 23060 4068 23112
rect 4120 23100 4126 23112
rect 4709 23103 4767 23109
rect 4709 23100 4721 23103
rect 4120 23072 4721 23100
rect 4120 23060 4126 23072
rect 4709 23069 4721 23072
rect 4755 23100 4767 23103
rect 4755 23072 4936 23100
rect 4755 23069 4767 23072
rect 4709 23063 4767 23069
rect 4798 23032 4804 23044
rect 3804 23004 4804 23032
rect 4798 22992 4804 23004
rect 4856 22992 4862 23044
rect 4908 23032 4936 23072
rect 8294 23060 8300 23112
rect 8352 23100 8358 23112
rect 8352 23086 8418 23100
rect 8352 23072 8432 23086
rect 8352 23060 8358 23072
rect 5534 23032 5540 23044
rect 4908 23004 5540 23032
rect 5534 22992 5540 23004
rect 5592 22992 5598 23044
rect 6486 23004 6868 23032
rect 2682 22924 2688 22976
rect 2740 22964 2746 22976
rect 2777 22967 2835 22973
rect 2777 22964 2789 22967
rect 2740 22936 2789 22964
rect 2740 22924 2746 22936
rect 2777 22933 2789 22936
rect 2823 22933 2835 22967
rect 2777 22927 2835 22933
rect 3418 22924 3424 22976
rect 3476 22964 3482 22976
rect 3881 22967 3939 22973
rect 3881 22964 3893 22967
rect 3476 22936 3893 22964
rect 3476 22924 3482 22936
rect 3881 22933 3893 22936
rect 3927 22933 3939 22967
rect 3881 22927 3939 22933
rect 5258 22924 5264 22976
rect 5316 22964 5322 22976
rect 6564 22964 6592 23004
rect 5316 22936 6592 22964
rect 6840 22964 6868 23004
rect 7282 22992 7288 23044
rect 7340 22992 7346 23044
rect 8404 22964 8432 23072
rect 9122 23060 9128 23112
rect 9180 23100 9186 23112
rect 9180 23072 9628 23100
rect 9180 23060 9186 23072
rect 9490 22992 9496 23044
rect 9548 22992 9554 23044
rect 9600 23032 9628 23072
rect 9674 23060 9680 23112
rect 9732 23060 9738 23112
rect 9766 23060 9772 23112
rect 9824 23060 9830 23112
rect 9858 23060 9864 23112
rect 9916 23060 9922 23112
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 9968 23032 9996 23063
rect 15286 23060 15292 23112
rect 15344 23060 15350 23112
rect 18524 23109 18552 23276
rect 23474 23264 23480 23276
rect 23532 23264 23538 23316
rect 30650 23264 30656 23316
rect 30708 23304 30714 23316
rect 31665 23307 31723 23313
rect 31665 23304 31677 23307
rect 30708 23276 31677 23304
rect 30708 23264 30714 23276
rect 31665 23273 31677 23276
rect 31711 23273 31723 23307
rect 31665 23267 31723 23273
rect 34422 23264 34428 23316
rect 34480 23264 34486 23316
rect 20456 23208 22968 23236
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 18690 23060 18696 23112
rect 18748 23060 18754 23112
rect 20456 23109 20484 23208
rect 22940 23180 22968 23208
rect 27522 23196 27528 23248
rect 27580 23236 27586 23248
rect 27580 23208 28764 23236
rect 27580 23196 27586 23208
rect 20717 23171 20775 23177
rect 20717 23137 20729 23171
rect 20763 23168 20775 23171
rect 21358 23168 21364 23180
rect 20763 23140 21364 23168
rect 20763 23137 20775 23140
rect 20717 23131 20775 23137
rect 21358 23128 21364 23140
rect 21416 23168 21422 23180
rect 21416 23140 21864 23168
rect 21416 23128 21422 23140
rect 18785 23103 18843 23109
rect 18785 23069 18797 23103
rect 18831 23100 18843 23103
rect 20441 23103 20499 23109
rect 18831 23072 20116 23100
rect 18831 23069 18843 23072
rect 18785 23063 18843 23069
rect 9600 23004 9996 23032
rect 10042 22992 10048 23044
rect 10100 23032 10106 23044
rect 10597 23035 10655 23041
rect 10597 23032 10609 23035
rect 10100 23004 10609 23032
rect 10100 22992 10106 23004
rect 10597 23001 10609 23004
rect 10643 23001 10655 23035
rect 10597 22995 10655 23001
rect 11054 22992 11060 23044
rect 11112 22992 11118 23044
rect 13814 23032 13820 23044
rect 13662 23004 13820 23032
rect 13814 22992 13820 23004
rect 13872 23032 13878 23044
rect 13872 23004 14688 23032
rect 13872 22992 13878 23004
rect 6840 22936 8432 22964
rect 9293 22967 9351 22973
rect 5316 22924 5322 22936
rect 9293 22933 9305 22967
rect 9339 22964 9351 22967
rect 10870 22964 10876 22976
rect 9339 22936 10876 22964
rect 9339 22933 9351 22936
rect 9293 22927 9351 22933
rect 10870 22924 10876 22936
rect 10928 22964 10934 22976
rect 12069 22967 12127 22973
rect 12069 22964 12081 22967
rect 10928 22936 12081 22964
rect 10928 22924 10934 22936
rect 12069 22933 12081 22936
rect 12115 22933 12127 22967
rect 12069 22927 12127 22933
rect 13998 22924 14004 22976
rect 14056 22964 14062 22976
rect 14093 22967 14151 22973
rect 14093 22964 14105 22967
rect 14056 22936 14105 22964
rect 14056 22924 14062 22936
rect 14093 22933 14105 22936
rect 14139 22933 14151 22967
rect 14093 22927 14151 22933
rect 14461 22967 14519 22973
rect 14461 22933 14473 22967
rect 14507 22964 14519 22967
rect 14550 22964 14556 22976
rect 14507 22936 14556 22964
rect 14507 22933 14519 22936
rect 14461 22927 14519 22933
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 14660 22964 14688 23004
rect 15562 22992 15568 23044
rect 15620 22992 15626 23044
rect 16850 23032 16856 23044
rect 16790 23004 16856 23032
rect 16850 22992 16856 23004
rect 16908 23032 16914 23044
rect 16908 23004 17172 23032
rect 16908 22992 16914 23004
rect 15838 22964 15844 22976
rect 14660 22936 15844 22964
rect 15838 22924 15844 22936
rect 15896 22924 15902 22976
rect 17034 22924 17040 22976
rect 17092 22924 17098 22976
rect 17144 22964 17172 23004
rect 18046 22992 18052 23044
rect 18104 22992 18110 23044
rect 19978 22992 19984 23044
rect 20036 22992 20042 23044
rect 20088 23032 20116 23072
rect 20441 23069 20453 23103
rect 20487 23069 20499 23103
rect 20441 23063 20499 23069
rect 20530 23060 20536 23112
rect 20588 23100 20594 23112
rect 21836 23109 21864 23140
rect 22922 23128 22928 23180
rect 22980 23128 22986 23180
rect 23658 23128 23664 23180
rect 23716 23168 23722 23180
rect 25225 23171 25283 23177
rect 25225 23168 25237 23171
rect 23716 23140 25237 23168
rect 23716 23128 23722 23140
rect 25225 23137 25237 23140
rect 25271 23168 25283 23171
rect 26234 23168 26240 23180
rect 25271 23140 26240 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 26234 23128 26240 23140
rect 26292 23168 26298 23180
rect 26970 23168 26976 23180
rect 26292 23140 26976 23168
rect 26292 23128 26298 23140
rect 26970 23128 26976 23140
rect 27028 23128 27034 23180
rect 28736 23177 28764 23208
rect 28721 23171 28779 23177
rect 28721 23137 28733 23171
rect 28767 23137 28779 23171
rect 28721 23131 28779 23137
rect 30190 23128 30196 23180
rect 30248 23128 30254 23180
rect 32122 23128 32128 23180
rect 32180 23168 32186 23180
rect 32677 23171 32735 23177
rect 32677 23168 32689 23171
rect 32180 23140 32689 23168
rect 32180 23128 32186 23140
rect 32677 23137 32689 23140
rect 32723 23137 32735 23171
rect 32677 23131 32735 23137
rect 20625 23103 20683 23109
rect 20625 23100 20637 23103
rect 20588 23072 20637 23100
rect 20588 23060 20594 23072
rect 20625 23069 20637 23072
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 21637 23103 21695 23109
rect 21637 23069 21649 23103
rect 21683 23069 21695 23103
rect 21637 23063 21695 23069
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 21913 23103 21971 23109
rect 21913 23069 21925 23103
rect 21959 23100 21971 23103
rect 22462 23100 22468 23112
rect 21959 23072 22468 23100
rect 21959 23069 21971 23072
rect 21913 23063 21971 23069
rect 20548 23032 20576 23060
rect 20088 23004 20576 23032
rect 21174 22992 21180 23044
rect 21232 22992 21238 23044
rect 21652 23032 21680 23063
rect 22462 23060 22468 23072
rect 22520 23100 22526 23112
rect 22833 23103 22891 23109
rect 22833 23100 22845 23103
rect 22520 23072 22845 23100
rect 22520 23060 22526 23072
rect 22833 23069 22845 23072
rect 22879 23069 22891 23103
rect 22833 23063 22891 23069
rect 27525 23103 27583 23109
rect 27525 23069 27537 23103
rect 27571 23100 27583 23103
rect 27614 23100 27620 23112
rect 27571 23072 27620 23100
rect 27571 23069 27583 23072
rect 27525 23063 27583 23069
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 27709 23103 27767 23109
rect 27709 23069 27721 23103
rect 27755 23069 27767 23103
rect 27709 23063 27767 23069
rect 27801 23103 27859 23109
rect 27801 23069 27813 23103
rect 27847 23100 27859 23103
rect 28626 23100 28632 23112
rect 27847 23072 28632 23100
rect 27847 23069 27859 23072
rect 27801 23063 27859 23069
rect 22741 23035 22799 23041
rect 21652 23004 22692 23032
rect 18138 22964 18144 22976
rect 17144 22936 18144 22964
rect 18138 22924 18144 22936
rect 18196 22924 18202 22976
rect 22186 22924 22192 22976
rect 22244 22964 22250 22976
rect 22373 22967 22431 22973
rect 22373 22964 22385 22967
rect 22244 22936 22385 22964
rect 22244 22924 22250 22936
rect 22373 22933 22385 22936
rect 22419 22933 22431 22967
rect 22664 22964 22692 23004
rect 22741 23001 22753 23035
rect 22787 23032 22799 23035
rect 23566 23032 23572 23044
rect 22787 23004 23572 23032
rect 22787 23001 22799 23004
rect 22741 22995 22799 23001
rect 23566 22992 23572 23004
rect 23624 22992 23630 23044
rect 25501 23035 25559 23041
rect 25501 23001 25513 23035
rect 25547 23001 25559 23035
rect 25501 22995 25559 23001
rect 23934 22964 23940 22976
rect 22664 22936 23940 22964
rect 22373 22927 22431 22933
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 25516 22964 25544 22995
rect 26142 22992 26148 23044
rect 26200 22992 26206 23044
rect 27065 23035 27123 23041
rect 27065 23001 27077 23035
rect 27111 23032 27123 23035
rect 27246 23032 27252 23044
rect 27111 23004 27252 23032
rect 27111 23001 27123 23004
rect 27065 22995 27123 23001
rect 27246 22992 27252 23004
rect 27304 22992 27310 23044
rect 26234 22964 26240 22976
rect 25516 22936 26240 22964
rect 26234 22924 26240 22936
rect 26292 22924 26298 22976
rect 26878 22924 26884 22976
rect 26936 22964 26942 22976
rect 26973 22967 27031 22973
rect 26973 22964 26985 22967
rect 26936 22936 26985 22964
rect 26936 22924 26942 22936
rect 26973 22933 26985 22936
rect 27019 22964 27031 22967
rect 27724 22964 27752 23063
rect 28626 23060 28632 23072
rect 28684 23060 28690 23112
rect 28994 23060 29000 23112
rect 29052 23100 29058 23112
rect 29546 23100 29552 23112
rect 29052 23072 29552 23100
rect 29052 23060 29058 23072
rect 29546 23060 29552 23072
rect 29604 23100 29610 23112
rect 29917 23103 29975 23109
rect 29917 23100 29929 23103
rect 29604 23072 29929 23100
rect 29604 23060 29610 23072
rect 29917 23069 29929 23072
rect 29963 23069 29975 23103
rect 29917 23063 29975 23069
rect 32953 23035 33011 23041
rect 31418 23004 31524 23032
rect 31496 22976 31524 23004
rect 32953 23001 32965 23035
rect 32999 23032 33011 23035
rect 33226 23032 33232 23044
rect 32999 23004 33232 23032
rect 32999 23001 33011 23004
rect 32953 22995 33011 23001
rect 33226 22992 33232 23004
rect 33284 22992 33290 23044
rect 33410 23032 33416 23044
rect 33336 23004 33416 23032
rect 27019 22936 27752 22964
rect 27019 22933 27031 22936
rect 26973 22927 27031 22933
rect 27890 22924 27896 22976
rect 27948 22964 27954 22976
rect 28169 22967 28227 22973
rect 28169 22964 28181 22967
rect 27948 22936 28181 22964
rect 27948 22924 27954 22936
rect 28169 22933 28181 22936
rect 28215 22933 28227 22967
rect 28169 22927 28227 22933
rect 28537 22967 28595 22973
rect 28537 22933 28549 22967
rect 28583 22964 28595 22967
rect 29362 22964 29368 22976
rect 28583 22936 29368 22964
rect 28583 22933 28595 22936
rect 28537 22927 28595 22933
rect 29362 22924 29368 22936
rect 29420 22924 29426 22976
rect 31478 22924 31484 22976
rect 31536 22964 31542 22976
rect 33336 22964 33364 23004
rect 33410 22992 33416 23004
rect 33468 22992 33474 23044
rect 31536 22936 33364 22964
rect 31536 22924 31542 22936
rect 1104 22874 37076 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 37076 22874
rect 1104 22800 37076 22822
rect 1118 22720 1124 22772
rect 1176 22760 1182 22772
rect 1176 22732 6408 22760
rect 1176 22720 1182 22732
rect 2682 22652 2688 22704
rect 2740 22652 2746 22704
rect 3418 22652 3424 22704
rect 3476 22652 3482 22704
rect 3694 22652 3700 22704
rect 3752 22692 3758 22704
rect 3752 22664 3910 22692
rect 3752 22652 3758 22664
rect 4798 22652 4804 22704
rect 4856 22692 4862 22704
rect 5169 22695 5227 22701
rect 5169 22692 5181 22695
rect 4856 22664 5181 22692
rect 4856 22652 4862 22664
rect 5169 22661 5181 22664
rect 5215 22661 5227 22695
rect 5169 22655 5227 22661
rect 5534 22652 5540 22704
rect 5592 22652 5598 22704
rect 5626 22652 5632 22704
rect 5684 22692 5690 22704
rect 5813 22695 5871 22701
rect 5813 22692 5825 22695
rect 5684 22664 5825 22692
rect 5684 22652 5690 22664
rect 5813 22661 5825 22664
rect 5859 22661 5871 22695
rect 5813 22655 5871 22661
rect 6029 22695 6087 22701
rect 6029 22661 6041 22695
rect 6075 22692 6087 22695
rect 6270 22692 6276 22704
rect 6075 22664 6276 22692
rect 6075 22661 6087 22664
rect 6029 22655 6087 22661
rect 6270 22652 6276 22664
rect 6328 22652 6334 22704
rect 6380 22701 6408 22732
rect 7282 22720 7288 22772
rect 7340 22760 7346 22772
rect 8205 22763 8263 22769
rect 8205 22760 8217 22763
rect 7340 22732 8217 22760
rect 7340 22720 7346 22732
rect 8205 22729 8217 22732
rect 8251 22729 8263 22763
rect 8205 22723 8263 22729
rect 8570 22720 8576 22772
rect 8628 22720 8634 22772
rect 8662 22720 8668 22772
rect 8720 22720 8726 22772
rect 9401 22763 9459 22769
rect 9401 22729 9413 22763
rect 9447 22760 9459 22763
rect 9447 22732 9720 22760
rect 9447 22729 9459 22732
rect 9401 22723 9459 22729
rect 6365 22695 6423 22701
rect 6365 22661 6377 22695
rect 6411 22661 6423 22695
rect 6365 22655 6423 22661
rect 9033 22695 9091 22701
rect 9033 22661 9045 22695
rect 9079 22661 9091 22695
rect 9033 22655 9091 22661
rect 2041 22627 2099 22633
rect 2041 22593 2053 22627
rect 2087 22624 2099 22627
rect 2087 22596 2360 22624
rect 2087 22593 2099 22596
rect 2041 22587 2099 22593
rect 2332 22497 2360 22596
rect 3142 22584 3148 22636
rect 3200 22584 3206 22636
rect 5353 22627 5411 22633
rect 5353 22593 5365 22627
rect 5399 22593 5411 22627
rect 5353 22587 5411 22593
rect 5445 22627 5503 22633
rect 5445 22593 5457 22627
rect 5491 22624 5503 22627
rect 6914 22624 6920 22636
rect 5491 22596 6920 22624
rect 5491 22593 5503 22596
rect 5445 22587 5503 22593
rect 2774 22516 2780 22568
rect 2832 22516 2838 22568
rect 2961 22559 3019 22565
rect 2961 22525 2973 22559
rect 3007 22556 3019 22559
rect 4062 22556 4068 22568
rect 3007 22528 4068 22556
rect 3007 22525 3019 22528
rect 2961 22519 3019 22525
rect 4062 22516 4068 22528
rect 4120 22516 4126 22568
rect 4798 22516 4804 22568
rect 4856 22556 4862 22568
rect 5258 22556 5264 22568
rect 4856 22528 5264 22556
rect 4856 22516 4862 22528
rect 5258 22516 5264 22528
rect 5316 22516 5322 22568
rect 5368 22556 5396 22587
rect 6914 22584 6920 22596
rect 6972 22624 6978 22636
rect 9048 22624 9076 22655
rect 9122 22652 9128 22704
rect 9180 22692 9186 22704
rect 9233 22695 9291 22701
rect 9233 22692 9245 22695
rect 9180 22664 9245 22692
rect 9180 22652 9186 22664
rect 9233 22661 9245 22664
rect 9279 22661 9291 22695
rect 9233 22655 9291 22661
rect 9692 22692 9720 22732
rect 10042 22720 10048 22772
rect 10100 22720 10106 22772
rect 10137 22763 10195 22769
rect 10137 22729 10149 22763
rect 10183 22760 10195 22763
rect 10502 22760 10508 22772
rect 10183 22732 10508 22760
rect 10183 22729 10195 22732
rect 10137 22723 10195 22729
rect 10502 22720 10508 22732
rect 10560 22720 10566 22772
rect 14090 22760 14096 22772
rect 12268 22732 14096 22760
rect 10778 22692 10784 22704
rect 9692 22664 10364 22692
rect 6972 22596 9076 22624
rect 6972 22584 6978 22596
rect 9398 22584 9404 22636
rect 9456 22624 9462 22636
rect 9692 22633 9720 22664
rect 10336 22633 10364 22664
rect 10612 22664 10784 22692
rect 9493 22627 9551 22633
rect 9493 22624 9505 22627
rect 9456 22596 9505 22624
rect 9456 22584 9462 22596
rect 9493 22593 9505 22596
rect 9539 22593 9551 22627
rect 9493 22587 9551 22593
rect 9677 22627 9735 22633
rect 9677 22593 9689 22627
rect 9723 22593 9735 22627
rect 9677 22587 9735 22593
rect 10229 22627 10287 22633
rect 10229 22593 10241 22627
rect 10275 22593 10287 22627
rect 10229 22587 10287 22593
rect 10321 22627 10379 22633
rect 10321 22593 10333 22627
rect 10367 22624 10379 22627
rect 10410 22624 10416 22636
rect 10367 22596 10416 22624
rect 10367 22593 10379 22596
rect 10321 22587 10379 22593
rect 6546 22556 6552 22568
rect 5368 22528 6552 22556
rect 2317 22491 2375 22497
rect 2317 22457 2329 22491
rect 2363 22457 2375 22491
rect 2317 22451 2375 22457
rect 5718 22448 5724 22500
rect 5776 22448 5782 22500
rect 1670 22380 1676 22432
rect 1728 22420 1734 22432
rect 1949 22423 2007 22429
rect 1949 22420 1961 22423
rect 1728 22392 1961 22420
rect 1728 22380 1734 22392
rect 1949 22389 1961 22392
rect 1995 22389 2007 22423
rect 1949 22383 2007 22389
rect 4890 22380 4896 22432
rect 4948 22420 4954 22432
rect 5442 22420 5448 22432
rect 4948 22392 5448 22420
rect 4948 22380 4954 22392
rect 5442 22380 5448 22392
rect 5500 22380 5506 22432
rect 6012 22429 6040 22528
rect 6546 22516 6552 22528
rect 6604 22516 6610 22568
rect 8849 22559 8907 22565
rect 8849 22525 8861 22559
rect 8895 22556 8907 22559
rect 9585 22559 9643 22565
rect 9585 22556 9597 22559
rect 8895 22528 9597 22556
rect 8895 22525 8907 22528
rect 8849 22519 8907 22525
rect 9585 22525 9597 22528
rect 9631 22556 9643 22559
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 9631 22528 9781 22556
rect 9631 22525 9643 22528
rect 9585 22519 9643 22525
rect 9769 22525 9781 22528
rect 9815 22525 9827 22559
rect 10244 22556 10272 22587
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 10502 22584 10508 22636
rect 10560 22584 10566 22636
rect 10612 22633 10640 22664
rect 10778 22652 10784 22664
rect 10836 22652 10842 22704
rect 10597 22627 10655 22633
rect 10597 22593 10609 22627
rect 10643 22593 10655 22627
rect 10597 22587 10655 22593
rect 10686 22584 10692 22636
rect 10744 22584 10750 22636
rect 10870 22584 10876 22636
rect 10928 22584 10934 22636
rect 12158 22584 12164 22636
rect 12216 22624 12222 22636
rect 12268 22633 12296 22732
rect 14090 22720 14096 22732
rect 14148 22760 14154 22772
rect 14458 22760 14464 22772
rect 14148 22732 14464 22760
rect 14148 22720 14154 22732
rect 14458 22720 14464 22732
rect 14516 22760 14522 22772
rect 15286 22760 15292 22772
rect 14516 22732 15292 22760
rect 14516 22720 14522 22732
rect 15286 22720 15292 22732
rect 15344 22720 15350 22772
rect 17221 22763 17279 22769
rect 17221 22729 17233 22763
rect 17267 22760 17279 22763
rect 17310 22760 17316 22772
rect 17267 22732 17316 22760
rect 17267 22729 17279 22732
rect 17221 22723 17279 22729
rect 17310 22720 17316 22732
rect 17368 22720 17374 22772
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 20622 22760 20628 22772
rect 19668 22732 20628 22760
rect 19668 22720 19674 22732
rect 20622 22720 20628 22732
rect 20680 22760 20686 22772
rect 20680 22732 21956 22760
rect 20680 22720 20686 22732
rect 13814 22692 13820 22704
rect 13754 22664 13820 22692
rect 13814 22652 13820 22664
rect 13872 22652 13878 22704
rect 15838 22692 15844 22704
rect 15594 22664 15844 22692
rect 15838 22652 15844 22664
rect 15896 22692 15902 22704
rect 16850 22692 16856 22704
rect 15896 22664 16856 22692
rect 15896 22652 15902 22664
rect 16850 22652 16856 22664
rect 16908 22652 16914 22704
rect 18046 22652 18052 22704
rect 18104 22652 18110 22704
rect 18138 22652 18144 22704
rect 18196 22692 18202 22704
rect 19889 22695 19947 22701
rect 18196 22664 18538 22692
rect 18196 22652 18202 22664
rect 19889 22661 19901 22695
rect 19935 22692 19947 22695
rect 19978 22692 19984 22704
rect 19935 22664 19984 22692
rect 19935 22661 19947 22664
rect 19889 22655 19947 22661
rect 19978 22652 19984 22664
rect 20036 22652 20042 22704
rect 12253 22627 12311 22633
rect 12253 22624 12265 22627
rect 12216 22596 12265 22624
rect 12216 22584 12222 22596
rect 12253 22593 12265 22596
rect 12299 22593 12311 22627
rect 12253 22587 12311 22593
rect 14090 22584 14096 22636
rect 14148 22584 14154 22636
rect 17034 22584 17040 22636
rect 17092 22624 17098 22636
rect 17313 22627 17371 22633
rect 17313 22624 17325 22627
rect 17092 22596 17325 22624
rect 17092 22584 17098 22596
rect 17313 22593 17325 22596
rect 17359 22593 17371 22627
rect 19610 22624 19616 22636
rect 17313 22587 17371 22593
rect 19444 22596 19616 22624
rect 10781 22559 10839 22565
rect 10781 22556 10793 22559
rect 10244 22528 10793 22556
rect 9769 22519 9827 22525
rect 10781 22525 10793 22528
rect 10827 22525 10839 22559
rect 10781 22519 10839 22525
rect 12529 22559 12587 22565
rect 12529 22525 12541 22559
rect 12575 22556 12587 22559
rect 13998 22556 14004 22568
rect 12575 22528 14004 22556
rect 12575 22525 12587 22528
rect 12529 22519 12587 22525
rect 13998 22516 14004 22528
rect 14056 22516 14062 22568
rect 14366 22516 14372 22568
rect 14424 22516 14430 22568
rect 17126 22516 17132 22568
rect 17184 22556 17190 22568
rect 17405 22559 17463 22565
rect 17405 22556 17417 22559
rect 17184 22528 17417 22556
rect 17184 22516 17190 22528
rect 17405 22525 17417 22528
rect 17451 22525 17463 22559
rect 17405 22519 17463 22525
rect 17773 22559 17831 22565
rect 17773 22525 17785 22559
rect 17819 22556 17831 22559
rect 19444 22556 19472 22596
rect 19610 22584 19616 22596
rect 19668 22584 19674 22636
rect 21928 22633 21956 22732
rect 23566 22720 23572 22772
rect 23624 22760 23630 22772
rect 23661 22763 23719 22769
rect 23661 22760 23673 22763
rect 23624 22732 23673 22760
rect 23624 22720 23630 22732
rect 23661 22729 23673 22732
rect 23707 22729 23719 22763
rect 23661 22723 23719 22729
rect 23934 22720 23940 22772
rect 23992 22760 23998 22772
rect 27062 22760 27068 22772
rect 23992 22732 27068 22760
rect 23992 22720 23998 22732
rect 27062 22720 27068 22732
rect 27120 22720 27126 22772
rect 27172 22732 27384 22760
rect 22186 22652 22192 22704
rect 22244 22652 22250 22704
rect 22646 22652 22652 22704
rect 22704 22652 22710 22704
rect 26142 22692 26148 22704
rect 25424 22664 26148 22692
rect 25424 22636 25452 22664
rect 26142 22652 26148 22664
rect 26200 22692 26206 22704
rect 27172 22692 27200 22732
rect 26200 22664 27200 22692
rect 26200 22652 26206 22664
rect 27246 22652 27252 22704
rect 27304 22652 27310 22704
rect 27356 22692 27384 22732
rect 28626 22720 28632 22772
rect 28684 22760 28690 22772
rect 28721 22763 28779 22769
rect 28721 22760 28733 22763
rect 28684 22732 28733 22760
rect 28684 22720 28690 22732
rect 28721 22729 28733 22732
rect 28767 22729 28779 22763
rect 28721 22723 28779 22729
rect 30742 22720 30748 22772
rect 30800 22720 30806 22772
rect 33870 22720 33876 22772
rect 33928 22720 33934 22772
rect 31478 22692 31484 22704
rect 27356 22664 27738 22692
rect 30498 22664 31484 22692
rect 31478 22652 31484 22664
rect 31536 22652 31542 22704
rect 32398 22652 32404 22704
rect 32456 22652 32462 22704
rect 33410 22652 33416 22704
rect 33468 22652 33474 22704
rect 21913 22627 21971 22633
rect 17819 22528 19472 22556
rect 19521 22559 19579 22565
rect 17819 22525 17831 22528
rect 17773 22519 17831 22525
rect 19521 22525 19533 22559
rect 19567 22556 19579 22559
rect 20530 22556 20536 22568
rect 19567 22528 20536 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 21008 22556 21036 22610
rect 21913 22593 21925 22627
rect 21959 22593 21971 22627
rect 21913 22587 21971 22593
rect 23658 22584 23664 22636
rect 23716 22624 23722 22636
rect 23753 22627 23811 22633
rect 23753 22624 23765 22627
rect 23716 22596 23765 22624
rect 23716 22584 23722 22596
rect 23753 22593 23765 22596
rect 23799 22593 23811 22627
rect 25406 22624 25412 22636
rect 25162 22596 25412 22624
rect 23753 22587 23811 22593
rect 25406 22584 25412 22596
rect 25464 22584 25470 22636
rect 25958 22584 25964 22636
rect 26016 22584 26022 22636
rect 28994 22584 29000 22636
rect 29052 22584 29058 22636
rect 32122 22584 32128 22636
rect 32180 22584 32186 22636
rect 22554 22556 22560 22568
rect 21008 22528 22560 22556
rect 22554 22516 22560 22528
rect 22612 22516 22618 22568
rect 24026 22516 24032 22568
rect 24084 22516 24090 22568
rect 26053 22559 26111 22565
rect 26053 22525 26065 22559
rect 26099 22525 26111 22559
rect 26053 22519 26111 22525
rect 21358 22448 21364 22500
rect 21416 22448 21422 22500
rect 25038 22448 25044 22500
rect 25096 22488 25102 22500
rect 25593 22491 25651 22497
rect 25593 22488 25605 22491
rect 25096 22460 25605 22488
rect 25096 22448 25102 22460
rect 25593 22457 25605 22460
rect 25639 22457 25651 22491
rect 25593 22451 25651 22457
rect 5997 22423 6055 22429
rect 5997 22389 6009 22423
rect 6043 22389 6055 22423
rect 5997 22383 6055 22389
rect 6181 22423 6239 22429
rect 6181 22389 6193 22423
rect 6227 22420 6239 22423
rect 7282 22420 7288 22432
rect 6227 22392 7288 22420
rect 6227 22389 6239 22392
rect 6181 22383 6239 22389
rect 7282 22380 7288 22392
rect 7340 22380 7346 22432
rect 7650 22380 7656 22432
rect 7708 22380 7714 22432
rect 8202 22380 8208 22432
rect 8260 22420 8266 22432
rect 8386 22420 8392 22432
rect 8260 22392 8392 22420
rect 8260 22380 8266 22392
rect 8386 22380 8392 22392
rect 8444 22420 8450 22432
rect 9217 22423 9275 22429
rect 9217 22420 9229 22423
rect 8444 22392 9229 22420
rect 8444 22380 8450 22392
rect 9217 22389 9229 22392
rect 9263 22389 9275 22423
rect 9217 22383 9275 22389
rect 9766 22380 9772 22432
rect 9824 22420 9830 22432
rect 10778 22420 10784 22432
rect 9824 22392 10784 22420
rect 9824 22380 9830 22392
rect 10778 22380 10784 22392
rect 10836 22380 10842 22432
rect 14001 22423 14059 22429
rect 14001 22389 14013 22423
rect 14047 22420 14059 22423
rect 14550 22420 14556 22432
rect 14047 22392 14556 22420
rect 14047 22389 14059 22392
rect 14001 22383 14059 22389
rect 14550 22380 14556 22392
rect 14608 22420 14614 22432
rect 15010 22420 15016 22432
rect 14608 22392 15016 22420
rect 14608 22380 14614 22392
rect 15010 22380 15016 22392
rect 15068 22380 15074 22432
rect 15838 22380 15844 22432
rect 15896 22380 15902 22432
rect 16850 22380 16856 22432
rect 16908 22380 16914 22432
rect 25498 22380 25504 22432
rect 25556 22420 25562 22432
rect 26068 22420 26096 22519
rect 26142 22516 26148 22568
rect 26200 22556 26206 22568
rect 26418 22556 26424 22568
rect 26200 22528 26424 22556
rect 26200 22516 26206 22528
rect 26418 22516 26424 22528
rect 26476 22516 26482 22568
rect 26970 22516 26976 22568
rect 27028 22516 27034 22568
rect 29270 22516 29276 22568
rect 29328 22516 29334 22568
rect 25556 22392 26096 22420
rect 25556 22380 25562 22392
rect 27062 22380 27068 22432
rect 27120 22420 27126 22432
rect 30006 22420 30012 22432
rect 27120 22392 30012 22420
rect 27120 22380 27126 22392
rect 30006 22380 30012 22392
rect 30064 22420 30070 22432
rect 30466 22420 30472 22432
rect 30064 22392 30472 22420
rect 30064 22380 30070 22392
rect 30466 22380 30472 22392
rect 30524 22380 30530 22432
rect 1104 22330 37076 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 37076 22330
rect 1104 22256 37076 22278
rect 1670 22225 1676 22228
rect 1660 22219 1676 22225
rect 1660 22185 1672 22219
rect 1660 22179 1676 22185
rect 1670 22176 1676 22179
rect 1728 22176 1734 22228
rect 3789 22219 3847 22225
rect 3789 22185 3801 22219
rect 3835 22216 3847 22219
rect 3970 22216 3976 22228
rect 3835 22188 3976 22216
rect 3835 22185 3847 22188
rect 3789 22179 3847 22185
rect 3970 22176 3976 22188
rect 4028 22176 4034 22228
rect 5442 22176 5448 22228
rect 5500 22216 5506 22228
rect 5629 22219 5687 22225
rect 5629 22216 5641 22219
rect 5500 22188 5641 22216
rect 5500 22176 5506 22188
rect 5629 22185 5641 22188
rect 5675 22185 5687 22219
rect 5629 22179 5687 22185
rect 2774 22108 2780 22160
rect 2832 22148 2838 22160
rect 3145 22151 3203 22157
rect 3145 22148 3157 22151
rect 2832 22120 3157 22148
rect 2832 22108 2838 22120
rect 3145 22117 3157 22120
rect 3191 22148 3203 22151
rect 5644 22148 5672 22179
rect 6270 22176 6276 22228
rect 6328 22216 6334 22228
rect 6549 22219 6607 22225
rect 6549 22216 6561 22219
rect 6328 22188 6561 22216
rect 6328 22176 6334 22188
rect 6549 22185 6561 22188
rect 6595 22185 6607 22219
rect 6549 22179 6607 22185
rect 6733 22219 6791 22225
rect 6733 22185 6745 22219
rect 6779 22185 6791 22219
rect 6733 22179 6791 22185
rect 6748 22148 6776 22179
rect 10594 22176 10600 22228
rect 10652 22216 10658 22228
rect 10762 22219 10820 22225
rect 10762 22216 10774 22219
rect 10652 22188 10774 22216
rect 10652 22176 10658 22188
rect 10762 22185 10774 22188
rect 10808 22185 10820 22219
rect 10762 22179 10820 22185
rect 14366 22176 14372 22228
rect 14424 22216 14430 22228
rect 14553 22219 14611 22225
rect 14553 22216 14565 22219
rect 14424 22188 14565 22216
rect 14424 22176 14430 22188
rect 14553 22185 14565 22188
rect 14599 22185 14611 22219
rect 14553 22179 14611 22185
rect 15562 22176 15568 22228
rect 15620 22176 15626 22228
rect 16656 22219 16714 22225
rect 16656 22185 16668 22219
rect 16702 22216 16714 22219
rect 16850 22216 16856 22228
rect 16702 22188 16856 22216
rect 16702 22185 16714 22188
rect 16656 22179 16714 22185
rect 16850 22176 16856 22188
rect 16908 22176 16914 22228
rect 20980 22219 21038 22225
rect 20980 22185 20992 22219
rect 21026 22216 21038 22219
rect 21174 22216 21180 22228
rect 21026 22188 21180 22216
rect 21026 22185 21038 22188
rect 20980 22179 21038 22185
rect 21174 22176 21180 22188
rect 21232 22176 21238 22228
rect 22462 22176 22468 22228
rect 22520 22176 22526 22228
rect 24660 22219 24718 22225
rect 24660 22185 24672 22219
rect 24706 22216 24718 22219
rect 25038 22216 25044 22228
rect 24706 22188 25044 22216
rect 24706 22185 24718 22188
rect 24660 22179 24718 22185
rect 25038 22176 25044 22188
rect 25096 22176 25102 22228
rect 25958 22176 25964 22228
rect 26016 22216 26022 22228
rect 26145 22219 26203 22225
rect 26145 22216 26157 22219
rect 26016 22188 26157 22216
rect 26016 22176 26022 22188
rect 26145 22185 26157 22188
rect 26191 22185 26203 22219
rect 26145 22179 26203 22185
rect 3191 22120 5028 22148
rect 5644 22120 6776 22148
rect 3191 22117 3203 22120
rect 3145 22111 3203 22117
rect 1394 21972 1400 22024
rect 1452 21972 1458 22024
rect 3804 22021 3832 22120
rect 4890 22080 4896 22092
rect 4080 22052 4896 22080
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 21981 3847 22015
rect 3789 21975 3847 21981
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 4080 22021 4108 22052
rect 4890 22040 4896 22052
rect 4948 22040 4954 22092
rect 5000 22080 5028 22120
rect 9674 22108 9680 22160
rect 9732 22148 9738 22160
rect 10502 22148 10508 22160
rect 9732 22120 10508 22148
rect 9732 22108 9738 22120
rect 10502 22108 10508 22120
rect 10560 22108 10566 22160
rect 15378 22148 15384 22160
rect 15120 22120 15384 22148
rect 5810 22080 5816 22092
rect 5000 22052 5816 22080
rect 5644 22021 5672 22052
rect 5810 22040 5816 22052
rect 5868 22080 5874 22092
rect 6822 22080 6828 22092
rect 5868 22052 6828 22080
rect 5868 22040 5874 22052
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 7098 22040 7104 22092
rect 7156 22080 7162 22092
rect 7469 22083 7527 22089
rect 7469 22080 7481 22083
rect 7156 22052 7481 22080
rect 7156 22040 7162 22052
rect 7469 22049 7481 22052
rect 7515 22049 7527 22083
rect 10520 22080 10548 22108
rect 12253 22083 12311 22089
rect 12253 22080 12265 22083
rect 10520 22052 12265 22080
rect 7469 22043 7527 22049
rect 12253 22049 12265 22052
rect 12299 22049 12311 22083
rect 12253 22043 12311 22049
rect 15010 22040 15016 22092
rect 15068 22040 15074 22092
rect 15120 22089 15148 22120
rect 15378 22108 15384 22120
rect 15436 22148 15442 22160
rect 15436 22120 16160 22148
rect 15436 22108 15442 22120
rect 15105 22083 15163 22089
rect 15105 22049 15117 22083
rect 15151 22049 15163 22083
rect 15838 22080 15844 22092
rect 15105 22043 15163 22049
rect 15212 22052 15844 22080
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 4162 22015 4220 22021
rect 4162 21981 4174 22015
rect 4208 22012 4220 22015
rect 4617 22015 4675 22021
rect 4617 22012 4629 22015
rect 4208 21984 4629 22012
rect 4208 21981 4220 21984
rect 4162 21975 4220 21981
rect 4617 21981 4629 21984
rect 4663 21981 4675 22015
rect 5537 22015 5595 22021
rect 5537 22012 5549 22015
rect 4617 21975 4675 21981
rect 4724 21984 5549 22012
rect 2958 21944 2964 21956
rect 2898 21916 2964 21944
rect 2958 21904 2964 21916
rect 3016 21904 3022 21956
rect 3878 21904 3884 21956
rect 3936 21944 3942 21956
rect 4172 21944 4200 21975
rect 3936 21916 4200 21944
rect 3936 21904 3942 21916
rect 4338 21904 4344 21956
rect 4396 21904 4402 21956
rect 4724 21888 4752 21984
rect 5537 21981 5549 21984
rect 5583 21981 5595 22015
rect 5537 21975 5595 21981
rect 5629 22015 5687 22021
rect 5629 21981 5641 22015
rect 5675 21981 5687 22015
rect 5629 21975 5687 21981
rect 5905 22015 5963 22021
rect 5905 21981 5917 22015
rect 5951 22012 5963 22015
rect 5951 21984 7144 22012
rect 5951 21981 5963 21984
rect 5905 21975 5963 21981
rect 5353 21947 5411 21953
rect 5353 21913 5365 21947
rect 5399 21913 5411 21947
rect 5552 21944 5580 21975
rect 6701 21947 6759 21953
rect 6701 21944 6713 21947
rect 5552 21916 6713 21944
rect 5353 21907 5411 21913
rect 6701 21913 6713 21916
rect 6747 21913 6759 21947
rect 6701 21907 6759 21913
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4439 21879 4497 21885
rect 4439 21876 4451 21879
rect 4212 21848 4451 21876
rect 4212 21836 4218 21848
rect 4439 21845 4451 21848
rect 4485 21845 4497 21879
rect 4439 21839 4497 21845
rect 4525 21879 4583 21885
rect 4525 21845 4537 21879
rect 4571 21876 4583 21879
rect 4706 21876 4712 21888
rect 4571 21848 4712 21876
rect 4571 21845 4583 21848
rect 4525 21839 4583 21845
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 5368 21876 5396 21907
rect 6822 21904 6828 21956
rect 6880 21944 6886 21956
rect 6917 21947 6975 21953
rect 6917 21944 6929 21947
rect 6880 21916 6929 21944
rect 6880 21904 6886 21916
rect 6917 21913 6929 21916
rect 6963 21913 6975 21947
rect 6917 21907 6975 21913
rect 7116 21888 7144 21984
rect 7282 21972 7288 22024
rect 7340 22012 7346 22024
rect 8202 22012 8208 22024
rect 7340 21984 8208 22012
rect 7340 21972 7346 21984
rect 8202 21972 8208 21984
rect 8260 21972 8266 22024
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10505 22015 10563 22021
rect 10505 22012 10517 22015
rect 10100 21984 10517 22012
rect 10100 21972 10106 21984
rect 10505 21981 10517 21984
rect 10551 21981 10563 22015
rect 10505 21975 10563 21981
rect 14921 22015 14979 22021
rect 14921 21981 14933 22015
rect 14967 22012 14979 22015
rect 15212 22012 15240 22052
rect 15838 22040 15844 22052
rect 15896 22080 15902 22092
rect 16132 22089 16160 22120
rect 16025 22083 16083 22089
rect 16025 22080 16037 22083
rect 15896 22052 16037 22080
rect 15896 22040 15902 22052
rect 16025 22049 16037 22052
rect 16071 22049 16083 22083
rect 16025 22043 16083 22049
rect 16117 22083 16175 22089
rect 16117 22049 16129 22083
rect 16163 22049 16175 22083
rect 16117 22043 16175 22049
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 18141 22083 18199 22089
rect 18141 22080 18153 22083
rect 17276 22052 18153 22080
rect 17276 22040 17282 22052
rect 18141 22049 18153 22052
rect 18187 22049 18199 22083
rect 18141 22043 18199 22049
rect 20622 22040 20628 22092
rect 20680 22080 20686 22092
rect 20717 22083 20775 22089
rect 20717 22080 20729 22083
rect 20680 22052 20729 22080
rect 20680 22040 20686 22052
rect 20717 22049 20729 22052
rect 20763 22049 20775 22083
rect 20717 22043 20775 22049
rect 23658 22040 23664 22092
rect 23716 22080 23722 22092
rect 24397 22083 24455 22089
rect 24397 22080 24409 22083
rect 23716 22052 24409 22080
rect 23716 22040 23722 22052
rect 24397 22049 24409 22052
rect 24443 22049 24455 22083
rect 24397 22043 24455 22049
rect 25406 22040 25412 22092
rect 25464 22080 25470 22092
rect 26160 22080 26188 22179
rect 26234 22176 26240 22228
rect 26292 22176 26298 22228
rect 27890 22225 27896 22228
rect 27880 22219 27896 22225
rect 27880 22185 27892 22219
rect 27880 22179 27896 22185
rect 27890 22176 27896 22179
rect 27948 22176 27954 22228
rect 29362 22176 29368 22228
rect 29420 22176 29426 22228
rect 26418 22108 26424 22160
rect 26476 22148 26482 22160
rect 29380 22148 29408 22176
rect 26476 22120 26832 22148
rect 29380 22120 30236 22148
rect 26476 22108 26482 22120
rect 26804 22094 26832 22120
rect 26804 22089 26869 22094
rect 26697 22083 26755 22089
rect 26697 22080 26709 22083
rect 25464 22052 25912 22080
rect 26160 22052 26709 22080
rect 25464 22040 25470 22052
rect 14967 21984 15240 22012
rect 14967 21981 14979 21984
rect 14921 21975 14979 21981
rect 15286 21972 15292 22024
rect 15344 22012 15350 22024
rect 16393 22015 16451 22021
rect 16393 22012 16405 22015
rect 15344 21984 16405 22012
rect 15344 21972 15350 21984
rect 16393 21981 16405 21984
rect 16439 21981 16451 22015
rect 16393 21975 16451 21981
rect 23477 22015 23535 22021
rect 23477 21981 23489 22015
rect 23523 21981 23535 22015
rect 23477 21975 23535 21981
rect 11054 21904 11060 21956
rect 11112 21944 11118 21956
rect 15933 21947 15991 21953
rect 11112 21916 11270 21944
rect 11112 21904 11118 21916
rect 15933 21913 15945 21947
rect 15979 21944 15991 21947
rect 16942 21944 16948 21956
rect 15979 21916 16948 21944
rect 15979 21913 15991 21916
rect 15933 21907 15991 21913
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 18138 21944 18144 21956
rect 17894 21916 18144 21944
rect 18138 21904 18144 21916
rect 18196 21904 18202 21956
rect 22554 21944 22560 21956
rect 22218 21916 22560 21944
rect 22554 21904 22560 21916
rect 22612 21904 22618 21956
rect 5534 21876 5540 21888
rect 5368 21848 5540 21876
rect 5534 21836 5540 21848
rect 5592 21836 5598 21888
rect 5813 21879 5871 21885
rect 5813 21845 5825 21879
rect 5859 21876 5871 21879
rect 5994 21876 6000 21888
rect 5859 21848 6000 21876
rect 5859 21845 5871 21848
rect 5813 21839 5871 21845
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 6178 21836 6184 21888
rect 6236 21876 6242 21888
rect 6273 21879 6331 21885
rect 6273 21876 6285 21879
rect 6236 21848 6285 21876
rect 6236 21836 6242 21848
rect 6273 21845 6285 21848
rect 6319 21845 6331 21879
rect 6273 21839 6331 21845
rect 6454 21836 6460 21888
rect 6512 21836 6518 21888
rect 7098 21836 7104 21888
rect 7156 21836 7162 21888
rect 23492 21876 23520 21975
rect 23566 21972 23572 22024
rect 23624 21972 23630 22024
rect 23750 21972 23756 22024
rect 23808 21972 23814 22024
rect 24026 21972 24032 22024
rect 24084 22012 24090 22024
rect 24213 22015 24271 22021
rect 24213 22012 24225 22015
rect 24084 21984 24225 22012
rect 24084 21972 24090 21984
rect 24213 21981 24225 21984
rect 24259 21981 24271 22015
rect 24213 21975 24271 21981
rect 25884 21944 25912 22052
rect 26697 22049 26709 22052
rect 26743 22049 26755 22083
rect 26697 22043 26755 22049
rect 26789 22083 26869 22089
rect 26789 22049 26801 22083
rect 26835 22066 26869 22083
rect 26835 22049 26847 22066
rect 26789 22043 26847 22049
rect 26970 22040 26976 22092
rect 27028 22080 27034 22092
rect 27617 22083 27675 22089
rect 27617 22080 27629 22083
rect 27028 22052 27629 22080
rect 27028 22040 27034 22052
rect 27617 22049 27629 22052
rect 27663 22049 27675 22083
rect 27617 22043 27675 22049
rect 29270 22040 29276 22092
rect 29328 22080 29334 22092
rect 29549 22083 29607 22089
rect 29549 22080 29561 22083
rect 29328 22052 29561 22080
rect 29328 22040 29334 22052
rect 29549 22049 29561 22052
rect 29595 22049 29607 22083
rect 29549 22043 29607 22049
rect 26605 22015 26663 22021
rect 26605 21981 26617 22015
rect 26651 22012 26663 22015
rect 26878 22012 26884 22024
rect 26651 21984 26884 22012
rect 26651 21981 26663 21984
rect 26605 21975 26663 21981
rect 26878 21972 26884 21984
rect 26936 21972 26942 22024
rect 30006 21972 30012 22024
rect 30064 21972 30070 22024
rect 30208 22021 30236 22120
rect 30285 22083 30343 22089
rect 30285 22049 30297 22083
rect 30331 22080 30343 22083
rect 30742 22080 30748 22092
rect 30331 22052 30748 22080
rect 30331 22049 30343 22052
rect 30285 22043 30343 22049
rect 30742 22040 30748 22052
rect 30800 22040 30806 22092
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 21981 30251 22015
rect 30193 21975 30251 21981
rect 26142 21944 26148 21956
rect 25884 21930 26148 21944
rect 25898 21916 26148 21930
rect 26142 21904 26148 21916
rect 26200 21904 26206 21956
rect 27982 21904 27988 21956
rect 28040 21944 28046 21956
rect 28040 21916 28382 21944
rect 28040 21904 28046 21916
rect 25498 21876 25504 21888
rect 23492 21848 25504 21876
rect 25498 21836 25504 21848
rect 25556 21836 25562 21888
rect 1104 21786 37076 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 37076 21786
rect 1104 21712 37076 21734
rect 5534 21632 5540 21684
rect 5592 21672 5598 21684
rect 6733 21675 6791 21681
rect 6733 21672 6745 21675
rect 5592 21644 6745 21672
rect 5592 21632 5598 21644
rect 6733 21641 6745 21644
rect 6779 21641 6791 21675
rect 6733 21635 6791 21641
rect 8018 21632 8024 21684
rect 8076 21672 8082 21684
rect 9674 21672 9680 21684
rect 8076 21644 9680 21672
rect 8076 21632 8082 21644
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 9950 21632 9956 21684
rect 10008 21632 10014 21684
rect 10410 21632 10416 21684
rect 10468 21672 10474 21684
rect 10505 21675 10563 21681
rect 10505 21672 10517 21675
rect 10468 21644 10517 21672
rect 10468 21632 10474 21644
rect 10505 21641 10517 21644
rect 10551 21641 10563 21675
rect 10505 21635 10563 21641
rect 2958 21564 2964 21616
rect 3016 21604 3022 21616
rect 3694 21604 3700 21616
rect 3016 21576 3700 21604
rect 3016 21564 3022 21576
rect 3694 21564 3700 21576
rect 3752 21604 3758 21616
rect 3752 21576 3910 21604
rect 3752 21564 3758 21576
rect 8754 21564 8760 21616
rect 8812 21604 8818 21616
rect 9125 21607 9183 21613
rect 9125 21604 9137 21607
rect 8812 21576 9137 21604
rect 8812 21564 8818 21576
rect 9125 21573 9137 21576
rect 9171 21573 9183 21607
rect 9125 21567 9183 21573
rect 9217 21607 9275 21613
rect 9217 21573 9229 21607
rect 9263 21604 9275 21607
rect 9493 21607 9551 21613
rect 9493 21604 9505 21607
rect 9263 21576 9505 21604
rect 9263 21573 9275 21576
rect 9217 21567 9275 21573
rect 9493 21573 9505 21576
rect 9539 21604 9551 21607
rect 9582 21604 9588 21616
rect 9539 21576 9588 21604
rect 9539 21573 9551 21576
rect 9493 21567 9551 21573
rect 6454 21496 6460 21548
rect 6512 21536 6518 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6512 21508 6561 21536
rect 6512 21496 6518 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21536 6883 21539
rect 6914 21536 6920 21548
rect 6871 21508 6920 21536
rect 6871 21505 6883 21508
rect 6825 21499 6883 21505
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 9140 21536 9168 21567
rect 9582 21564 9588 21576
rect 9640 21564 9646 21616
rect 9677 21539 9735 21545
rect 9677 21536 9689 21539
rect 9140 21508 9689 21536
rect 9677 21505 9689 21508
rect 9723 21505 9735 21539
rect 9677 21499 9735 21505
rect 9769 21539 9827 21545
rect 9769 21505 9781 21539
rect 9815 21505 9827 21539
rect 9769 21499 9827 21505
rect 1394 21428 1400 21480
rect 1452 21468 1458 21480
rect 3145 21471 3203 21477
rect 3145 21468 3157 21471
rect 1452 21440 3157 21468
rect 1452 21428 1458 21440
rect 3145 21437 3157 21440
rect 3191 21437 3203 21471
rect 3145 21431 3203 21437
rect 3418 21428 3424 21480
rect 3476 21428 3482 21480
rect 9122 21428 9128 21480
rect 9180 21468 9186 21480
rect 9401 21471 9459 21477
rect 9401 21468 9413 21471
rect 9180 21440 9413 21468
rect 9180 21428 9186 21440
rect 9401 21437 9413 21440
rect 9447 21437 9459 21471
rect 9401 21431 9459 21437
rect 8202 21360 8208 21412
rect 8260 21400 8266 21412
rect 8849 21403 8907 21409
rect 8849 21400 8861 21403
rect 8260 21372 8861 21400
rect 8260 21360 8266 21372
rect 8849 21369 8861 21372
rect 8895 21400 8907 21403
rect 9306 21400 9312 21412
rect 8895 21372 9312 21400
rect 8895 21369 8907 21372
rect 8849 21363 8907 21369
rect 9306 21360 9312 21372
rect 9364 21400 9370 21412
rect 9784 21400 9812 21499
rect 28350 21496 28356 21548
rect 28408 21536 28414 21548
rect 28537 21539 28595 21545
rect 28537 21536 28549 21539
rect 28408 21508 28549 21536
rect 28408 21496 28414 21508
rect 28537 21505 28549 21508
rect 28583 21505 28595 21539
rect 28537 21499 28595 21505
rect 28629 21539 28687 21545
rect 28629 21505 28641 21539
rect 28675 21536 28687 21539
rect 29546 21536 29552 21548
rect 28675 21508 29552 21536
rect 28675 21505 28687 21508
rect 28629 21499 28687 21505
rect 29546 21496 29552 21508
rect 29604 21536 29610 21548
rect 30653 21539 30711 21545
rect 30653 21536 30665 21539
rect 29604 21508 30665 21536
rect 29604 21496 29610 21508
rect 30653 21505 30665 21508
rect 30699 21505 30711 21539
rect 31481 21539 31539 21545
rect 31481 21536 31493 21539
rect 30653 21499 30711 21505
rect 30760 21508 31493 21536
rect 9950 21428 9956 21480
rect 10008 21468 10014 21480
rect 10597 21471 10655 21477
rect 10597 21468 10609 21471
rect 10008 21440 10609 21468
rect 10008 21428 10014 21440
rect 10597 21437 10609 21440
rect 10643 21437 10655 21471
rect 10597 21431 10655 21437
rect 10778 21428 10784 21480
rect 10836 21428 10842 21480
rect 28718 21428 28724 21480
rect 28776 21428 28782 21480
rect 30558 21428 30564 21480
rect 30616 21468 30622 21480
rect 30760 21477 30788 21508
rect 31481 21505 31493 21508
rect 31527 21505 31539 21539
rect 32677 21539 32735 21545
rect 32677 21536 32689 21539
rect 31481 21499 31539 21505
rect 31588 21508 32689 21536
rect 31588 21480 31616 21508
rect 32677 21505 32689 21508
rect 32723 21505 32735 21539
rect 32677 21499 32735 21505
rect 30745 21471 30803 21477
rect 30745 21468 30757 21471
rect 30616 21440 30757 21468
rect 30616 21428 30622 21440
rect 30745 21437 30757 21440
rect 30791 21437 30803 21471
rect 30745 21431 30803 21437
rect 30837 21471 30895 21477
rect 30837 21437 30849 21471
rect 30883 21437 30895 21471
rect 30837 21431 30895 21437
rect 9364 21372 9812 21400
rect 28736 21400 28764 21428
rect 30852 21400 30880 21431
rect 31570 21428 31576 21480
rect 31628 21428 31634 21480
rect 31665 21471 31723 21477
rect 31665 21437 31677 21471
rect 31711 21437 31723 21471
rect 31665 21431 31723 21437
rect 31680 21400 31708 21431
rect 32766 21428 32772 21480
rect 32824 21428 32830 21480
rect 32861 21471 32919 21477
rect 32861 21437 32873 21471
rect 32907 21437 32919 21471
rect 32861 21431 32919 21437
rect 32876 21400 32904 21431
rect 28736 21372 31708 21400
rect 9364 21360 9370 21372
rect 31680 21344 31708 21372
rect 32048 21372 32904 21400
rect 3878 21292 3884 21344
rect 3936 21332 3942 21344
rect 4706 21332 4712 21344
rect 3936 21304 4712 21332
rect 3936 21292 3942 21304
rect 4706 21292 4712 21304
rect 4764 21332 4770 21344
rect 4893 21335 4951 21341
rect 4893 21332 4905 21335
rect 4764 21304 4905 21332
rect 4764 21292 4770 21304
rect 4893 21301 4905 21304
rect 4939 21301 4951 21335
rect 4893 21295 4951 21301
rect 6086 21292 6092 21344
rect 6144 21332 6150 21344
rect 6365 21335 6423 21341
rect 6365 21332 6377 21335
rect 6144 21304 6377 21332
rect 6144 21292 6150 21304
rect 6365 21301 6377 21304
rect 6411 21301 6423 21335
rect 6365 21295 6423 21301
rect 7466 21292 7472 21344
rect 7524 21332 7530 21344
rect 8018 21332 8024 21344
rect 7524 21304 8024 21332
rect 7524 21292 7530 21304
rect 8018 21292 8024 21304
rect 8076 21292 8082 21344
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 9493 21335 9551 21341
rect 9493 21332 9505 21335
rect 9088 21304 9505 21332
rect 9088 21292 9094 21304
rect 9493 21301 9505 21304
rect 9539 21301 9551 21335
rect 9493 21295 9551 21301
rect 10137 21335 10195 21341
rect 10137 21301 10149 21335
rect 10183 21332 10195 21335
rect 10318 21332 10324 21344
rect 10183 21304 10324 21332
rect 10183 21301 10195 21304
rect 10137 21295 10195 21301
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 27614 21292 27620 21344
rect 27672 21332 27678 21344
rect 28169 21335 28227 21341
rect 28169 21332 28181 21335
rect 27672 21304 28181 21332
rect 27672 21292 27678 21304
rect 28169 21301 28181 21304
rect 28215 21301 28227 21335
rect 28169 21295 28227 21301
rect 30285 21335 30343 21341
rect 30285 21301 30297 21335
rect 30331 21332 30343 21335
rect 31018 21332 31024 21344
rect 30331 21304 31024 21332
rect 30331 21301 30343 21304
rect 30285 21295 30343 21301
rect 31018 21292 31024 21304
rect 31076 21292 31082 21344
rect 31110 21292 31116 21344
rect 31168 21292 31174 21344
rect 31662 21292 31668 21344
rect 31720 21332 31726 21344
rect 32048 21332 32076 21372
rect 31720 21304 32076 21332
rect 32309 21335 32367 21341
rect 31720 21292 31726 21304
rect 32309 21301 32321 21335
rect 32355 21332 32367 21335
rect 32950 21332 32956 21344
rect 32355 21304 32956 21332
rect 32355 21301 32367 21304
rect 32309 21295 32367 21301
rect 32950 21292 32956 21304
rect 33008 21292 33014 21344
rect 1104 21242 37076 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 37076 21242
rect 1104 21168 37076 21190
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 4065 21131 4123 21137
rect 4065 21128 4077 21131
rect 3476 21100 4077 21128
rect 3476 21088 3482 21100
rect 4065 21097 4077 21100
rect 4111 21097 4123 21131
rect 4065 21091 4123 21097
rect 4617 21131 4675 21137
rect 4617 21097 4629 21131
rect 4663 21128 4675 21131
rect 5534 21128 5540 21140
rect 4663 21100 5540 21128
rect 4663 21097 4675 21100
rect 4617 21091 4675 21097
rect 5534 21088 5540 21100
rect 5592 21088 5598 21140
rect 7006 21088 7012 21140
rect 7064 21128 7070 21140
rect 7064 21100 7880 21128
rect 7064 21088 7070 21100
rect 7285 21063 7343 21069
rect 7285 21060 7297 21063
rect 6932 21032 7297 21060
rect 6932 21004 6960 21032
rect 7285 21029 7297 21032
rect 7331 21029 7343 21063
rect 7285 21023 7343 21029
rect 1394 20952 1400 21004
rect 1452 20952 1458 21004
rect 4614 20992 4620 21004
rect 3804 20964 4620 20992
rect 3804 20933 3832 20964
rect 4614 20952 4620 20964
rect 4672 20952 4678 21004
rect 6086 20952 6092 21004
rect 6144 20952 6150 21004
rect 6914 20952 6920 21004
rect 6972 20952 6978 21004
rect 7006 20952 7012 21004
rect 7064 20952 7070 21004
rect 7852 21001 7880 21100
rect 8294 21088 8300 21140
rect 8352 21128 8358 21140
rect 8352 21100 9260 21128
rect 8352 21088 8358 21100
rect 7926 21020 7932 21072
rect 7984 21060 7990 21072
rect 9122 21060 9128 21072
rect 7984 21032 9128 21060
rect 7984 21020 7990 21032
rect 7837 20995 7895 21001
rect 7300 20964 7696 20992
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 3878 20884 3884 20936
rect 3936 20884 3942 20936
rect 4062 20884 4068 20936
rect 4120 20884 4126 20936
rect 6362 20884 6368 20936
rect 6420 20884 6426 20936
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20924 6883 20927
rect 7098 20924 7104 20936
rect 6871 20896 7104 20924
rect 6871 20893 6883 20896
rect 6825 20887 6883 20893
rect 7098 20884 7104 20896
rect 7156 20924 7162 20936
rect 7300 20933 7328 20964
rect 7285 20927 7343 20933
rect 7285 20924 7297 20927
rect 7156 20896 7297 20924
rect 7156 20884 7162 20896
rect 7285 20893 7297 20896
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 7466 20884 7472 20936
rect 7524 20884 7530 20936
rect 7668 20933 7696 20964
rect 7837 20961 7849 20995
rect 7883 20992 7895 20995
rect 8202 20992 8208 21004
rect 7883 20964 8208 20992
rect 7883 20961 7895 20964
rect 7837 20955 7895 20961
rect 8202 20952 8208 20964
rect 8260 20992 8266 21004
rect 8260 20964 8432 20992
rect 8260 20952 8266 20964
rect 7653 20927 7711 20933
rect 7653 20893 7665 20927
rect 7699 20924 7711 20927
rect 7926 20924 7932 20936
rect 7699 20896 7932 20924
rect 7699 20893 7711 20896
rect 7653 20887 7711 20893
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 8018 20884 8024 20936
rect 8076 20884 8082 20936
rect 8294 20884 8300 20936
rect 8352 20884 8358 20936
rect 8404 20933 8432 20964
rect 8588 20933 8616 21032
rect 9122 21020 9128 21032
rect 9180 21020 9186 21072
rect 9232 21060 9260 21100
rect 9950 21088 9956 21140
rect 10008 21088 10014 21140
rect 10410 21128 10416 21140
rect 10060 21100 10416 21128
rect 9858 21060 9864 21072
rect 9232 21032 9864 21060
rect 8754 20952 8760 21004
rect 8812 20992 8818 21004
rect 9033 20995 9091 21001
rect 9033 20992 9045 20995
rect 8812 20964 9045 20992
rect 8812 20952 8818 20964
rect 9033 20961 9045 20964
rect 9079 20961 9091 20995
rect 9033 20955 9091 20961
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20893 8447 20927
rect 8389 20887 8447 20893
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20893 8631 20927
rect 8573 20887 8631 20893
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20924 8999 20927
rect 9232 20924 9260 21032
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 10060 21060 10088 21100
rect 10410 21088 10416 21100
rect 10468 21088 10474 21140
rect 10778 21088 10784 21140
rect 10836 21128 10842 21140
rect 11793 21131 11851 21137
rect 11793 21128 11805 21131
rect 10836 21100 11805 21128
rect 10836 21088 10842 21100
rect 11793 21097 11805 21100
rect 11839 21097 11851 21131
rect 11793 21091 11851 21097
rect 29546 21088 29552 21140
rect 29604 21088 29610 21140
rect 31481 21131 31539 21137
rect 31481 21097 31493 21131
rect 31527 21128 31539 21131
rect 31570 21128 31576 21140
rect 31527 21100 31576 21128
rect 31527 21097 31539 21100
rect 31481 21091 31539 21097
rect 31570 21088 31576 21100
rect 31628 21088 31634 21140
rect 32766 21088 32772 21140
rect 32824 21128 32830 21140
rect 32824 21100 34100 21128
rect 32824 21088 32830 21100
rect 23566 21060 23572 21072
rect 9968 21032 10088 21060
rect 21376 21032 23572 21060
rect 9306 20952 9312 21004
rect 9364 20952 9370 21004
rect 8987 20896 9260 20924
rect 9401 20927 9459 20933
rect 8987 20893 8999 20896
rect 8941 20887 8999 20893
rect 9401 20893 9413 20927
rect 9447 20924 9459 20927
rect 9582 20924 9588 20936
rect 9447 20896 9588 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 9582 20884 9588 20896
rect 9640 20884 9646 20936
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 9968 20933 9996 21032
rect 10042 20952 10048 21004
rect 10100 20952 10106 21004
rect 10318 20952 10324 21004
rect 10376 20952 10382 21004
rect 21376 21001 21404 21032
rect 23566 21020 23572 21032
rect 23624 21020 23630 21072
rect 21361 20995 21419 21001
rect 21361 20961 21373 20995
rect 21407 20961 21419 20995
rect 23658 20992 23664 21004
rect 21361 20955 21419 20961
rect 22756 20964 23664 20992
rect 9769 20927 9827 20933
rect 9769 20924 9781 20927
rect 9732 20896 9781 20924
rect 9732 20884 9738 20896
rect 9769 20893 9781 20896
rect 9815 20893 9827 20927
rect 9769 20887 9827 20893
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20893 10011 20927
rect 9953 20887 10011 20893
rect 16761 20927 16819 20933
rect 16761 20893 16773 20927
rect 16807 20924 16819 20927
rect 16850 20924 16856 20936
rect 16807 20896 16856 20924
rect 16807 20893 16819 20896
rect 16761 20887 16819 20893
rect 16850 20884 16856 20896
rect 16908 20884 16914 20936
rect 22756 20933 22784 20964
rect 23658 20952 23664 20964
rect 23716 20992 23722 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 23716 20964 25145 20992
rect 23716 20952 23722 20964
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 27614 20952 27620 21004
rect 27672 20952 27678 21004
rect 27982 20952 27988 21004
rect 28040 20992 28046 21004
rect 28040 20964 28948 20992
rect 28040 20952 28046 20964
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20893 22615 20927
rect 22557 20887 22615 20893
rect 22741 20927 22799 20933
rect 22741 20893 22753 20927
rect 22787 20893 22799 20927
rect 22741 20887 22799 20893
rect 1670 20816 1676 20868
rect 1728 20816 1734 20868
rect 2958 20856 2964 20868
rect 2898 20828 2964 20856
rect 2958 20816 2964 20828
rect 3016 20856 3022 20868
rect 4798 20856 4804 20868
rect 3016 20828 4804 20856
rect 3016 20816 3022 20828
rect 4798 20816 4804 20828
rect 4856 20856 4862 20868
rect 6380 20856 6408 20884
rect 10042 20856 10048 20868
rect 4856 20828 4922 20856
rect 6380 20828 10048 20856
rect 4856 20816 4862 20828
rect 10042 20816 10048 20828
rect 10100 20816 10106 20868
rect 11054 20816 11060 20868
rect 11112 20816 11118 20868
rect 16022 20816 16028 20868
rect 16080 20856 16086 20868
rect 16485 20859 16543 20865
rect 16080 20828 16252 20856
rect 16080 20816 16086 20828
rect 3142 20748 3148 20800
rect 3200 20748 3206 20800
rect 6457 20791 6515 20797
rect 6457 20757 6469 20791
rect 6503 20788 6515 20791
rect 6638 20788 6644 20800
rect 6503 20760 6644 20788
rect 6503 20757 6515 20760
rect 6457 20751 6515 20757
rect 6638 20748 6644 20760
rect 6696 20748 6702 20800
rect 7745 20791 7803 20797
rect 7745 20757 7757 20791
rect 7791 20788 7803 20791
rect 7834 20788 7840 20800
rect 7791 20760 7840 20788
rect 7791 20757 7803 20760
rect 7745 20751 7803 20757
rect 7834 20748 7840 20760
rect 7892 20748 7898 20800
rect 7929 20791 7987 20797
rect 7929 20757 7941 20791
rect 7975 20788 7987 20791
rect 8294 20788 8300 20800
rect 7975 20760 8300 20788
rect 7975 20757 7987 20760
rect 7929 20751 7987 20757
rect 8294 20748 8300 20760
rect 8352 20748 8358 20800
rect 8757 20791 8815 20797
rect 8757 20757 8769 20791
rect 8803 20788 8815 20791
rect 8938 20788 8944 20800
rect 8803 20760 8944 20788
rect 8803 20757 8815 20760
rect 8757 20751 8815 20757
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 9122 20748 9128 20800
rect 9180 20748 9186 20800
rect 9585 20791 9643 20797
rect 9585 20757 9597 20791
rect 9631 20788 9643 20791
rect 9766 20788 9772 20800
rect 9631 20760 9772 20788
rect 9631 20757 9643 20760
rect 9585 20751 9643 20757
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 15013 20791 15071 20797
rect 15013 20757 15025 20791
rect 15059 20788 15071 20791
rect 16114 20788 16120 20800
rect 15059 20760 16120 20788
rect 15059 20757 15071 20760
rect 15013 20751 15071 20757
rect 16114 20748 16120 20760
rect 16172 20748 16178 20800
rect 16224 20788 16252 20828
rect 16485 20825 16497 20859
rect 16531 20856 16543 20859
rect 16574 20856 16580 20868
rect 16531 20828 16580 20856
rect 16531 20825 16543 20828
rect 16485 20819 16543 20825
rect 16574 20816 16580 20828
rect 16632 20816 16638 20868
rect 17126 20816 17132 20868
rect 17184 20816 17190 20868
rect 18138 20816 18144 20868
rect 18196 20816 18202 20868
rect 22094 20816 22100 20868
rect 22152 20816 22158 20868
rect 22572 20856 22600 20887
rect 22830 20884 22836 20936
rect 22888 20884 22894 20936
rect 24857 20927 24915 20933
rect 24857 20924 24869 20927
rect 24320 20896 24869 20924
rect 24320 20856 24348 20896
rect 24857 20893 24869 20896
rect 24903 20893 24915 20927
rect 24857 20887 24915 20893
rect 22572 20828 24348 20856
rect 24397 20859 24455 20865
rect 24397 20825 24409 20859
rect 24443 20825 24455 20859
rect 24872 20856 24900 20887
rect 24946 20884 24952 20936
rect 25004 20924 25010 20936
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 25004 20896 25053 20924
rect 25004 20884 25010 20896
rect 25041 20893 25053 20896
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 26970 20884 26976 20936
rect 27028 20924 27034 20936
rect 27341 20927 27399 20933
rect 27341 20924 27353 20927
rect 27028 20896 27353 20924
rect 27028 20884 27034 20896
rect 27341 20893 27353 20896
rect 27387 20893 27399 20927
rect 27341 20887 27399 20893
rect 27062 20856 27068 20868
rect 24872 20828 27068 20856
rect 24397 20819 24455 20825
rect 17954 20788 17960 20800
rect 16224 20760 17960 20788
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 18046 20748 18052 20800
rect 18104 20788 18110 20800
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18104 20760 18613 20788
rect 18104 20748 18110 20760
rect 18601 20757 18613 20760
rect 18647 20757 18659 20791
rect 18601 20751 18659 20757
rect 20714 20748 20720 20800
rect 20772 20748 20778 20800
rect 20806 20748 20812 20800
rect 20864 20788 20870 20800
rect 21085 20791 21143 20797
rect 21085 20788 21097 20791
rect 20864 20760 21097 20788
rect 20864 20748 20870 20760
rect 21085 20757 21097 20760
rect 21131 20757 21143 20791
rect 21085 20751 21143 20757
rect 21177 20791 21235 20797
rect 21177 20757 21189 20791
rect 21223 20788 21235 20791
rect 22830 20788 22836 20800
rect 21223 20760 22836 20788
rect 21223 20757 21235 20760
rect 21177 20751 21235 20757
rect 22830 20748 22836 20760
rect 22888 20748 22894 20800
rect 24412 20788 24440 20819
rect 27062 20816 27068 20828
rect 27120 20816 27126 20868
rect 28920 20856 28948 20964
rect 31018 20952 31024 21004
rect 31076 20952 31082 21004
rect 31297 20995 31355 21001
rect 31297 20961 31309 20995
rect 31343 20992 31355 20995
rect 31754 20992 31760 21004
rect 31343 20964 31760 20992
rect 31343 20961 31355 20964
rect 31297 20955 31355 20961
rect 31754 20952 31760 20964
rect 31812 20992 31818 21004
rect 33229 20995 33287 21001
rect 33229 20992 33241 20995
rect 31812 20964 33241 20992
rect 31812 20952 31818 20964
rect 33229 20961 33241 20964
rect 33275 20992 33287 20995
rect 33275 20964 33916 20992
rect 33275 20961 33287 20964
rect 33229 20955 33287 20961
rect 33410 20884 33416 20936
rect 33468 20924 33474 20936
rect 33781 20927 33839 20933
rect 33781 20924 33793 20927
rect 33468 20896 33793 20924
rect 33468 20884 33474 20896
rect 33781 20893 33793 20896
rect 33827 20893 33839 20927
rect 33781 20887 33839 20893
rect 30742 20856 30748 20868
rect 28842 20828 29224 20856
rect 30590 20828 30748 20856
rect 25130 20788 25136 20800
rect 24412 20760 25136 20788
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 28350 20748 28356 20800
rect 28408 20788 28414 20800
rect 29089 20791 29147 20797
rect 29089 20788 29101 20791
rect 28408 20760 29101 20788
rect 28408 20748 28414 20760
rect 29089 20757 29101 20760
rect 29135 20757 29147 20791
rect 29196 20788 29224 20828
rect 30668 20788 30696 20828
rect 30742 20816 30748 20828
rect 30800 20856 30806 20868
rect 32858 20856 32864 20868
rect 30800 20828 30972 20856
rect 32522 20828 32864 20856
rect 30800 20816 30806 20828
rect 29196 20760 30696 20788
rect 30944 20788 30972 20828
rect 32600 20788 32628 20828
rect 32858 20816 32864 20828
rect 32916 20816 32922 20868
rect 32950 20816 32956 20868
rect 33008 20816 33014 20868
rect 33321 20859 33379 20865
rect 33321 20825 33333 20859
rect 33367 20856 33379 20859
rect 33502 20856 33508 20868
rect 33367 20828 33508 20856
rect 33367 20825 33379 20828
rect 33321 20819 33379 20825
rect 33502 20816 33508 20828
rect 33560 20816 33566 20868
rect 33888 20856 33916 20964
rect 33962 20884 33968 20936
rect 34020 20884 34026 20936
rect 34072 20933 34100 21100
rect 34057 20927 34115 20933
rect 34057 20893 34069 20927
rect 34103 20893 34115 20927
rect 34057 20887 34115 20893
rect 34146 20884 34152 20936
rect 34204 20924 34210 20936
rect 34701 20927 34759 20933
rect 34701 20924 34713 20927
rect 34204 20896 34713 20924
rect 34204 20884 34210 20896
rect 34701 20893 34713 20896
rect 34747 20893 34759 20927
rect 34701 20887 34759 20893
rect 34164 20856 34192 20884
rect 33888 20828 34192 20856
rect 34974 20816 34980 20868
rect 35032 20816 35038 20868
rect 35434 20816 35440 20868
rect 35492 20816 35498 20868
rect 30944 20760 32628 20788
rect 29089 20751 29147 20757
rect 33962 20748 33968 20800
rect 34020 20788 34026 20800
rect 34422 20788 34428 20800
rect 34020 20760 34428 20788
rect 34020 20748 34026 20760
rect 34422 20748 34428 20760
rect 34480 20788 34486 20800
rect 36449 20791 36507 20797
rect 36449 20788 36461 20791
rect 34480 20760 36461 20788
rect 34480 20748 34486 20760
rect 36449 20757 36461 20760
rect 36495 20757 36507 20791
rect 36449 20751 36507 20757
rect 1104 20698 37076 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 37076 20698
rect 1104 20624 37076 20646
rect 4798 20544 4804 20596
rect 4856 20584 4862 20596
rect 6822 20584 6828 20596
rect 4856 20556 6828 20584
rect 4856 20544 4862 20556
rect 6822 20544 6828 20556
rect 6880 20584 6886 20596
rect 8113 20587 8171 20593
rect 6880 20556 7052 20584
rect 6880 20544 6886 20556
rect 6638 20476 6644 20528
rect 6696 20476 6702 20528
rect 7024 20516 7052 20556
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8202 20584 8208 20596
rect 8159 20556 8208 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 8294 20544 8300 20596
rect 8352 20584 8358 20596
rect 8665 20587 8723 20593
rect 8665 20584 8677 20587
rect 8352 20556 8677 20584
rect 8352 20544 8358 20556
rect 8665 20553 8677 20556
rect 8711 20553 8723 20587
rect 8665 20547 8723 20553
rect 7024 20488 7130 20516
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20448 2283 20451
rect 3142 20448 3148 20460
rect 2271 20420 3148 20448
rect 2271 20417 2283 20420
rect 2225 20411 2283 20417
rect 3142 20408 3148 20420
rect 3200 20408 3206 20460
rect 8110 20408 8116 20460
rect 8168 20448 8174 20460
rect 8573 20451 8631 20457
rect 8573 20448 8585 20451
rect 8168 20420 8585 20448
rect 8168 20408 8174 20420
rect 8573 20417 8585 20420
rect 8619 20417 8631 20451
rect 8680 20448 8708 20547
rect 9582 20544 9588 20596
rect 9640 20544 9646 20596
rect 10042 20544 10048 20596
rect 10100 20584 10106 20596
rect 10100 20556 11284 20584
rect 10100 20544 10106 20556
rect 11054 20516 11060 20528
rect 10626 20488 11060 20516
rect 11054 20476 11060 20488
rect 11112 20476 11118 20528
rect 11256 20516 11284 20556
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 20456 20556 22508 20584
rect 15930 20516 15936 20528
rect 11256 20488 11376 20516
rect 15318 20488 15936 20516
rect 8680 20420 8892 20448
rect 8573 20411 8631 20417
rect 1670 20340 1676 20392
rect 1728 20380 1734 20392
rect 1857 20383 1915 20389
rect 1857 20380 1869 20383
rect 1728 20352 1869 20380
rect 1728 20340 1734 20352
rect 1857 20349 1869 20352
rect 1903 20349 1915 20383
rect 1857 20343 1915 20349
rect 2317 20383 2375 20389
rect 2317 20349 2329 20383
rect 2363 20380 2375 20383
rect 2958 20380 2964 20392
rect 2363 20352 2964 20380
rect 2363 20349 2375 20352
rect 2317 20343 2375 20349
rect 2958 20340 2964 20352
rect 3016 20340 3022 20392
rect 6362 20340 6368 20392
rect 6420 20340 6426 20392
rect 8754 20340 8760 20392
rect 8812 20340 8818 20392
rect 8864 20380 8892 20420
rect 8938 20408 8944 20460
rect 8996 20448 9002 20460
rect 11348 20457 11376 20488
rect 15930 20476 15936 20488
rect 15988 20476 15994 20528
rect 17126 20476 17132 20528
rect 17184 20516 17190 20528
rect 17497 20519 17555 20525
rect 17497 20516 17509 20519
rect 17184 20488 17509 20516
rect 17184 20476 17190 20488
rect 17497 20485 17509 20488
rect 17543 20485 17555 20519
rect 17497 20479 17555 20485
rect 19242 20476 19248 20528
rect 19300 20516 19306 20528
rect 20456 20516 20484 20556
rect 19300 20488 20562 20516
rect 19300 20476 19306 20488
rect 22094 20476 22100 20528
rect 22152 20476 22158 20528
rect 22480 20516 22508 20556
rect 22830 20544 22836 20596
rect 22888 20584 22894 20596
rect 23569 20587 23627 20593
rect 23569 20584 23581 20587
rect 22888 20556 23581 20584
rect 22888 20544 22894 20556
rect 23569 20553 23581 20556
rect 23615 20553 23627 20587
rect 23569 20547 23627 20553
rect 23658 20544 23664 20596
rect 23716 20544 23722 20596
rect 26142 20584 26148 20596
rect 23860 20556 26148 20584
rect 22554 20516 22560 20528
rect 22480 20488 22560 20516
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 23860 20516 23888 20556
rect 24780 20516 24808 20556
rect 26142 20544 26148 20556
rect 26200 20544 26206 20596
rect 26970 20544 26976 20596
rect 27028 20584 27034 20596
rect 29733 20587 29791 20593
rect 27028 20556 28672 20584
rect 27028 20544 27034 20556
rect 23322 20502 23888 20516
rect 23308 20488 23888 20502
rect 24702 20488 24808 20516
rect 9217 20451 9275 20457
rect 9217 20448 9229 20451
rect 8996 20420 9229 20448
rect 8996 20408 9002 20420
rect 9217 20417 9229 20420
rect 9263 20417 9275 20451
rect 9217 20411 9275 20417
rect 11333 20451 11391 20457
rect 11333 20417 11345 20451
rect 11379 20417 11391 20451
rect 11333 20411 11391 20417
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15620 20420 16037 20448
rect 15620 20408 15626 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20417 18015 20451
rect 17957 20411 18015 20417
rect 18141 20451 18199 20457
rect 18141 20417 18153 20451
rect 18187 20448 18199 20451
rect 18414 20448 18420 20460
rect 18187 20420 18420 20448
rect 18187 20417 18199 20420
rect 18141 20411 18199 20417
rect 9033 20383 9091 20389
rect 9033 20380 9045 20383
rect 8864 20352 9045 20380
rect 9033 20349 9045 20352
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 11054 20340 11060 20392
rect 11112 20340 11118 20392
rect 13814 20340 13820 20392
rect 13872 20340 13878 20392
rect 14093 20383 14151 20389
rect 14093 20349 14105 20383
rect 14139 20380 14151 20383
rect 14139 20352 15700 20380
rect 14139 20349 14151 20352
rect 14093 20343 14151 20349
rect 7742 20272 7748 20324
rect 7800 20312 7806 20324
rect 8205 20315 8263 20321
rect 8205 20312 8217 20315
rect 7800 20284 8217 20312
rect 7800 20272 7806 20284
rect 8205 20281 8217 20284
rect 8251 20281 8263 20315
rect 8205 20275 8263 20281
rect 9401 20315 9459 20321
rect 9401 20281 9413 20315
rect 9447 20312 9459 20315
rect 9674 20312 9680 20324
rect 9447 20284 9680 20312
rect 9447 20281 9459 20284
rect 9401 20275 9459 20281
rect 9674 20272 9680 20284
rect 9732 20272 9738 20324
rect 15672 20321 15700 20352
rect 16298 20340 16304 20392
rect 16356 20340 16362 20392
rect 15657 20315 15715 20321
rect 15657 20281 15669 20315
rect 15703 20281 15715 20315
rect 17972 20312 18000 20411
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 18046 20340 18052 20392
rect 18104 20380 18110 20392
rect 18233 20383 18291 20389
rect 18233 20380 18245 20383
rect 18104 20352 18245 20380
rect 18104 20340 18110 20352
rect 18233 20349 18245 20352
rect 18279 20349 18291 20383
rect 18233 20343 18291 20349
rect 19797 20383 19855 20389
rect 19797 20349 19809 20383
rect 19843 20349 19855 20383
rect 19797 20343 19855 20349
rect 20073 20383 20131 20389
rect 20073 20349 20085 20383
rect 20119 20380 20131 20383
rect 20714 20380 20720 20392
rect 20119 20352 20720 20380
rect 20119 20349 20131 20352
rect 20073 20343 20131 20349
rect 19150 20312 19156 20324
rect 17972 20284 19156 20312
rect 15657 20275 15715 20281
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 15562 20204 15568 20256
rect 15620 20204 15626 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19812 20244 19840 20343
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 20806 20340 20812 20392
rect 20864 20380 20870 20392
rect 21545 20383 21603 20389
rect 21545 20380 21557 20383
rect 20864 20352 21557 20380
rect 20864 20340 20870 20352
rect 21545 20349 21557 20352
rect 21591 20349 21603 20383
rect 21545 20343 21603 20349
rect 21821 20383 21879 20389
rect 21821 20349 21833 20383
rect 21867 20349 21879 20383
rect 21821 20343 21879 20349
rect 21836 20312 21864 20343
rect 22554 20340 22560 20392
rect 22612 20380 22618 20392
rect 23308 20380 23336 20488
rect 25130 20476 25136 20528
rect 25188 20476 25194 20528
rect 26237 20519 26295 20525
rect 26237 20485 26249 20519
rect 26283 20516 26295 20519
rect 26283 20488 27016 20516
rect 26283 20485 26295 20488
rect 26237 20479 26295 20485
rect 26145 20451 26203 20457
rect 26145 20417 26157 20451
rect 26191 20448 26203 20451
rect 26510 20448 26516 20460
rect 26191 20420 26516 20448
rect 26191 20417 26203 20420
rect 26145 20411 26203 20417
rect 26510 20408 26516 20420
rect 26568 20408 26574 20460
rect 22612 20352 23336 20380
rect 22612 20340 22618 20352
rect 23658 20340 23664 20392
rect 23716 20380 23722 20392
rect 23716 20352 25360 20380
rect 23716 20340 23722 20352
rect 21100 20284 21864 20312
rect 25332 20312 25360 20352
rect 25406 20340 25412 20392
rect 25464 20340 25470 20392
rect 26329 20383 26387 20389
rect 26329 20380 26341 20383
rect 26206 20352 26341 20380
rect 26206 20312 26234 20352
rect 26329 20349 26341 20352
rect 26375 20349 26387 20383
rect 26329 20343 26387 20349
rect 25332 20284 26234 20312
rect 21100 20244 21128 20284
rect 19576 20216 21128 20244
rect 21836 20244 21864 20284
rect 22278 20244 22284 20256
rect 21836 20216 22284 20244
rect 19576 20204 19582 20216
rect 22278 20204 22284 20216
rect 22336 20204 22342 20256
rect 25038 20204 25044 20256
rect 25096 20244 25102 20256
rect 26988 20253 27016 20488
rect 27982 20476 27988 20528
rect 28040 20476 28046 20528
rect 28644 20516 28672 20556
rect 29733 20553 29745 20587
rect 29779 20584 29791 20587
rect 30558 20584 30564 20596
rect 29779 20556 30564 20584
rect 29779 20553 29791 20556
rect 29733 20547 29791 20553
rect 30558 20544 30564 20556
rect 30616 20544 30622 20596
rect 32309 20587 32367 20593
rect 32309 20553 32321 20587
rect 32355 20584 32367 20587
rect 32766 20584 32772 20596
rect 32355 20556 32772 20584
rect 32355 20553 32367 20556
rect 32309 20547 32367 20553
rect 32766 20544 32772 20556
rect 32824 20544 32830 20596
rect 32858 20544 32864 20596
rect 32916 20584 32922 20596
rect 35434 20584 35440 20596
rect 32916 20556 35440 20584
rect 32916 20544 32922 20556
rect 28644 20488 28764 20516
rect 28736 20457 28764 20488
rect 30742 20476 30748 20528
rect 30800 20476 30806 20528
rect 31110 20476 31116 20528
rect 31168 20516 31174 20528
rect 31205 20519 31263 20525
rect 31205 20516 31217 20519
rect 31168 20488 31217 20516
rect 31168 20476 31174 20488
rect 31205 20485 31217 20488
rect 31251 20485 31263 20519
rect 31205 20479 31263 20485
rect 33318 20476 33324 20528
rect 33376 20516 33382 20528
rect 33428 20516 33456 20556
rect 35434 20544 35440 20556
rect 35492 20544 35498 20596
rect 33376 20488 33456 20516
rect 33376 20476 33382 20488
rect 33502 20476 33508 20528
rect 33560 20516 33566 20528
rect 33781 20519 33839 20525
rect 33781 20516 33793 20519
rect 33560 20488 33793 20516
rect 33560 20476 33566 20488
rect 33781 20485 33793 20488
rect 33827 20485 33839 20519
rect 33781 20479 33839 20485
rect 34974 20476 34980 20528
rect 35032 20516 35038 20528
rect 35161 20519 35219 20525
rect 35161 20516 35173 20519
rect 35032 20488 35173 20516
rect 35032 20476 35038 20488
rect 35161 20485 35173 20488
rect 35207 20485 35219 20519
rect 35161 20479 35219 20485
rect 28721 20451 28779 20457
rect 28721 20417 28733 20451
rect 28767 20417 28779 20451
rect 28721 20411 28779 20417
rect 34057 20451 34115 20457
rect 34057 20417 34069 20451
rect 34103 20448 34115 20451
rect 34146 20448 34152 20460
rect 34103 20420 34152 20448
rect 34103 20417 34115 20420
rect 34057 20411 34115 20417
rect 34146 20408 34152 20420
rect 34204 20408 34210 20460
rect 34422 20408 34428 20460
rect 34480 20408 34486 20460
rect 34514 20408 34520 20460
rect 34572 20408 34578 20460
rect 34701 20451 34759 20457
rect 34701 20417 34713 20451
rect 34747 20417 34759 20451
rect 34701 20411 34759 20417
rect 27706 20340 27712 20392
rect 27764 20380 27770 20392
rect 28445 20383 28503 20389
rect 28445 20380 28457 20383
rect 27764 20352 28457 20380
rect 27764 20340 27770 20352
rect 28445 20349 28457 20352
rect 28491 20349 28503 20383
rect 28445 20343 28503 20349
rect 31481 20383 31539 20389
rect 31481 20349 31493 20383
rect 31527 20380 31539 20383
rect 31754 20380 31760 20392
rect 31527 20352 31760 20380
rect 31527 20349 31539 20352
rect 31481 20343 31539 20349
rect 31754 20340 31760 20352
rect 31812 20340 31818 20392
rect 33226 20340 33232 20392
rect 33284 20380 33290 20392
rect 34716 20380 34744 20411
rect 33284 20352 34744 20380
rect 33284 20340 33290 20352
rect 25777 20247 25835 20253
rect 25777 20244 25789 20247
rect 25096 20216 25789 20244
rect 25096 20204 25102 20216
rect 25777 20213 25789 20216
rect 25823 20213 25835 20247
rect 25777 20207 25835 20213
rect 26973 20247 27031 20253
rect 26973 20213 26985 20247
rect 27019 20244 27031 20247
rect 28442 20244 28448 20256
rect 27019 20216 28448 20244
rect 27019 20213 27031 20216
rect 26973 20207 27031 20213
rect 28442 20204 28448 20216
rect 28500 20204 28506 20256
rect 1104 20154 37076 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 37076 20154
rect 1104 20080 37076 20102
rect 1946 20000 1952 20052
rect 2004 20040 2010 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2004 20012 2973 20040
rect 2004 20000 2010 20012
rect 2961 20009 2973 20012
rect 3007 20040 3019 20043
rect 4062 20040 4068 20052
rect 3007 20012 4068 20040
rect 3007 20009 3019 20012
rect 2961 20003 3019 20009
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 7834 20000 7840 20052
rect 7892 20040 7898 20052
rect 7929 20043 7987 20049
rect 7929 20040 7941 20043
rect 7892 20012 7941 20040
rect 7892 20000 7898 20012
rect 7929 20009 7941 20012
rect 7975 20040 7987 20043
rect 8018 20040 8024 20052
rect 7975 20012 8024 20040
rect 7975 20009 7987 20012
rect 7929 20003 7987 20009
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 8110 20000 8116 20052
rect 8168 20000 8174 20052
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 11054 20040 11060 20052
rect 10183 20012 11060 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 18414 20000 18420 20052
rect 18472 20000 18478 20052
rect 24029 20043 24087 20049
rect 24029 20009 24041 20043
rect 24075 20040 24087 20043
rect 24854 20040 24860 20052
rect 24075 20012 24860 20040
rect 24075 20009 24087 20012
rect 24029 20003 24087 20009
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 26510 20000 26516 20052
rect 26568 20000 26574 20052
rect 26528 19972 26556 20000
rect 26528 19944 27292 19972
rect 9766 19864 9772 19916
rect 9824 19864 9830 19916
rect 19245 19907 19303 19913
rect 19245 19873 19257 19907
rect 19291 19904 19303 19907
rect 19518 19904 19524 19916
rect 19291 19876 19524 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 24765 19907 24823 19913
rect 24765 19873 24777 19907
rect 24811 19904 24823 19907
rect 25406 19904 25412 19916
rect 24811 19876 25412 19904
rect 24811 19873 24823 19876
rect 24765 19867 24823 19873
rect 25406 19864 25412 19876
rect 25464 19904 25470 19916
rect 26970 19904 26976 19916
rect 25464 19876 26976 19904
rect 25464 19864 25470 19876
rect 26970 19864 26976 19876
rect 27028 19864 27034 19916
rect 2406 19796 2412 19848
rect 2464 19796 2470 19848
rect 2590 19796 2596 19848
rect 2648 19796 2654 19848
rect 8202 19836 8208 19848
rect 7760 19808 8208 19836
rect 1762 19728 1768 19780
rect 1820 19768 1826 19780
rect 3142 19768 3148 19780
rect 1820 19740 3148 19768
rect 1820 19728 1826 19740
rect 3142 19728 3148 19740
rect 3200 19768 3206 19780
rect 3878 19768 3884 19780
rect 3200 19740 3884 19768
rect 3200 19728 3206 19740
rect 3878 19728 3884 19740
rect 3936 19728 3942 19780
rect 7760 19777 7788 19808
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9916 19808 9965 19836
rect 9916 19796 9922 19808
rect 9953 19805 9965 19808
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19805 16727 19839
rect 16669 19799 16727 19805
rect 7745 19771 7803 19777
rect 7745 19737 7757 19771
rect 7791 19737 7803 19771
rect 7745 19731 7803 19737
rect 7926 19728 7932 19780
rect 7984 19777 7990 19780
rect 7984 19771 8003 19777
rect 7991 19737 8003 19771
rect 16684 19768 16712 19799
rect 22278 19796 22284 19848
rect 22336 19796 22342 19848
rect 26142 19796 26148 19848
rect 26200 19796 26206 19848
rect 27062 19796 27068 19848
rect 27120 19796 27126 19848
rect 27264 19845 27292 19944
rect 27706 19864 27712 19916
rect 27764 19864 27770 19916
rect 28442 19864 28448 19916
rect 28500 19864 28506 19916
rect 30300 19876 31340 19904
rect 30300 19848 30328 19876
rect 27249 19839 27307 19845
rect 27249 19805 27261 19839
rect 27295 19805 27307 19839
rect 27249 19799 27307 19805
rect 27341 19839 27399 19845
rect 27341 19805 27353 19839
rect 27387 19805 27399 19839
rect 27341 19799 27399 19805
rect 28169 19839 28227 19845
rect 28169 19805 28181 19839
rect 28215 19805 28227 19839
rect 28169 19799 28227 19805
rect 16850 19768 16856 19780
rect 16684 19740 16856 19768
rect 7984 19731 8003 19737
rect 7984 19728 7990 19731
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 16945 19771 17003 19777
rect 16945 19737 16957 19771
rect 16991 19737 17003 19771
rect 19242 19768 19248 19780
rect 18170 19740 19248 19768
rect 16945 19731 17003 19737
rect 2314 19660 2320 19712
rect 2372 19700 2378 19712
rect 2501 19703 2559 19709
rect 2501 19700 2513 19703
rect 2372 19672 2513 19700
rect 2372 19660 2378 19672
rect 2501 19669 2513 19672
rect 2547 19669 2559 19703
rect 2501 19663 2559 19669
rect 2590 19660 2596 19712
rect 2648 19700 2654 19712
rect 2958 19709 2964 19712
rect 2777 19703 2835 19709
rect 2777 19700 2789 19703
rect 2648 19672 2789 19700
rect 2648 19660 2654 19672
rect 2777 19669 2789 19672
rect 2823 19669 2835 19703
rect 2777 19663 2835 19669
rect 2945 19703 2964 19709
rect 2945 19669 2957 19703
rect 3016 19700 3022 19712
rect 3970 19700 3976 19712
rect 3016 19672 3976 19700
rect 2945 19663 2964 19669
rect 2958 19660 2964 19663
rect 3016 19660 3022 19672
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 16960 19700 16988 19731
rect 19242 19728 19248 19740
rect 19300 19768 19306 19780
rect 19521 19771 19579 19777
rect 19300 19740 19472 19768
rect 19300 19728 19306 19740
rect 17770 19700 17776 19712
rect 16960 19672 17776 19700
rect 17770 19660 17776 19672
rect 17828 19660 17834 19712
rect 19444 19700 19472 19740
rect 19521 19737 19533 19771
rect 19567 19768 19579 19771
rect 19794 19768 19800 19780
rect 19567 19740 19800 19768
rect 19567 19737 19579 19740
rect 19521 19731 19579 19737
rect 19794 19728 19800 19740
rect 19852 19728 19858 19780
rect 19904 19740 20010 19768
rect 19904 19700 19932 19740
rect 22554 19728 22560 19780
rect 22612 19728 22618 19780
rect 23782 19740 24992 19768
rect 20898 19700 20904 19712
rect 19444 19672 20904 19700
rect 20898 19660 20904 19672
rect 20956 19660 20962 19712
rect 20990 19660 20996 19712
rect 21048 19660 21054 19712
rect 24964 19700 24992 19740
rect 25038 19728 25044 19780
rect 25096 19728 25102 19780
rect 26602 19728 26608 19780
rect 26660 19728 26666 19780
rect 25130 19700 25136 19712
rect 24964 19672 25136 19700
rect 25130 19660 25136 19672
rect 25188 19660 25194 19712
rect 26050 19660 26056 19712
rect 26108 19700 26114 19712
rect 27356 19700 27384 19799
rect 26108 19672 27384 19700
rect 28184 19700 28212 19799
rect 28350 19796 28356 19848
rect 28408 19796 28414 19848
rect 30009 19839 30067 19845
rect 30009 19805 30021 19839
rect 30055 19805 30067 19839
rect 30009 19799 30067 19805
rect 29086 19728 29092 19780
rect 29144 19768 29150 19780
rect 29549 19771 29607 19777
rect 29549 19768 29561 19771
rect 29144 19740 29561 19768
rect 29144 19728 29150 19740
rect 29549 19737 29561 19740
rect 29595 19737 29607 19771
rect 29549 19731 29607 19737
rect 30024 19700 30052 19799
rect 30190 19796 30196 19848
rect 30248 19796 30254 19848
rect 30282 19796 30288 19848
rect 30340 19796 30346 19848
rect 31110 19796 31116 19848
rect 31168 19796 31174 19848
rect 31312 19845 31340 19876
rect 34514 19864 34520 19916
rect 34572 19904 34578 19916
rect 35437 19907 35495 19913
rect 35437 19904 35449 19907
rect 34572 19876 35449 19904
rect 34572 19864 34578 19876
rect 35437 19873 35449 19876
rect 35483 19873 35495 19907
rect 35437 19867 35495 19873
rect 31297 19839 31355 19845
rect 31297 19805 31309 19839
rect 31343 19805 31355 19839
rect 31297 19799 31355 19805
rect 31386 19796 31392 19848
rect 31444 19796 31450 19848
rect 35161 19839 35219 19845
rect 35161 19836 35173 19839
rect 31726 19808 35173 19836
rect 30374 19728 30380 19780
rect 30432 19768 30438 19780
rect 30653 19771 30711 19777
rect 30653 19768 30665 19771
rect 30432 19740 30665 19768
rect 30432 19728 30438 19740
rect 30653 19737 30665 19740
rect 30699 19737 30711 19771
rect 30653 19731 30711 19737
rect 31128 19768 31156 19796
rect 31726 19768 31754 19808
rect 35161 19805 35173 19808
rect 35207 19805 35219 19839
rect 35161 19799 35219 19805
rect 35342 19796 35348 19848
rect 35400 19796 35406 19848
rect 31128 19740 31754 19768
rect 31128 19700 31156 19740
rect 34698 19728 34704 19780
rect 34756 19728 34762 19780
rect 28184 19672 31156 19700
rect 26108 19660 26114 19672
rect 1104 19610 37076 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 37076 19610
rect 1104 19536 37076 19558
rect 1850 19499 1908 19505
rect 1850 19465 1862 19499
rect 1896 19496 1908 19499
rect 2406 19496 2412 19508
rect 1896 19468 2412 19496
rect 1896 19465 1908 19468
rect 1850 19459 1908 19465
rect 2406 19456 2412 19468
rect 2464 19456 2470 19508
rect 2958 19496 2964 19508
rect 2516 19468 2964 19496
rect 1762 19388 1768 19440
rect 1820 19388 1826 19440
rect 1946 19388 1952 19440
rect 2004 19388 2010 19440
rect 2516 19428 2544 19468
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 8018 19456 8024 19508
rect 8076 19496 8082 19508
rect 8205 19499 8263 19505
rect 8205 19496 8217 19499
rect 8076 19468 8217 19496
rect 8076 19456 8082 19468
rect 8205 19465 8217 19468
rect 8251 19465 8263 19499
rect 8205 19459 8263 19465
rect 8312 19468 9352 19496
rect 2056 19400 2544 19428
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 2056 19360 2084 19400
rect 3050 19388 3056 19440
rect 3108 19388 3114 19440
rect 6822 19388 6828 19440
rect 6880 19428 6886 19440
rect 6914 19428 6920 19440
rect 6880 19400 6920 19428
rect 6880 19388 6886 19400
rect 6914 19388 6920 19400
rect 6972 19428 6978 19440
rect 8312 19428 8340 19468
rect 9324 19428 9352 19468
rect 16114 19456 16120 19508
rect 16172 19496 16178 19508
rect 18414 19496 18420 19508
rect 16172 19468 17448 19496
rect 16172 19456 16178 19468
rect 9398 19428 9404 19440
rect 6972 19400 8340 19428
rect 9246 19400 9404 19428
rect 6972 19388 6978 19400
rect 9398 19388 9404 19400
rect 9456 19388 9462 19440
rect 16022 19428 16028 19440
rect 15594 19400 16028 19428
rect 16022 19388 16028 19400
rect 16080 19388 16086 19440
rect 16574 19388 16580 19440
rect 16632 19428 16638 19440
rect 16669 19431 16727 19437
rect 16669 19428 16681 19431
rect 16632 19400 16681 19428
rect 16632 19388 16638 19400
rect 16669 19397 16681 19400
rect 16715 19397 16727 19431
rect 16669 19391 16727 19397
rect 1719 19332 2084 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 3970 19320 3976 19372
rect 4028 19360 4034 19372
rect 4157 19363 4215 19369
rect 4157 19360 4169 19363
rect 4028 19332 4169 19360
rect 4028 19320 4034 19332
rect 4157 19329 4169 19332
rect 4203 19329 4215 19363
rect 4157 19323 4215 19329
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 4614 19360 4620 19372
rect 4387 19332 4620 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 4614 19320 4620 19332
rect 4672 19320 4678 19372
rect 4798 19320 4804 19372
rect 4856 19320 4862 19372
rect 6181 19363 6239 19369
rect 6181 19329 6193 19363
rect 6227 19360 6239 19363
rect 6362 19360 6368 19372
rect 6227 19332 6368 19360
rect 6227 19329 6239 19332
rect 6181 19323 6239 19329
rect 6362 19320 6368 19332
rect 6420 19320 6426 19372
rect 9953 19363 10011 19369
rect 9953 19329 9965 19363
rect 9999 19360 10011 19363
rect 10042 19360 10048 19372
rect 9999 19332 10048 19360
rect 9999 19329 10011 19332
rect 9953 19323 10011 19329
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 14093 19363 14151 19369
rect 14093 19360 14105 19363
rect 13872 19332 14105 19360
rect 13872 19320 13878 19332
rect 14093 19329 14105 19332
rect 14139 19329 14151 19363
rect 14093 19323 14151 19329
rect 17126 19320 17132 19372
rect 17184 19320 17190 19372
rect 17420 19369 17448 19468
rect 18156 19468 18420 19496
rect 18046 19428 18052 19440
rect 17512 19400 18052 19428
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19329 17463 19363
rect 17405 19323 17463 19329
rect 1394 19252 1400 19304
rect 1452 19292 1458 19304
rect 2041 19295 2099 19301
rect 2041 19292 2053 19295
rect 1452 19264 2053 19292
rect 1452 19252 1458 19264
rect 2041 19261 2053 19264
rect 2087 19261 2099 19295
rect 2041 19255 2099 19261
rect 2314 19252 2320 19304
rect 2372 19252 2378 19304
rect 4249 19295 4307 19301
rect 4249 19261 4261 19295
rect 4295 19292 4307 19295
rect 5905 19295 5963 19301
rect 5905 19292 5917 19295
rect 4295 19264 5917 19292
rect 4295 19261 4307 19264
rect 4249 19255 4307 19261
rect 5905 19261 5917 19264
rect 5951 19261 5963 19295
rect 5905 19255 5963 19261
rect 9674 19252 9680 19304
rect 9732 19252 9738 19304
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19292 14427 19295
rect 15010 19292 15016 19304
rect 14415 19264 15016 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 17328 19292 17356 19323
rect 17512 19292 17540 19400
rect 18046 19388 18052 19400
rect 18104 19388 18110 19440
rect 18156 19437 18184 19468
rect 18414 19456 18420 19468
rect 18472 19456 18478 19508
rect 22554 19456 22560 19508
rect 22612 19496 22618 19508
rect 23293 19499 23351 19505
rect 23293 19496 23305 19499
rect 22612 19468 23305 19496
rect 22612 19456 22618 19468
rect 23293 19465 23305 19468
rect 23339 19465 23351 19499
rect 23293 19459 23351 19465
rect 23661 19499 23719 19505
rect 23661 19465 23673 19499
rect 23707 19496 23719 19499
rect 24854 19496 24860 19508
rect 23707 19468 24860 19496
rect 23707 19465 23719 19468
rect 23661 19459 23719 19465
rect 24854 19456 24860 19468
rect 24912 19456 24918 19508
rect 25130 19456 25136 19508
rect 25188 19496 25194 19508
rect 26142 19496 26148 19508
rect 25188 19468 26148 19496
rect 25188 19456 25194 19468
rect 26142 19456 26148 19468
rect 26200 19496 26206 19508
rect 27982 19496 27988 19508
rect 26200 19468 27988 19496
rect 26200 19456 26234 19468
rect 27982 19456 27988 19468
rect 28040 19456 28046 19508
rect 30466 19456 30472 19508
rect 30524 19496 30530 19508
rect 31205 19499 31263 19505
rect 31205 19496 31217 19499
rect 30524 19468 31217 19496
rect 30524 19456 30530 19468
rect 31205 19465 31217 19468
rect 31251 19465 31263 19499
rect 31205 19459 31263 19465
rect 34146 19456 34152 19508
rect 34204 19456 34210 19508
rect 34514 19456 34520 19508
rect 34572 19496 34578 19508
rect 35805 19499 35863 19505
rect 35805 19496 35817 19499
rect 34572 19468 35817 19496
rect 34572 19456 34578 19468
rect 35805 19465 35817 19468
rect 35851 19465 35863 19499
rect 35805 19459 35863 19465
rect 18141 19431 18199 19437
rect 18141 19397 18153 19431
rect 18187 19397 18199 19431
rect 18141 19391 18199 19397
rect 18322 19388 18328 19440
rect 18380 19388 18386 19440
rect 19794 19388 19800 19440
rect 19852 19428 19858 19440
rect 20165 19431 20223 19437
rect 20165 19428 20177 19431
rect 19852 19400 20177 19428
rect 19852 19388 19858 19400
rect 20165 19397 20177 19400
rect 20211 19397 20223 19431
rect 26206 19428 26234 19456
rect 26082 19400 26234 19428
rect 26513 19431 26571 19437
rect 20165 19391 20223 19397
rect 26513 19397 26525 19431
rect 26559 19428 26571 19431
rect 26602 19428 26608 19440
rect 26559 19400 26608 19428
rect 26559 19397 26571 19400
rect 26513 19391 26571 19397
rect 26602 19388 26608 19400
rect 26660 19388 26666 19440
rect 34164 19428 34192 19456
rect 34072 19400 34192 19428
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 20625 19363 20683 19369
rect 17828 19332 17908 19360
rect 17828 19320 17834 19332
rect 17328 19264 17540 19292
rect 17880 19233 17908 19332
rect 20625 19329 20637 19363
rect 20671 19360 20683 19363
rect 20714 19360 20720 19372
rect 20671 19332 20720 19360
rect 20671 19329 20683 19332
rect 20625 19323 20683 19329
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 20806 19320 20812 19372
rect 20864 19320 20870 19372
rect 20901 19363 20959 19369
rect 20901 19329 20913 19363
rect 20947 19360 20959 19363
rect 20990 19360 20996 19372
rect 20947 19332 20996 19360
rect 20947 19329 20959 19332
rect 20901 19323 20959 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 29270 19320 29276 19372
rect 29328 19360 29334 19372
rect 29641 19363 29699 19369
rect 29641 19360 29653 19363
rect 29328 19332 29653 19360
rect 29328 19320 29334 19332
rect 29641 19329 29653 19332
rect 29687 19360 29699 19363
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 29687 19332 29745 19360
rect 29687 19329 29699 19332
rect 29641 19323 29699 19329
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 30929 19363 30987 19369
rect 30929 19329 30941 19363
rect 30975 19360 30987 19363
rect 31110 19360 31116 19372
rect 30975 19332 31116 19360
rect 30975 19329 30987 19332
rect 30929 19323 30987 19329
rect 31110 19320 31116 19332
rect 31168 19320 31174 19372
rect 31573 19363 31631 19369
rect 31573 19329 31585 19363
rect 31619 19360 31631 19363
rect 31938 19360 31944 19372
rect 31619 19332 31944 19360
rect 31619 19329 31631 19332
rect 31573 19323 31631 19329
rect 31938 19320 31944 19332
rect 31996 19320 32002 19372
rect 34072 19369 34100 19400
rect 34057 19363 34115 19369
rect 34057 19329 34069 19363
rect 34103 19329 34115 19363
rect 34057 19323 34115 19329
rect 35434 19320 35440 19372
rect 35492 19320 35498 19372
rect 18417 19295 18475 19301
rect 18417 19261 18429 19295
rect 18463 19292 18475 19295
rect 18598 19292 18604 19304
rect 18463 19264 18604 19292
rect 18463 19261 18475 19264
rect 18417 19255 18475 19261
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 23750 19252 23756 19304
rect 23808 19252 23814 19304
rect 23845 19295 23903 19301
rect 23845 19261 23857 19295
rect 23891 19261 23903 19295
rect 23845 19255 23903 19261
rect 25041 19295 25099 19301
rect 25041 19261 25053 19295
rect 25087 19292 25099 19295
rect 26050 19292 26056 19304
rect 25087 19264 26056 19292
rect 25087 19261 25099 19264
rect 25041 19255 25099 19261
rect 17865 19227 17923 19233
rect 17865 19193 17877 19227
rect 17911 19193 17923 19227
rect 17865 19187 17923 19193
rect 23658 19184 23664 19236
rect 23716 19224 23722 19236
rect 23860 19224 23888 19255
rect 26050 19252 26056 19264
rect 26108 19252 26114 19304
rect 26789 19295 26847 19301
rect 26789 19261 26801 19295
rect 26835 19292 26847 19295
rect 26970 19292 26976 19304
rect 26835 19264 26976 19292
rect 26835 19261 26847 19264
rect 26789 19255 26847 19261
rect 26970 19252 26976 19264
rect 27028 19252 27034 19304
rect 31294 19252 31300 19304
rect 31352 19292 31358 19304
rect 31665 19295 31723 19301
rect 31665 19292 31677 19295
rect 31352 19264 31677 19292
rect 31352 19252 31358 19264
rect 31665 19261 31677 19264
rect 31711 19261 31723 19295
rect 31665 19255 31723 19261
rect 31754 19252 31760 19304
rect 31812 19292 31818 19304
rect 31849 19295 31907 19301
rect 31849 19292 31861 19295
rect 31812 19264 31861 19292
rect 31812 19252 31818 19264
rect 31849 19261 31861 19264
rect 31895 19292 31907 19295
rect 33134 19292 33140 19304
rect 31895 19264 33140 19292
rect 31895 19261 31907 19264
rect 31849 19255 31907 19261
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 34333 19295 34391 19301
rect 34333 19261 34345 19295
rect 34379 19292 34391 19295
rect 34698 19292 34704 19304
rect 34379 19264 34704 19292
rect 34379 19261 34391 19264
rect 34333 19255 34391 19261
rect 34698 19252 34704 19264
rect 34756 19252 34762 19304
rect 23716 19196 23888 19224
rect 23716 19184 23722 19196
rect 3789 19159 3847 19165
rect 3789 19125 3801 19159
rect 3835 19156 3847 19159
rect 4062 19156 4068 19168
rect 3835 19128 4068 19156
rect 3835 19125 3847 19128
rect 3789 19119 3847 19125
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 4433 19159 4491 19165
rect 4433 19125 4445 19159
rect 4479 19156 4491 19159
rect 4614 19156 4620 19168
rect 4479 19128 4620 19156
rect 4479 19125 4491 19128
rect 4433 19119 4491 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 15838 19116 15844 19168
rect 15896 19116 15902 19168
rect 27062 19116 27068 19168
rect 27120 19156 27126 19168
rect 28353 19159 28411 19165
rect 28353 19156 28365 19159
rect 27120 19128 28365 19156
rect 27120 19116 27126 19128
rect 28353 19125 28365 19128
rect 28399 19156 28411 19159
rect 29454 19156 29460 19168
rect 28399 19128 29460 19156
rect 28399 19125 28411 19128
rect 28353 19119 28411 19125
rect 29454 19116 29460 19128
rect 29512 19156 29518 19168
rect 33226 19156 33232 19168
rect 29512 19128 33232 19156
rect 29512 19116 29518 19128
rect 33226 19116 33232 19128
rect 33284 19116 33290 19168
rect 1104 19066 37076 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 37076 19066
rect 1104 18992 37076 19014
rect 8754 18912 8760 18964
rect 8812 18912 8818 18964
rect 18322 18912 18328 18964
rect 18380 18952 18386 18964
rect 18693 18955 18751 18961
rect 18693 18952 18705 18955
rect 18380 18924 18705 18952
rect 18380 18912 18386 18924
rect 18693 18921 18705 18924
rect 18739 18921 18751 18955
rect 27062 18952 27068 18964
rect 18693 18915 18751 18921
rect 24964 18924 27068 18952
rect 16298 18844 16304 18896
rect 16356 18884 16362 18896
rect 16356 18856 16712 18884
rect 16356 18844 16362 18856
rect 1394 18776 1400 18828
rect 1452 18776 1458 18828
rect 4062 18776 4068 18828
rect 4120 18776 4126 18828
rect 4522 18776 4528 18828
rect 4580 18816 4586 18828
rect 4617 18819 4675 18825
rect 4617 18816 4629 18819
rect 4580 18788 4629 18816
rect 4580 18776 4586 18788
rect 4617 18785 4629 18788
rect 4663 18785 4675 18819
rect 4617 18779 4675 18785
rect 5077 18819 5135 18825
rect 5077 18785 5089 18819
rect 5123 18816 5135 18819
rect 6641 18819 6699 18825
rect 6641 18816 6653 18819
rect 5123 18788 6653 18816
rect 5123 18785 5135 18788
rect 5077 18779 5135 18785
rect 6641 18785 6653 18788
rect 6687 18785 6699 18819
rect 6641 18779 6699 18785
rect 7285 18819 7343 18825
rect 7285 18785 7297 18819
rect 7331 18816 7343 18819
rect 7742 18816 7748 18828
rect 7331 18788 7748 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 15010 18776 15016 18828
rect 15068 18776 15074 18828
rect 15749 18819 15807 18825
rect 15749 18785 15761 18819
rect 15795 18816 15807 18819
rect 15838 18816 15844 18828
rect 15795 18788 15844 18816
rect 15795 18785 15807 18788
rect 15749 18779 15807 18785
rect 15838 18776 15844 18788
rect 15896 18816 15902 18828
rect 16684 18825 16712 18856
rect 20898 18844 20904 18896
rect 20956 18884 20962 18896
rect 21453 18887 21511 18893
rect 21453 18884 21465 18887
rect 20956 18856 21465 18884
rect 20956 18844 20962 18856
rect 21453 18853 21465 18856
rect 21499 18853 21511 18887
rect 21453 18847 21511 18853
rect 16577 18819 16635 18825
rect 16577 18816 16589 18819
rect 15896 18788 16589 18816
rect 15896 18776 15902 18788
rect 16577 18785 16589 18788
rect 16623 18785 16635 18819
rect 16577 18779 16635 18785
rect 16669 18819 16727 18825
rect 16669 18785 16681 18819
rect 16715 18785 16727 18819
rect 16669 18779 16727 18785
rect 19518 18776 19524 18828
rect 19576 18776 19582 18828
rect 21913 18819 21971 18825
rect 21913 18785 21925 18819
rect 21959 18816 21971 18819
rect 22370 18816 22376 18828
rect 21959 18788 22376 18816
rect 21959 18785 21971 18788
rect 21913 18779 21971 18785
rect 22370 18776 22376 18788
rect 22428 18776 22434 18828
rect 3789 18751 3847 18757
rect 3789 18748 3801 18751
rect 3160 18720 3801 18748
rect 1670 18640 1676 18692
rect 1728 18640 1734 18692
rect 3050 18680 3056 18692
rect 2898 18652 3056 18680
rect 3050 18640 3056 18652
rect 3108 18640 3114 18692
rect 3160 18624 3188 18720
rect 3789 18717 3801 18720
rect 3835 18717 3847 18751
rect 3789 18711 3847 18717
rect 3878 18708 3884 18760
rect 3936 18748 3942 18760
rect 4157 18751 4215 18757
rect 4157 18748 4169 18751
rect 3936 18720 4169 18748
rect 3936 18708 3942 18720
rect 4157 18717 4169 18720
rect 4203 18717 4215 18751
rect 4157 18711 4215 18717
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 6917 18751 6975 18757
rect 4755 18720 5212 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4246 18640 4252 18692
rect 4304 18689 4310 18692
rect 4304 18683 4332 18689
rect 4320 18680 4332 18683
rect 4614 18680 4620 18692
rect 4320 18652 4620 18680
rect 4320 18649 4332 18652
rect 4304 18643 4332 18649
rect 4304 18640 4310 18643
rect 4614 18640 4620 18652
rect 4672 18640 4678 18692
rect 3142 18572 3148 18624
rect 3200 18572 3206 18624
rect 4433 18615 4491 18621
rect 4433 18581 4445 18615
rect 4479 18612 4491 18615
rect 4798 18612 4804 18624
rect 4479 18584 4804 18612
rect 4479 18581 4491 18584
rect 4433 18575 4491 18581
rect 4798 18572 4804 18584
rect 4856 18572 4862 18624
rect 5184 18621 5212 18720
rect 6917 18717 6929 18751
rect 6963 18748 6975 18751
rect 7009 18751 7067 18757
rect 7009 18748 7021 18751
rect 6963 18720 7021 18748
rect 6963 18717 6975 18720
rect 6917 18711 6975 18717
rect 7009 18717 7021 18720
rect 7055 18717 7067 18751
rect 7009 18711 7067 18717
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 6730 18680 6736 18692
rect 6210 18652 6736 18680
rect 5169 18615 5227 18621
rect 5169 18581 5181 18615
rect 5215 18612 5227 18615
rect 5258 18612 5264 18624
rect 5215 18584 5264 18612
rect 5215 18581 5227 18584
rect 5169 18575 5227 18581
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 5626 18572 5632 18624
rect 5684 18612 5690 18624
rect 6288 18612 6316 18652
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 5684 18584 6316 18612
rect 5684 18572 5690 18584
rect 6822 18572 6828 18624
rect 6880 18612 6886 18624
rect 6914 18612 6920 18624
rect 6880 18584 6920 18612
rect 6880 18572 6886 18584
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7024 18612 7052 18711
rect 9398 18680 9404 18692
rect 8510 18652 9404 18680
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 15488 18680 15516 18711
rect 15562 18708 15568 18760
rect 15620 18748 15626 18760
rect 15657 18751 15715 18757
rect 15657 18748 15669 18751
rect 15620 18720 15669 18748
rect 15620 18708 15626 18720
rect 15657 18717 15669 18720
rect 15703 18717 15715 18751
rect 15657 18711 15715 18717
rect 16850 18708 16856 18760
rect 16908 18748 16914 18760
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16908 18720 16957 18748
rect 16908 18708 16914 18720
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 24118 18708 24124 18760
rect 24176 18748 24182 18760
rect 24673 18751 24731 18757
rect 24673 18748 24685 18751
rect 24176 18720 24685 18748
rect 24176 18708 24182 18720
rect 24673 18717 24685 18720
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 24762 18708 24768 18760
rect 24820 18757 24826 18760
rect 24964 18757 24992 18924
rect 27062 18912 27068 18924
rect 27120 18912 27126 18964
rect 29273 18955 29331 18961
rect 29273 18921 29285 18955
rect 29319 18952 29331 18955
rect 30282 18952 30288 18964
rect 29319 18924 30288 18952
rect 29319 18921 29331 18924
rect 29273 18915 29331 18921
rect 30282 18912 30288 18924
rect 30340 18912 30346 18964
rect 31294 18912 31300 18964
rect 31352 18912 31358 18964
rect 35342 18844 35348 18896
rect 35400 18844 35406 18896
rect 29549 18819 29607 18825
rect 29549 18816 29561 18819
rect 27540 18788 29561 18816
rect 24820 18751 24849 18757
rect 24837 18717 24849 18751
rect 24820 18711 24849 18717
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 24820 18708 24826 18711
rect 26142 18708 26148 18760
rect 26200 18708 26206 18760
rect 26234 18708 26240 18760
rect 26292 18708 26298 18760
rect 26970 18708 26976 18760
rect 27028 18748 27034 18760
rect 27540 18757 27568 18788
rect 29549 18785 29561 18788
rect 29595 18785 29607 18819
rect 29549 18779 29607 18785
rect 29825 18819 29883 18825
rect 29825 18785 29837 18819
rect 29871 18816 29883 18819
rect 30374 18816 30380 18828
rect 29871 18788 30380 18816
rect 29871 18785 29883 18788
rect 29825 18779 29883 18785
rect 30374 18776 30380 18788
rect 30432 18776 30438 18828
rect 31846 18776 31852 18828
rect 31904 18816 31910 18828
rect 32033 18819 32091 18825
rect 32033 18816 32045 18819
rect 31904 18788 32045 18816
rect 31904 18776 31910 18788
rect 32033 18785 32045 18788
rect 32079 18785 32091 18819
rect 32033 18779 32091 18785
rect 32309 18819 32367 18825
rect 32309 18785 32321 18819
rect 32355 18816 32367 18819
rect 33318 18816 33324 18828
rect 32355 18788 33324 18816
rect 32355 18785 32367 18788
rect 32309 18779 32367 18785
rect 33318 18776 33324 18788
rect 33376 18776 33382 18828
rect 27525 18751 27583 18757
rect 27525 18748 27537 18751
rect 27028 18720 27537 18748
rect 27028 18708 27034 18720
rect 27525 18717 27537 18720
rect 27571 18717 27583 18751
rect 27525 18711 27583 18717
rect 35069 18751 35127 18757
rect 35069 18717 35081 18751
rect 35115 18748 35127 18751
rect 35250 18748 35256 18760
rect 35115 18720 35256 18748
rect 35115 18717 35127 18720
rect 35069 18711 35127 18717
rect 35250 18708 35256 18720
rect 35308 18708 35314 18760
rect 16206 18680 16212 18692
rect 15488 18652 16212 18680
rect 16206 18640 16212 18652
rect 16264 18640 16270 18692
rect 17218 18640 17224 18692
rect 17276 18640 17282 18692
rect 17954 18640 17960 18692
rect 18012 18640 18018 18692
rect 19794 18640 19800 18692
rect 19852 18640 19858 18692
rect 20806 18640 20812 18692
rect 20864 18640 20870 18692
rect 22005 18683 22063 18689
rect 22005 18680 22017 18683
rect 21100 18652 22017 18680
rect 7926 18612 7932 18624
rect 7024 18584 7932 18612
rect 7926 18572 7932 18584
rect 7984 18572 7990 18624
rect 14918 18572 14924 18624
rect 14976 18612 14982 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 14976 18584 16129 18612
rect 14976 18572 14982 18584
rect 16117 18581 16129 18584
rect 16163 18581 16175 18615
rect 16117 18575 16175 18581
rect 16482 18572 16488 18624
rect 16540 18572 16546 18624
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 21100 18612 21128 18652
rect 22005 18649 22017 18652
rect 22051 18649 22063 18683
rect 22005 18643 22063 18649
rect 25409 18683 25467 18689
rect 25409 18649 25421 18683
rect 25455 18649 25467 18683
rect 25409 18643 25467 18649
rect 25501 18683 25559 18689
rect 25501 18649 25513 18683
rect 25547 18680 25559 18683
rect 26007 18683 26065 18689
rect 25547 18652 25912 18680
rect 25547 18649 25559 18652
rect 25501 18643 25559 18649
rect 20772 18584 21128 18612
rect 20772 18572 20778 18584
rect 21266 18572 21272 18624
rect 21324 18612 21330 18624
rect 21913 18615 21971 18621
rect 21913 18612 21925 18615
rect 21324 18584 21925 18612
rect 21324 18572 21330 18584
rect 21913 18581 21925 18584
rect 21959 18581 21971 18615
rect 25424 18612 25452 18643
rect 25590 18612 25596 18624
rect 25424 18584 25596 18612
rect 21913 18575 21971 18581
rect 25590 18572 25596 18584
rect 25648 18572 25654 18624
rect 25884 18612 25912 18652
rect 26007 18649 26019 18683
rect 26053 18680 26065 18683
rect 27062 18680 27068 18692
rect 26053 18652 27068 18680
rect 26053 18649 26065 18652
rect 26007 18643 26065 18649
rect 27062 18640 27068 18652
rect 27120 18640 27126 18692
rect 27801 18683 27859 18689
rect 27801 18649 27813 18683
rect 27847 18649 27859 18683
rect 27801 18643 27859 18649
rect 26326 18612 26332 18624
rect 25884 18584 26332 18612
rect 26326 18572 26332 18584
rect 26384 18572 26390 18624
rect 27816 18612 27844 18643
rect 28258 18640 28264 18692
rect 28316 18640 28322 18692
rect 30834 18640 30840 18692
rect 30892 18640 30898 18692
rect 33594 18680 33600 18692
rect 33534 18652 33600 18680
rect 33594 18640 33600 18652
rect 33652 18640 33658 18692
rect 34790 18640 34796 18692
rect 34848 18640 34854 18692
rect 29086 18612 29092 18624
rect 27816 18584 29092 18612
rect 29086 18572 29092 18584
rect 29144 18572 29150 18624
rect 33778 18572 33784 18624
rect 33836 18612 33842 18624
rect 34885 18615 34943 18621
rect 34885 18612 34897 18615
rect 33836 18584 34897 18612
rect 33836 18572 33842 18584
rect 34885 18581 34897 18584
rect 34931 18581 34943 18615
rect 34885 18575 34943 18581
rect 1104 18522 37076 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 37076 18522
rect 1104 18448 37076 18470
rect 3970 18368 3976 18420
rect 4028 18368 4034 18420
rect 4141 18411 4199 18417
rect 4141 18377 4153 18411
rect 4187 18408 4199 18411
rect 4522 18408 4528 18420
rect 4187 18380 4528 18408
rect 4187 18377 4199 18380
rect 4141 18371 4199 18377
rect 4522 18368 4528 18380
rect 4580 18408 4586 18420
rect 4890 18408 4896 18420
rect 4580 18380 4896 18408
rect 4580 18368 4586 18380
rect 4890 18368 4896 18380
rect 4948 18368 4954 18420
rect 10042 18368 10048 18420
rect 10100 18368 10106 18420
rect 16393 18411 16451 18417
rect 16393 18377 16405 18411
rect 16439 18408 16451 18411
rect 16482 18408 16488 18420
rect 16439 18380 16488 18408
rect 16439 18377 16451 18380
rect 16393 18371 16451 18377
rect 16482 18368 16488 18380
rect 16540 18368 16546 18420
rect 17218 18368 17224 18420
rect 17276 18408 17282 18420
rect 18031 18411 18089 18417
rect 18031 18408 18043 18411
rect 17276 18380 18043 18408
rect 17276 18368 17282 18380
rect 18031 18377 18043 18380
rect 18077 18377 18089 18411
rect 28721 18411 28779 18417
rect 18031 18371 18089 18377
rect 22296 18380 25912 18408
rect 4341 18343 4399 18349
rect 4341 18309 4353 18343
rect 4387 18340 4399 18343
rect 5258 18340 5264 18352
rect 4387 18312 5264 18340
rect 4387 18309 4399 18312
rect 4341 18303 4399 18309
rect 5258 18300 5264 18312
rect 5316 18300 5322 18352
rect 6181 18343 6239 18349
rect 6181 18309 6193 18343
rect 6227 18340 6239 18343
rect 7650 18340 7656 18352
rect 6227 18312 7656 18340
rect 6227 18309 6239 18312
rect 6181 18303 6239 18309
rect 7650 18300 7656 18312
rect 7708 18340 7714 18352
rect 7745 18343 7803 18349
rect 7745 18340 7757 18343
rect 7708 18312 7757 18340
rect 7708 18300 7714 18312
rect 7745 18309 7757 18312
rect 7791 18309 7803 18343
rect 7745 18303 7803 18309
rect 7926 18300 7932 18352
rect 7984 18340 7990 18352
rect 9493 18343 9551 18349
rect 9493 18340 9505 18343
rect 7984 18312 9505 18340
rect 7984 18300 7990 18312
rect 9493 18309 9505 18312
rect 9539 18340 9551 18343
rect 10060 18340 10088 18368
rect 9539 18312 10088 18340
rect 9539 18309 9551 18312
rect 9493 18303 9551 18309
rect 1578 18232 1584 18284
rect 1636 18232 1642 18284
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18272 2283 18275
rect 3142 18272 3148 18284
rect 2271 18244 3148 18272
rect 2271 18241 2283 18244
rect 2225 18235 2283 18241
rect 3142 18232 3148 18244
rect 3200 18232 3206 18284
rect 9600 18281 9628 18312
rect 14918 18300 14924 18352
rect 14976 18300 14982 18352
rect 15654 18300 15660 18352
rect 15712 18300 15718 18352
rect 18322 18300 18328 18352
rect 18380 18300 18386 18352
rect 18509 18343 18567 18349
rect 18509 18309 18521 18343
rect 18555 18340 18567 18343
rect 19058 18340 19064 18352
rect 18555 18312 19064 18340
rect 18555 18309 18567 18312
rect 18509 18303 18567 18309
rect 19058 18300 19064 18312
rect 19116 18300 19122 18352
rect 19794 18300 19800 18352
rect 19852 18340 19858 18352
rect 20257 18343 20315 18349
rect 20257 18340 20269 18343
rect 19852 18312 20269 18340
rect 19852 18300 19858 18312
rect 20257 18309 20269 18312
rect 20303 18309 20315 18343
rect 20990 18340 20996 18352
rect 20257 18303 20315 18309
rect 20916 18312 20996 18340
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 1670 18164 1676 18216
rect 1728 18204 1734 18216
rect 1857 18207 1915 18213
rect 1857 18204 1869 18207
rect 1728 18176 1869 18204
rect 1728 18164 1734 18176
rect 1857 18173 1869 18176
rect 1903 18173 1915 18207
rect 1857 18167 1915 18173
rect 2317 18207 2375 18213
rect 2317 18173 2329 18207
rect 2363 18204 2375 18207
rect 2590 18204 2596 18216
rect 2363 18176 2596 18204
rect 2363 18173 2375 18176
rect 2317 18167 2375 18173
rect 2590 18164 2596 18176
rect 2648 18164 2654 18216
rect 9858 18164 9864 18216
rect 9916 18164 9922 18216
rect 4246 18136 4252 18148
rect 4172 18108 4252 18136
rect 1394 18028 1400 18080
rect 1452 18028 1458 18080
rect 4172 18077 4200 18108
rect 4246 18096 4252 18108
rect 4304 18136 4310 18148
rect 5074 18136 5080 18148
rect 4304 18108 5080 18136
rect 4304 18096 4310 18108
rect 5074 18096 5080 18108
rect 5132 18096 5138 18148
rect 4157 18071 4215 18077
rect 4157 18037 4169 18071
rect 4203 18037 4215 18071
rect 4157 18031 4215 18037
rect 4614 18028 4620 18080
rect 4672 18068 4678 18080
rect 4709 18071 4767 18077
rect 4709 18068 4721 18071
rect 4672 18040 4721 18068
rect 4672 18028 4678 18040
rect 4709 18037 4721 18040
rect 4755 18037 4767 18071
rect 4709 18031 4767 18037
rect 9398 18028 9404 18080
rect 9456 18068 9462 18080
rect 10980 18068 11008 18258
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14274 18272 14280 18284
rect 13872 18244 14280 18272
rect 13872 18232 13878 18244
rect 14274 18232 14280 18244
rect 14332 18272 14338 18284
rect 20916 18281 20944 18312
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 22296 18284 22324 18380
rect 23782 18326 24426 18340
rect 23782 18312 24440 18326
rect 14645 18275 14703 18281
rect 14645 18272 14657 18275
rect 14332 18244 14657 18272
rect 14332 18232 14338 18244
rect 14645 18241 14657 18244
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18241 20775 18275
rect 20717 18235 20775 18241
rect 20901 18275 20959 18281
rect 20901 18241 20913 18275
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 18598 18164 18604 18216
rect 18656 18164 18662 18216
rect 20732 18136 20760 18235
rect 22278 18232 22284 18284
rect 22336 18232 22342 18284
rect 20993 18207 21051 18213
rect 20993 18173 21005 18207
rect 21039 18204 21051 18207
rect 21266 18204 21272 18216
rect 21039 18176 21272 18204
rect 21039 18173 21051 18176
rect 20993 18167 21051 18173
rect 21266 18164 21272 18176
rect 21324 18164 21330 18216
rect 22554 18164 22560 18216
rect 22612 18164 22618 18216
rect 23750 18164 23756 18216
rect 23808 18204 23814 18216
rect 24029 18207 24087 18213
rect 24029 18204 24041 18207
rect 23808 18176 24041 18204
rect 23808 18164 23814 18176
rect 24029 18173 24041 18176
rect 24075 18173 24087 18207
rect 24029 18167 24087 18173
rect 24118 18164 24124 18216
rect 24176 18164 24182 18216
rect 24412 18204 24440 18312
rect 25590 18300 25596 18352
rect 25648 18300 25654 18352
rect 25884 18281 25912 18380
rect 28721 18377 28733 18411
rect 28767 18408 28779 18411
rect 28994 18408 29000 18420
rect 28767 18380 29000 18408
rect 28767 18377 28779 18380
rect 28721 18371 28779 18377
rect 28994 18368 29000 18380
rect 29052 18408 29058 18420
rect 30190 18408 30196 18420
rect 29052 18380 30196 18408
rect 29052 18368 29058 18380
rect 30190 18368 30196 18380
rect 30248 18368 30254 18420
rect 35342 18408 35348 18420
rect 32876 18380 35348 18408
rect 28258 18300 28264 18352
rect 28316 18300 28322 18352
rect 31938 18340 31944 18352
rect 31312 18312 31944 18340
rect 25869 18275 25927 18281
rect 25869 18241 25881 18275
rect 25915 18241 25927 18275
rect 25869 18235 25927 18241
rect 30561 18275 30619 18281
rect 30561 18241 30573 18275
rect 30607 18272 30619 18275
rect 30926 18272 30932 18284
rect 30607 18244 30932 18272
rect 30607 18241 30619 18244
rect 30561 18235 30619 18241
rect 30926 18232 30932 18244
rect 30984 18232 30990 18284
rect 31312 18281 31340 18312
rect 31938 18300 31944 18312
rect 31996 18300 32002 18352
rect 32876 18349 32904 18380
rect 35342 18368 35348 18380
rect 35400 18368 35406 18420
rect 32861 18343 32919 18349
rect 32861 18309 32873 18343
rect 32907 18309 32919 18343
rect 32861 18303 32919 18309
rect 33594 18300 33600 18352
rect 33652 18300 33658 18352
rect 31297 18275 31355 18281
rect 31297 18241 31309 18275
rect 31343 18241 31355 18275
rect 31297 18235 31355 18241
rect 31481 18275 31539 18281
rect 31481 18241 31493 18275
rect 31527 18272 31539 18275
rect 31527 18244 31616 18272
rect 31527 18241 31539 18244
rect 31481 18235 31539 18241
rect 25130 18204 25136 18216
rect 24412 18176 25136 18204
rect 25130 18164 25136 18176
rect 25188 18164 25194 18216
rect 26970 18164 26976 18216
rect 27028 18164 27034 18216
rect 27249 18207 27307 18213
rect 27249 18173 27261 18207
rect 27295 18204 27307 18207
rect 27614 18204 27620 18216
rect 27295 18176 27620 18204
rect 27295 18173 27307 18176
rect 27249 18167 27307 18173
rect 27614 18164 27620 18176
rect 27672 18164 27678 18216
rect 31202 18164 31208 18216
rect 31260 18164 31266 18216
rect 31588 18148 31616 18244
rect 31754 18164 31760 18216
rect 31812 18204 31818 18216
rect 31941 18207 31999 18213
rect 31941 18204 31953 18207
rect 31812 18176 31953 18204
rect 31812 18164 31818 18176
rect 31941 18173 31953 18176
rect 31987 18173 31999 18207
rect 31941 18167 31999 18173
rect 32122 18164 32128 18216
rect 32180 18204 32186 18216
rect 32585 18207 32643 18213
rect 32585 18204 32597 18207
rect 32180 18176 32597 18204
rect 32180 18164 32186 18176
rect 32585 18173 32597 18176
rect 32631 18173 32643 18207
rect 33410 18204 33416 18216
rect 32585 18167 32643 18173
rect 32692 18176 33416 18204
rect 22002 18136 22008 18148
rect 20732 18108 22008 18136
rect 22002 18096 22008 18108
rect 22060 18096 22066 18148
rect 31570 18096 31576 18148
rect 31628 18136 31634 18148
rect 32692 18136 32720 18176
rect 33410 18164 33416 18176
rect 33468 18164 33474 18216
rect 34333 18207 34391 18213
rect 34333 18173 34345 18207
rect 34379 18204 34391 18207
rect 35250 18204 35256 18216
rect 34379 18176 35256 18204
rect 34379 18173 34391 18176
rect 34333 18167 34391 18173
rect 35250 18164 35256 18176
rect 35308 18164 35314 18216
rect 31628 18108 32720 18136
rect 31628 18096 31634 18108
rect 9456 18040 11008 18068
rect 9456 18028 9462 18040
rect 11330 18028 11336 18080
rect 11388 18028 11394 18080
rect 23658 18028 23664 18080
rect 23716 18068 23722 18080
rect 27890 18068 27896 18080
rect 23716 18040 27896 18068
rect 23716 18028 23722 18040
rect 27890 18028 27896 18040
rect 27948 18068 27954 18080
rect 28718 18068 28724 18080
rect 27948 18040 28724 18068
rect 27948 18028 27954 18040
rect 28718 18028 28724 18040
rect 28776 18068 28782 18080
rect 29089 18071 29147 18077
rect 29089 18068 29101 18071
rect 28776 18040 29101 18068
rect 28776 18028 28782 18040
rect 29089 18037 29101 18040
rect 29135 18037 29147 18071
rect 29089 18031 29147 18037
rect 1104 17978 37076 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 37076 17978
rect 1104 17904 37076 17926
rect 1578 17824 1584 17876
rect 1636 17864 1642 17876
rect 1857 17867 1915 17873
rect 1857 17864 1869 17867
rect 1636 17836 1869 17864
rect 1636 17824 1642 17836
rect 1857 17833 1869 17836
rect 1903 17833 1915 17867
rect 1857 17827 1915 17833
rect 4706 17824 4712 17876
rect 4764 17864 4770 17876
rect 5077 17867 5135 17873
rect 5077 17864 5089 17867
rect 4764 17836 5089 17864
rect 4764 17824 4770 17836
rect 5077 17833 5089 17836
rect 5123 17833 5135 17867
rect 5077 17827 5135 17833
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 10229 17867 10287 17873
rect 10229 17864 10241 17867
rect 9916 17836 10241 17864
rect 9916 17824 9922 17836
rect 10229 17833 10241 17836
rect 10275 17833 10287 17867
rect 10229 17827 10287 17833
rect 10689 17867 10747 17873
rect 10689 17833 10701 17867
rect 10735 17864 10747 17867
rect 11330 17864 11336 17876
rect 10735 17836 11336 17864
rect 10735 17833 10747 17836
rect 10689 17827 10747 17833
rect 11330 17824 11336 17836
rect 11388 17824 11394 17876
rect 19058 17824 19064 17876
rect 19116 17824 19122 17876
rect 22370 17824 22376 17876
rect 22428 17824 22434 17876
rect 22554 17824 22560 17876
rect 22612 17864 22618 17876
rect 23385 17867 23443 17873
rect 23385 17864 23397 17867
rect 22612 17836 23397 17864
rect 22612 17824 22618 17836
rect 23385 17833 23397 17836
rect 23431 17833 23443 17867
rect 23385 17827 23443 17833
rect 24762 17824 24768 17876
rect 24820 17864 24826 17876
rect 26234 17864 26240 17876
rect 24820 17836 26240 17864
rect 24820 17824 24826 17836
rect 26234 17824 26240 17836
rect 26292 17824 26298 17876
rect 27614 17824 27620 17876
rect 27672 17864 27678 17876
rect 28353 17867 28411 17873
rect 28353 17864 28365 17867
rect 27672 17836 28365 17864
rect 27672 17824 27678 17836
rect 28353 17833 28365 17836
rect 28399 17833 28411 17867
rect 28353 17827 28411 17833
rect 31849 17867 31907 17873
rect 31849 17833 31861 17867
rect 31895 17864 31907 17867
rect 31938 17864 31944 17876
rect 31895 17836 31944 17864
rect 31895 17833 31907 17836
rect 31849 17827 31907 17833
rect 31938 17824 31944 17836
rect 31996 17824 32002 17876
rect 33318 17824 33324 17876
rect 33376 17824 33382 17876
rect 4249 17799 4307 17805
rect 4249 17765 4261 17799
rect 4295 17765 4307 17799
rect 4249 17759 4307 17765
rect 11241 17799 11299 17805
rect 11241 17765 11253 17799
rect 11287 17765 11299 17799
rect 11241 17759 11299 17765
rect 1486 17620 1492 17672
rect 1544 17660 1550 17672
rect 2041 17663 2099 17669
rect 2041 17660 2053 17663
rect 1544 17632 2053 17660
rect 1544 17620 1550 17632
rect 2041 17629 2053 17632
rect 2087 17629 2099 17663
rect 2041 17623 2099 17629
rect 3878 17620 3884 17672
rect 3936 17660 3942 17672
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3936 17632 3985 17660
rect 3936 17620 3942 17632
rect 3973 17629 3985 17632
rect 4019 17629 4031 17663
rect 4264 17660 4292 17759
rect 4890 17728 4896 17740
rect 4540 17700 4896 17728
rect 4540 17672 4568 17700
rect 4890 17688 4896 17700
rect 4948 17728 4954 17740
rect 6273 17731 6331 17737
rect 4948 17700 5396 17728
rect 4948 17688 4954 17700
rect 4341 17663 4399 17669
rect 4341 17660 4353 17663
rect 4264 17632 4353 17660
rect 3973 17623 4031 17629
rect 4341 17629 4353 17632
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 4522 17620 4528 17672
rect 4580 17620 4586 17672
rect 4614 17620 4620 17672
rect 4672 17620 4678 17672
rect 5074 17620 5080 17672
rect 5132 17620 5138 17672
rect 5368 17669 5396 17700
rect 6273 17697 6285 17731
rect 6319 17728 6331 17731
rect 6914 17728 6920 17740
rect 6319 17700 6920 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 6914 17688 6920 17700
rect 6972 17688 6978 17740
rect 11256 17728 11284 17759
rect 10244 17700 11284 17728
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 9858 17620 9864 17672
rect 9916 17660 9922 17672
rect 10244 17669 10272 17700
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 16850 17728 16856 17740
rect 14332 17700 16856 17728
rect 14332 17688 14338 17700
rect 16850 17688 16856 17700
rect 16908 17728 16914 17740
rect 17313 17731 17371 17737
rect 17313 17728 17325 17731
rect 16908 17700 17325 17728
rect 16908 17688 16914 17700
rect 17313 17697 17325 17700
rect 17359 17697 17371 17731
rect 17313 17691 17371 17697
rect 20625 17731 20683 17737
rect 20625 17697 20637 17731
rect 20671 17728 20683 17731
rect 22278 17728 22284 17740
rect 20671 17700 22284 17728
rect 20671 17697 20683 17700
rect 20625 17691 20683 17697
rect 22278 17688 22284 17700
rect 22336 17688 22342 17740
rect 23658 17688 23664 17740
rect 23716 17728 23722 17740
rect 23937 17731 23995 17737
rect 23937 17728 23949 17731
rect 23716 17700 23949 17728
rect 23716 17688 23722 17700
rect 23937 17697 23949 17700
rect 23983 17697 23995 17731
rect 23937 17691 23995 17697
rect 26234 17688 26240 17740
rect 26292 17728 26298 17740
rect 26513 17731 26571 17737
rect 26513 17728 26525 17731
rect 26292 17700 26525 17728
rect 26292 17688 26298 17700
rect 26513 17697 26525 17700
rect 26559 17697 26571 17731
rect 26513 17691 26571 17697
rect 28813 17731 28871 17737
rect 28813 17697 28825 17731
rect 28859 17728 28871 17731
rect 28994 17728 29000 17740
rect 28859 17700 29000 17728
rect 28859 17697 28871 17700
rect 28813 17691 28871 17697
rect 10045 17663 10103 17669
rect 10045 17660 10057 17663
rect 9916 17632 10057 17660
rect 9916 17620 9922 17632
rect 10045 17629 10057 17632
rect 10091 17629 10103 17663
rect 10045 17623 10103 17629
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 4249 17595 4307 17601
rect 4249 17561 4261 17595
rect 4295 17592 4307 17595
rect 4706 17592 4712 17604
rect 4295 17564 4712 17592
rect 4295 17561 4307 17564
rect 4249 17555 4307 17561
rect 4706 17552 4712 17564
rect 4764 17552 4770 17604
rect 6546 17552 6552 17604
rect 6604 17552 6610 17604
rect 6822 17552 6828 17604
rect 6880 17592 6886 17604
rect 6880 17564 7038 17592
rect 6880 17552 6886 17564
rect 3418 17484 3424 17536
rect 3476 17524 3482 17536
rect 4065 17527 4123 17533
rect 4065 17524 4077 17527
rect 3476 17496 4077 17524
rect 3476 17484 3482 17496
rect 4065 17493 4077 17496
rect 4111 17493 4123 17527
rect 4065 17487 4123 17493
rect 4338 17484 4344 17536
rect 4396 17524 4402 17536
rect 4433 17527 4491 17533
rect 4433 17524 4445 17527
rect 4396 17496 4445 17524
rect 4396 17484 4402 17496
rect 4433 17493 4445 17496
rect 4479 17493 4491 17527
rect 4433 17487 4491 17493
rect 5258 17484 5264 17536
rect 5316 17484 5322 17536
rect 7466 17484 7472 17536
rect 7524 17524 7530 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7524 17496 8033 17524
rect 7524 17484 7530 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 10060 17524 10088 17623
rect 10502 17620 10508 17672
rect 10560 17660 10566 17672
rect 10965 17663 11023 17669
rect 10965 17660 10977 17663
rect 10560 17632 10977 17660
rect 10560 17620 10566 17632
rect 10704 17601 10732 17632
rect 10965 17629 10977 17632
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17660 11299 17663
rect 11330 17660 11336 17672
rect 11287 17632 11336 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 10673 17595 10732 17601
rect 10673 17561 10685 17595
rect 10719 17564 10732 17595
rect 10873 17595 10931 17601
rect 10719 17561 10731 17564
rect 10673 17555 10731 17561
rect 10873 17561 10885 17595
rect 10919 17561 10931 17595
rect 10873 17555 10931 17561
rect 10505 17527 10563 17533
rect 10505 17524 10517 17527
rect 10060 17496 10517 17524
rect 8021 17487 8079 17493
rect 10505 17493 10517 17496
rect 10551 17493 10563 17527
rect 10888 17524 10916 17555
rect 14550 17552 14556 17604
rect 14608 17592 14614 17604
rect 15289 17595 15347 17601
rect 15289 17592 15301 17595
rect 14608 17564 15301 17592
rect 14608 17552 14614 17564
rect 15289 17561 15301 17564
rect 15335 17561 15347 17595
rect 15289 17555 15347 17561
rect 11054 17524 11060 17536
rect 10888 17496 11060 17524
rect 10505 17487 10563 17493
rect 11054 17484 11060 17496
rect 11112 17484 11118 17536
rect 15764 17524 15792 17623
rect 15948 17592 15976 17623
rect 16022 17620 16028 17672
rect 16080 17620 16086 17672
rect 23750 17620 23756 17672
rect 23808 17620 23814 17672
rect 23845 17663 23903 17669
rect 23845 17629 23857 17663
rect 23891 17660 23903 17663
rect 24118 17660 24124 17672
rect 23891 17632 24124 17660
rect 23891 17629 23903 17632
rect 23845 17623 23903 17629
rect 24118 17620 24124 17632
rect 24176 17620 24182 17672
rect 26528 17660 26556 17691
rect 28994 17688 29000 17700
rect 29052 17688 29058 17740
rect 30101 17731 30159 17737
rect 30101 17697 30113 17731
rect 30147 17728 30159 17731
rect 31846 17728 31852 17740
rect 30147 17700 31852 17728
rect 30147 17697 30159 17700
rect 30101 17691 30159 17697
rect 31846 17688 31852 17700
rect 31904 17728 31910 17740
rect 31904 17700 32444 17728
rect 31904 17688 31910 17700
rect 26789 17663 26847 17669
rect 26789 17660 26801 17663
rect 26528 17632 26801 17660
rect 26789 17629 26801 17632
rect 26835 17660 26847 17663
rect 26970 17660 26976 17672
rect 26835 17632 26976 17660
rect 26835 17629 26847 17632
rect 26789 17623 26847 17629
rect 26970 17620 26976 17632
rect 27028 17660 27034 17672
rect 32416 17669 32444 17700
rect 33778 17688 33784 17740
rect 33836 17688 33842 17740
rect 33873 17731 33931 17737
rect 33873 17697 33885 17731
rect 33919 17728 33931 17731
rect 34790 17728 34796 17740
rect 33919 17700 34796 17728
rect 33919 17697 33931 17700
rect 33873 17691 33931 17697
rect 27341 17663 27399 17669
rect 27341 17660 27353 17663
rect 27028 17632 27353 17660
rect 27028 17620 27034 17632
rect 27341 17629 27353 17632
rect 27387 17629 27399 17663
rect 27341 17623 27399 17629
rect 32401 17663 32459 17669
rect 32401 17629 32413 17663
rect 32447 17660 32459 17663
rect 33042 17660 33048 17672
rect 32447 17632 33048 17660
rect 32447 17629 32459 17632
rect 32401 17623 32459 17629
rect 33042 17620 33048 17632
rect 33100 17620 33106 17672
rect 33410 17620 33416 17672
rect 33468 17660 33474 17672
rect 33888 17660 33916 17691
rect 34790 17688 34796 17700
rect 34848 17688 34854 17740
rect 33468 17632 33916 17660
rect 33468 17620 33474 17632
rect 16482 17592 16488 17604
rect 15948 17564 16488 17592
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 17589 17595 17647 17601
rect 17589 17561 17601 17595
rect 17635 17592 17647 17595
rect 17862 17592 17868 17604
rect 17635 17564 17868 17592
rect 17635 17561 17647 17564
rect 17589 17555 17647 17561
rect 17862 17552 17868 17564
rect 17920 17552 17926 17604
rect 18046 17552 18052 17604
rect 18104 17552 18110 17604
rect 20898 17552 20904 17604
rect 20956 17552 20962 17604
rect 20990 17552 20996 17604
rect 21048 17592 21054 17604
rect 21048 17564 21390 17592
rect 21048 17552 21054 17564
rect 25590 17552 25596 17604
rect 25648 17552 25654 17604
rect 26237 17595 26295 17601
rect 26237 17561 26249 17595
rect 26283 17592 26295 17595
rect 26326 17592 26332 17604
rect 26283 17564 26332 17592
rect 26283 17561 26295 17564
rect 26237 17555 26295 17561
rect 26326 17552 26332 17564
rect 26384 17552 26390 17604
rect 28166 17552 28172 17604
rect 28224 17552 28230 17604
rect 28718 17552 28724 17604
rect 28776 17592 28782 17604
rect 28905 17595 28963 17601
rect 28905 17592 28917 17595
rect 28776 17564 28917 17592
rect 28776 17552 28782 17564
rect 28905 17561 28917 17564
rect 28951 17561 28963 17595
rect 28905 17555 28963 17561
rect 30377 17595 30435 17601
rect 30377 17561 30389 17595
rect 30423 17592 30435 17595
rect 30466 17592 30472 17604
rect 30423 17564 30472 17592
rect 30423 17561 30435 17564
rect 30377 17555 30435 17561
rect 30466 17552 30472 17564
rect 30524 17552 30530 17604
rect 30834 17552 30840 17604
rect 30892 17552 30898 17604
rect 18598 17524 18604 17536
rect 15764 17496 18604 17524
rect 18598 17484 18604 17496
rect 18656 17524 18662 17536
rect 21634 17524 21640 17536
rect 18656 17496 21640 17524
rect 18656 17484 18662 17496
rect 21634 17484 21640 17496
rect 21692 17484 21698 17536
rect 26878 17484 26884 17536
rect 26936 17524 26942 17536
rect 28813 17527 28871 17533
rect 28813 17524 28825 17527
rect 26936 17496 28825 17524
rect 26936 17484 26942 17496
rect 28813 17493 28825 17496
rect 28859 17493 28871 17527
rect 28813 17487 28871 17493
rect 33781 17527 33839 17533
rect 33781 17493 33793 17527
rect 33827 17524 33839 17527
rect 34054 17524 34060 17536
rect 33827 17496 34060 17524
rect 33827 17493 33839 17496
rect 33781 17487 33839 17493
rect 34054 17484 34060 17496
rect 34112 17484 34118 17536
rect 1104 17434 37076 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 37076 17434
rect 1104 17360 37076 17382
rect 4614 17320 4620 17332
rect 1688 17292 3280 17320
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 1688 17193 1716 17292
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 1544 17156 1685 17184
rect 1544 17144 1550 17156
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 3252 17184 3280 17292
rect 4080 17292 4620 17320
rect 3418 17212 3424 17264
rect 3476 17252 3482 17264
rect 3605 17255 3663 17261
rect 3605 17252 3617 17255
rect 3476 17224 3617 17252
rect 3476 17212 3482 17224
rect 3605 17221 3617 17224
rect 3651 17221 3663 17255
rect 3605 17215 3663 17221
rect 3786 17212 3792 17264
rect 3844 17261 3850 17264
rect 3844 17255 3863 17261
rect 3851 17221 3863 17255
rect 3844 17215 3863 17221
rect 3844 17212 3850 17215
rect 4080 17193 4108 17292
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 4706 17280 4712 17332
rect 4764 17320 4770 17332
rect 5813 17323 5871 17329
rect 5813 17320 5825 17323
rect 4764 17292 5825 17320
rect 4764 17280 4770 17292
rect 5813 17289 5825 17292
rect 5859 17289 5871 17323
rect 5813 17283 5871 17289
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 7101 17323 7159 17329
rect 7101 17320 7113 17323
rect 6604 17292 7113 17320
rect 6604 17280 6610 17292
rect 7101 17289 7113 17292
rect 7147 17289 7159 17323
rect 7101 17283 7159 17289
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 18693 17323 18751 17329
rect 18693 17320 18705 17323
rect 17920 17292 18705 17320
rect 17920 17280 17926 17292
rect 18693 17289 18705 17292
rect 18739 17289 18751 17323
rect 18693 17283 18751 17289
rect 19058 17280 19064 17332
rect 19116 17280 19122 17332
rect 22370 17280 22376 17332
rect 22428 17320 22434 17332
rect 23385 17323 23443 17329
rect 23385 17320 23397 17323
rect 22428 17292 23397 17320
rect 22428 17280 22434 17292
rect 23385 17289 23397 17292
rect 23431 17289 23443 17323
rect 26234 17320 26240 17332
rect 23385 17283 23443 17289
rect 25056 17292 26240 17320
rect 4338 17212 4344 17264
rect 4396 17212 4402 17264
rect 5626 17252 5632 17264
rect 5566 17224 5632 17252
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 6914 17212 6920 17264
rect 6972 17252 6978 17264
rect 7926 17252 7932 17264
rect 6972 17224 7932 17252
rect 6972 17212 6978 17224
rect 4065 17187 4123 17193
rect 4065 17184 4077 17187
rect 3252 17156 4077 17184
rect 4065 17153 4077 17156
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 7466 17144 7472 17196
rect 7524 17144 7530 17196
rect 7760 17193 7788 17224
rect 7926 17212 7932 17224
rect 7984 17212 7990 17264
rect 9398 17252 9404 17264
rect 9246 17224 9404 17252
rect 9398 17212 9404 17224
rect 9456 17212 9462 17264
rect 14550 17212 14556 17264
rect 14608 17212 14614 17264
rect 17586 17252 17592 17264
rect 16546 17224 17592 17252
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17153 7803 17187
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 7745 17147 7803 17153
rect 9508 17156 9781 17184
rect 1946 17076 1952 17128
rect 2004 17076 2010 17128
rect 4706 17116 4712 17128
rect 3804 17088 4712 17116
rect 3418 16940 3424 16992
rect 3476 16940 3482 16992
rect 3804 16989 3832 17088
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 7561 17119 7619 17125
rect 7561 17085 7573 17119
rect 7607 17116 7619 17119
rect 7607 17088 7880 17116
rect 7607 17085 7619 17088
rect 7561 17079 7619 17085
rect 3789 16983 3847 16989
rect 3789 16949 3801 16983
rect 3835 16949 3847 16983
rect 3789 16943 3847 16949
rect 3973 16983 4031 16989
rect 3973 16949 3985 16983
rect 4019 16980 4031 16983
rect 4522 16980 4528 16992
rect 4019 16952 4528 16980
rect 4019 16949 4031 16952
rect 3973 16943 4031 16949
rect 4522 16940 4528 16952
rect 4580 16940 4586 16992
rect 7852 16980 7880 17088
rect 8018 17076 8024 17128
rect 8076 17076 8082 17128
rect 9508 16992 9536 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 9858 17144 9864 17196
rect 9916 17184 9922 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9916 17156 9965 17184
rect 9916 17144 9922 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 11054 17184 11060 17196
rect 10459 17156 11060 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 14090 17144 14096 17196
rect 14148 17184 14154 17196
rect 14274 17184 14280 17196
rect 14148 17156 14280 17184
rect 14148 17144 14154 17156
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 16546 17184 16574 17224
rect 17586 17212 17592 17224
rect 17644 17212 17650 17264
rect 20625 17255 20683 17261
rect 20625 17221 20637 17255
rect 20671 17252 20683 17255
rect 20806 17252 20812 17264
rect 20671 17224 20812 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 20806 17212 20812 17224
rect 20864 17212 20870 17264
rect 22278 17212 22284 17264
rect 22336 17252 22342 17264
rect 22557 17255 22615 17261
rect 22557 17252 22569 17255
rect 22336 17224 22569 17252
rect 22336 17212 22342 17224
rect 22557 17221 22569 17224
rect 22603 17221 22615 17255
rect 22557 17215 22615 17221
rect 15712 17156 16574 17184
rect 15712 17144 15718 17156
rect 20438 17144 20444 17196
rect 20496 17184 20502 17196
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 20496 17156 20729 17184
rect 20496 17144 20502 17156
rect 20717 17153 20729 17156
rect 20763 17184 20775 17187
rect 20763 17156 21496 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 10502 17076 10508 17128
rect 10560 17076 10566 17128
rect 16850 17076 16856 17128
rect 16908 17076 16914 17128
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17116 17187 17119
rect 17770 17116 17776 17128
rect 17175 17088 17776 17116
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 17770 17076 17776 17088
rect 17828 17076 17834 17128
rect 18506 17076 18512 17128
rect 18564 17116 18570 17128
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 18564 17088 18613 17116
rect 18564 17076 18570 17088
rect 18601 17085 18613 17088
rect 18647 17116 18659 17119
rect 19153 17119 19211 17125
rect 19153 17116 19165 17119
rect 18647 17088 19165 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 19153 17085 19165 17088
rect 19199 17085 19211 17119
rect 19153 17079 19211 17085
rect 19337 17119 19395 17125
rect 19337 17085 19349 17119
rect 19383 17116 19395 17119
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 19383 17088 20821 17116
rect 19383 17085 19395 17088
rect 19337 17079 19395 17085
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 21468 17116 21496 17156
rect 21818 17144 21824 17196
rect 21876 17144 21882 17196
rect 25056 17193 25084 17292
rect 26234 17280 26240 17292
rect 26292 17280 26298 17332
rect 26789 17323 26847 17329
rect 26789 17289 26801 17323
rect 26835 17320 26847 17323
rect 26878 17320 26884 17332
rect 26835 17292 26884 17320
rect 26835 17289 26847 17292
rect 26789 17283 26847 17289
rect 26878 17280 26884 17292
rect 26936 17280 26942 17332
rect 34054 17280 34060 17332
rect 34112 17320 34118 17332
rect 35713 17323 35771 17329
rect 35713 17320 35725 17323
rect 34112 17292 35725 17320
rect 34112 17280 34118 17292
rect 35713 17289 35725 17292
rect 35759 17289 35771 17323
rect 35713 17283 35771 17289
rect 25590 17212 25596 17264
rect 25648 17252 25654 17264
rect 25648 17224 25806 17252
rect 25648 17212 25654 17224
rect 28810 17212 28816 17264
rect 28868 17252 28874 17264
rect 29733 17255 29791 17261
rect 29733 17252 29745 17255
rect 28868 17224 29745 17252
rect 28868 17212 28874 17224
rect 29733 17221 29745 17224
rect 29779 17221 29791 17255
rect 29733 17215 29791 17221
rect 30650 17212 30656 17264
rect 30708 17212 30714 17264
rect 31665 17255 31723 17261
rect 31665 17221 31677 17255
rect 31711 17252 31723 17255
rect 31754 17252 31760 17264
rect 31711 17224 31760 17252
rect 31711 17221 31723 17224
rect 31665 17215 31723 17221
rect 31754 17212 31760 17224
rect 31812 17212 31818 17264
rect 33704 17224 34730 17252
rect 25041 17187 25099 17193
rect 25041 17153 25053 17187
rect 25087 17153 25099 17187
rect 25041 17147 25099 17153
rect 28994 17144 29000 17196
rect 29052 17144 29058 17196
rect 29546 17144 29552 17196
rect 29604 17144 29610 17196
rect 31938 17144 31944 17196
rect 31996 17144 32002 17196
rect 33502 17144 33508 17196
rect 33560 17184 33566 17196
rect 33704 17184 33732 17224
rect 33560 17156 33732 17184
rect 33560 17144 33566 17156
rect 23293 17119 23351 17125
rect 23293 17116 23305 17119
rect 21468 17088 23305 17116
rect 20809 17079 20867 17085
rect 23293 17085 23305 17088
rect 23339 17085 23351 17119
rect 23293 17079 23351 17085
rect 23477 17119 23535 17125
rect 23477 17085 23489 17119
rect 23523 17085 23535 17119
rect 23477 17079 23535 17085
rect 25317 17119 25375 17125
rect 25317 17085 25329 17119
rect 25363 17116 25375 17119
rect 26786 17116 26792 17128
rect 25363 17088 26792 17116
rect 25363 17085 25375 17088
rect 25317 17079 25375 17085
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 19352 17048 19380 17079
rect 18288 17020 19380 17048
rect 18288 17008 18294 17020
rect 21634 17008 21640 17060
rect 21692 17048 21698 17060
rect 23492 17048 23520 17079
rect 26786 17076 26792 17088
rect 26844 17076 26850 17128
rect 29822 17076 29828 17128
rect 29880 17116 29886 17128
rect 29880 17088 32076 17116
rect 29880 17076 29886 17088
rect 21692 17020 23520 17048
rect 21692 17008 21698 17020
rect 8570 16980 8576 16992
rect 7852 16952 8576 16980
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9490 16940 9496 16992
rect 9548 16940 9554 16992
rect 9582 16940 9588 16992
rect 9640 16940 9646 16992
rect 10781 16983 10839 16989
rect 10781 16949 10793 16983
rect 10827 16980 10839 16983
rect 10870 16980 10876 16992
rect 10827 16952 10876 16980
rect 10827 16949 10839 16952
rect 10781 16943 10839 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16390 16980 16396 16992
rect 16080 16952 16396 16980
rect 16080 16940 16086 16952
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 16482 16940 16488 16992
rect 16540 16980 16546 16992
rect 18248 16980 18276 17008
rect 16540 16952 18276 16980
rect 16540 16940 16546 16952
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 20257 16983 20315 16989
rect 20257 16980 20269 16983
rect 19392 16952 20269 16980
rect 19392 16940 19398 16952
rect 20257 16949 20269 16952
rect 20303 16949 20315 16983
rect 20257 16943 20315 16949
rect 21910 16940 21916 16992
rect 21968 16980 21974 16992
rect 22925 16983 22983 16989
rect 22925 16980 22937 16983
rect 21968 16952 22937 16980
rect 21968 16940 21974 16952
rect 22925 16949 22937 16952
rect 22971 16949 22983 16983
rect 22925 16943 22983 16949
rect 27798 16940 27804 16992
rect 27856 16980 27862 16992
rect 29273 16983 29331 16989
rect 29273 16980 29285 16983
rect 27856 16952 29285 16980
rect 27856 16940 27862 16952
rect 29273 16949 29285 16952
rect 29319 16949 29331 16983
rect 29273 16943 29331 16949
rect 30193 16983 30251 16989
rect 30193 16949 30205 16983
rect 30239 16980 30251 16983
rect 31202 16980 31208 16992
rect 30239 16952 31208 16980
rect 30239 16949 30251 16952
rect 30193 16943 30251 16949
rect 31202 16940 31208 16952
rect 31260 16980 31266 16992
rect 31938 16980 31944 16992
rect 31260 16952 31944 16980
rect 31260 16940 31266 16952
rect 31938 16940 31944 16952
rect 31996 16940 32002 16992
rect 32048 16980 32076 17088
rect 32122 17076 32128 17128
rect 32180 17076 32186 17128
rect 32398 17076 32404 17128
rect 32456 17076 32462 17128
rect 33042 17076 33048 17128
rect 33100 17116 33106 17128
rect 33965 17119 34023 17125
rect 33965 17116 33977 17119
rect 33100 17088 33977 17116
rect 33100 17076 33106 17088
rect 33965 17085 33977 17088
rect 34011 17085 34023 17119
rect 33965 17079 34023 17085
rect 34238 17076 34244 17128
rect 34296 17076 34302 17128
rect 33410 16980 33416 16992
rect 32048 16952 33416 16980
rect 33410 16940 33416 16952
rect 33468 16940 33474 16992
rect 33502 16940 33508 16992
rect 33560 16980 33566 16992
rect 33873 16983 33931 16989
rect 33873 16980 33885 16983
rect 33560 16952 33885 16980
rect 33560 16940 33566 16952
rect 33873 16949 33885 16952
rect 33919 16949 33931 16983
rect 33873 16943 33931 16949
rect 1104 16890 37076 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 37076 16890
rect 1104 16816 37076 16838
rect 1765 16779 1823 16785
rect 1765 16745 1777 16779
rect 1811 16776 1823 16779
rect 1946 16776 1952 16788
rect 1811 16748 1952 16776
rect 1811 16745 1823 16748
rect 1765 16739 1823 16745
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 4430 16736 4436 16788
rect 4488 16776 4494 16788
rect 5258 16776 5264 16788
rect 4488 16748 5264 16776
rect 4488 16736 4494 16748
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 8297 16779 8355 16785
rect 8297 16776 8309 16779
rect 8076 16748 8309 16776
rect 8076 16736 8082 16748
rect 8297 16745 8309 16748
rect 8343 16745 8355 16779
rect 9582 16776 9588 16788
rect 8297 16739 8355 16745
rect 8496 16748 9588 16776
rect 4798 16708 4804 16720
rect 4172 16680 4804 16708
rect 2222 16600 2228 16652
rect 2280 16600 2286 16652
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 3418 16572 3424 16584
rect 2179 16544 3424 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 3418 16532 3424 16544
rect 3476 16532 3482 16584
rect 3789 16575 3847 16581
rect 3789 16541 3801 16575
rect 3835 16572 3847 16575
rect 3970 16572 3976 16584
rect 3835 16544 3976 16572
rect 3835 16541 3847 16544
rect 3789 16535 3847 16541
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4062 16532 4068 16584
rect 4120 16532 4126 16584
rect 4172 16581 4200 16680
rect 4798 16668 4804 16680
rect 4856 16668 4862 16720
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 4264 16612 4537 16640
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 3881 16507 3939 16513
rect 3881 16473 3893 16507
rect 3927 16504 3939 16507
rect 4264 16504 4292 16612
rect 4525 16609 4537 16612
rect 4571 16609 4583 16643
rect 4525 16603 4583 16609
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 5169 16643 5227 16649
rect 5169 16640 5181 16643
rect 4672 16612 5181 16640
rect 4672 16600 4678 16612
rect 5169 16609 5181 16612
rect 5215 16609 5227 16643
rect 5169 16603 5227 16609
rect 4430 16532 4436 16584
rect 4488 16532 4494 16584
rect 8496 16581 8524 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 12345 16779 12403 16785
rect 12345 16776 12357 16779
rect 11112 16748 12357 16776
rect 11112 16736 11118 16748
rect 12345 16745 12357 16748
rect 12391 16745 12403 16779
rect 12345 16739 12403 16745
rect 20438 16736 20444 16788
rect 20496 16736 20502 16788
rect 25120 16779 25178 16785
rect 25120 16745 25132 16779
rect 25166 16776 25178 16779
rect 25682 16776 25688 16788
rect 25166 16748 25688 16776
rect 25166 16745 25178 16748
rect 25120 16739 25178 16745
rect 25682 16736 25688 16748
rect 25740 16736 25746 16788
rect 26786 16736 26792 16788
rect 26844 16736 26850 16788
rect 27062 16736 27068 16788
rect 27120 16776 27126 16788
rect 29273 16779 29331 16785
rect 27120 16748 28994 16776
rect 27120 16736 27126 16748
rect 9490 16708 9496 16720
rect 8956 16680 9496 16708
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 4801 16575 4859 16581
rect 4801 16572 4813 16575
rect 4755 16544 4813 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 4801 16541 4813 16544
rect 4847 16541 4859 16575
rect 4801 16535 4859 16541
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 8956 16581 8984 16680
rect 9490 16668 9496 16680
rect 9548 16668 9554 16720
rect 28966 16708 28994 16748
rect 29273 16745 29285 16779
rect 29319 16776 29331 16779
rect 29546 16776 29552 16788
rect 29319 16748 29552 16776
rect 29319 16745 29331 16748
rect 29273 16739 29331 16745
rect 29546 16736 29552 16748
rect 29604 16736 29610 16788
rect 33502 16776 33508 16788
rect 31680 16748 33508 16776
rect 30837 16711 30895 16717
rect 30837 16708 30849 16711
rect 28966 16680 30849 16708
rect 30837 16677 30849 16680
rect 30883 16677 30895 16711
rect 30837 16671 30895 16677
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 10594 16640 10600 16652
rect 10100 16612 10600 16640
rect 10100 16600 10106 16612
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10870 16600 10876 16652
rect 10928 16600 10934 16652
rect 14090 16600 14096 16652
rect 14148 16600 14154 16652
rect 14369 16643 14427 16649
rect 14369 16609 14381 16643
rect 14415 16640 14427 16643
rect 15930 16640 15936 16652
rect 14415 16612 15936 16640
rect 14415 16609 14427 16612
rect 14369 16603 14427 16609
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16640 16635 16643
rect 18966 16640 18972 16652
rect 16623 16612 18972 16640
rect 16623 16609 16635 16612
rect 16577 16603 16635 16609
rect 18966 16600 18972 16612
rect 19024 16600 19030 16652
rect 21910 16600 21916 16652
rect 21968 16600 21974 16652
rect 22189 16643 22247 16649
rect 22189 16609 22201 16643
rect 22235 16640 22247 16643
rect 22278 16640 22284 16652
rect 22235 16612 22284 16640
rect 22235 16609 22247 16612
rect 22189 16603 22247 16609
rect 22278 16600 22284 16612
rect 22336 16640 22342 16652
rect 22373 16643 22431 16649
rect 22373 16640 22385 16643
rect 22336 16612 22385 16640
rect 22336 16600 22342 16612
rect 22373 16609 22385 16612
rect 22419 16609 22431 16643
rect 22373 16603 22431 16609
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16640 24915 16643
rect 26142 16640 26148 16652
rect 24903 16612 26148 16640
rect 24903 16609 24915 16612
rect 24857 16603 24915 16609
rect 26142 16600 26148 16612
rect 26200 16640 26206 16652
rect 27522 16640 27528 16652
rect 26200 16612 27528 16640
rect 26200 16600 26206 16612
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 27798 16600 27804 16652
rect 27856 16600 27862 16652
rect 29012 16612 29316 16640
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16572 9183 16575
rect 9858 16572 9864 16584
rect 9171 16544 9864 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 17770 16532 17776 16584
rect 17828 16532 17834 16584
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 3927 16476 4292 16504
rect 4893 16507 4951 16513
rect 3927 16473 3939 16476
rect 3881 16467 3939 16473
rect 4893 16473 4905 16507
rect 4939 16504 4951 16507
rect 5445 16507 5503 16513
rect 5445 16504 5457 16507
rect 4939 16476 5457 16504
rect 4939 16473 4951 16476
rect 4893 16467 4951 16473
rect 5445 16473 5457 16476
rect 5491 16473 5503 16507
rect 5445 16467 5503 16473
rect 5534 16464 5540 16516
rect 5592 16504 5598 16516
rect 7193 16507 7251 16513
rect 5592 16476 5934 16504
rect 5592 16464 5598 16476
rect 7193 16473 7205 16507
rect 7239 16504 7251 16507
rect 7282 16504 7288 16516
rect 7239 16476 7288 16504
rect 7239 16473 7251 16476
rect 7193 16467 7251 16473
rect 7282 16464 7288 16476
rect 7340 16464 7346 16516
rect 8588 16504 8616 16532
rect 9033 16507 9091 16513
rect 9033 16504 9045 16507
rect 8588 16476 9045 16504
rect 9033 16473 9045 16476
rect 9079 16473 9091 16507
rect 9033 16467 9091 16473
rect 9398 16464 9404 16516
rect 9456 16504 9462 16516
rect 11330 16504 11336 16516
rect 9456 16476 11336 16504
rect 9456 16464 9462 16476
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 15654 16504 15660 16516
rect 15594 16476 15660 16504
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 17310 16464 17316 16516
rect 17368 16464 17374 16516
rect 18248 16504 18276 16535
rect 18414 16532 18420 16584
rect 18472 16532 18478 16584
rect 18506 16532 18512 16584
rect 18564 16532 18570 16584
rect 26878 16532 26884 16584
rect 26936 16572 26942 16584
rect 27065 16575 27123 16581
rect 27065 16572 27077 16575
rect 26936 16544 27077 16572
rect 26936 16532 26942 16544
rect 27065 16541 27077 16544
rect 27111 16541 27123 16575
rect 29012 16572 29040 16612
rect 28934 16544 29040 16572
rect 29288 16572 29316 16612
rect 30650 16572 30656 16584
rect 29288 16544 30656 16572
rect 27065 16535 27123 16541
rect 30650 16532 30656 16544
rect 30708 16532 30714 16584
rect 20622 16504 20628 16516
rect 18248 16476 20628 16504
rect 20622 16464 20628 16476
rect 20680 16464 20686 16516
rect 20898 16464 20904 16516
rect 20956 16464 20962 16516
rect 22646 16464 22652 16516
rect 22704 16464 22710 16516
rect 23934 16504 23940 16516
rect 23874 16476 23940 16504
rect 23934 16464 23940 16476
rect 23992 16504 23998 16516
rect 25590 16504 25596 16516
rect 23992 16476 25176 16504
rect 23992 16464 23998 16476
rect 4341 16439 4399 16445
rect 4341 16405 4353 16439
rect 4387 16436 4399 16439
rect 4706 16436 4712 16448
rect 4387 16408 4712 16436
rect 4387 16405 4399 16408
rect 4341 16399 4399 16405
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 15838 16396 15844 16448
rect 15896 16396 15902 16448
rect 24121 16439 24179 16445
rect 24121 16405 24133 16439
rect 24167 16436 24179 16439
rect 25038 16436 25044 16448
rect 24167 16408 25044 16436
rect 24167 16405 24179 16408
rect 24121 16399 24179 16405
rect 25038 16396 25044 16408
rect 25096 16396 25102 16448
rect 25148 16436 25176 16476
rect 25516 16476 25596 16504
rect 25516 16436 25544 16476
rect 25590 16464 25596 16476
rect 25648 16464 25654 16516
rect 27341 16507 27399 16513
rect 27341 16473 27353 16507
rect 27387 16473 27399 16507
rect 27341 16467 27399 16473
rect 25148 16408 25544 16436
rect 25958 16396 25964 16448
rect 26016 16436 26022 16448
rect 26605 16439 26663 16445
rect 26605 16436 26617 16439
rect 26016 16408 26617 16436
rect 26016 16396 26022 16408
rect 26605 16405 26617 16408
rect 26651 16436 26663 16439
rect 27249 16439 27307 16445
rect 27249 16436 27261 16439
rect 26651 16408 27261 16436
rect 26651 16405 26663 16408
rect 26605 16399 26663 16405
rect 27249 16405 27261 16408
rect 27295 16405 27307 16439
rect 27356 16436 27384 16467
rect 29270 16464 29276 16516
rect 29328 16504 29334 16516
rect 29549 16507 29607 16513
rect 29549 16504 29561 16507
rect 29328 16476 29561 16504
rect 29328 16464 29334 16476
rect 29549 16473 29561 16476
rect 29595 16473 29607 16507
rect 30852 16504 30880 16671
rect 31680 16649 31708 16748
rect 33502 16736 33508 16748
rect 33560 16736 33566 16788
rect 31754 16668 31760 16720
rect 31812 16708 31818 16720
rect 32122 16708 32128 16720
rect 31812 16680 32128 16708
rect 31812 16668 31818 16680
rect 32122 16668 32128 16680
rect 32180 16708 32186 16720
rect 32180 16680 34284 16708
rect 32180 16668 32186 16680
rect 31665 16643 31723 16649
rect 31665 16609 31677 16643
rect 31711 16609 31723 16643
rect 32030 16640 32036 16652
rect 31665 16603 31723 16609
rect 31772 16612 32036 16640
rect 31772 16581 31800 16612
rect 32030 16600 32036 16612
rect 32088 16600 32094 16652
rect 32398 16600 32404 16652
rect 32456 16600 32462 16652
rect 32677 16643 32735 16649
rect 32677 16609 32689 16643
rect 32723 16640 32735 16643
rect 33042 16640 33048 16652
rect 32723 16612 33048 16640
rect 32723 16609 32735 16612
rect 32677 16603 32735 16609
rect 33042 16600 33048 16612
rect 33100 16600 33106 16652
rect 34256 16649 34284 16680
rect 34241 16643 34299 16649
rect 34241 16609 34253 16643
rect 34287 16609 34299 16643
rect 34241 16603 34299 16609
rect 36446 16600 36452 16652
rect 36504 16600 36510 16652
rect 31757 16575 31815 16581
rect 31757 16541 31769 16575
rect 31803 16541 31815 16575
rect 31757 16535 31815 16541
rect 31938 16532 31944 16584
rect 31996 16532 32002 16584
rect 31662 16504 31668 16516
rect 30852 16476 31668 16504
rect 29549 16467 29607 16473
rect 31662 16464 31668 16476
rect 31720 16464 31726 16516
rect 33413 16507 33471 16513
rect 33413 16473 33425 16507
rect 33459 16504 33471 16507
rect 33505 16507 33563 16513
rect 33505 16504 33517 16507
rect 33459 16476 33517 16504
rect 33459 16473 33471 16476
rect 33413 16467 33471 16473
rect 33505 16473 33517 16476
rect 33551 16473 33563 16507
rect 33505 16467 33563 16473
rect 29822 16436 29828 16448
rect 27356 16408 29828 16436
rect 27249 16399 27307 16405
rect 29822 16396 29828 16408
rect 29880 16396 29886 16448
rect 29914 16396 29920 16448
rect 29972 16436 29978 16448
rect 33428 16436 33456 16467
rect 36630 16464 36636 16516
rect 36688 16464 36694 16516
rect 29972 16408 33456 16436
rect 29972 16396 29978 16408
rect 1104 16346 37076 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 37076 16346
rect 1104 16272 37076 16294
rect 3418 16192 3424 16244
rect 3476 16232 3482 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 3476 16204 3893 16232
rect 3476 16192 3482 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 4062 16192 4068 16244
rect 4120 16192 4126 16244
rect 17126 16232 17132 16244
rect 15212 16204 17132 16232
rect 2332 16136 3924 16164
rect 2222 16056 2228 16108
rect 2280 16105 2286 16108
rect 2280 16096 2289 16105
rect 2332 16096 2360 16136
rect 3896 16108 3924 16136
rect 10502 16124 10508 16176
rect 10560 16124 10566 16176
rect 2280 16068 2360 16096
rect 2409 16099 2467 16105
rect 2280 16059 2289 16068
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 3418 16096 3424 16108
rect 2455 16068 3424 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2280 16056 2286 16059
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 3694 16056 3700 16108
rect 3752 16056 3758 16108
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16065 3847 16099
rect 3789 16059 3847 16065
rect 3804 16028 3832 16059
rect 3878 16056 3884 16108
rect 3936 16056 3942 16108
rect 14274 16056 14280 16108
rect 14332 16096 14338 16108
rect 15212 16105 15240 16204
rect 17126 16192 17132 16204
rect 17184 16192 17190 16244
rect 19518 16232 19524 16244
rect 19076 16204 19524 16232
rect 15654 16124 15660 16176
rect 15712 16164 15718 16176
rect 15712 16136 16974 16164
rect 15712 16124 15718 16136
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 14332 16068 14657 16096
rect 14332 16056 14338 16068
rect 14645 16065 14657 16068
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15286 16096 15292 16108
rect 15243 16068 15292 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 15838 16096 15844 16108
rect 15427 16068 15844 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16096 18475 16099
rect 18598 16096 18604 16108
rect 18463 16068 18604 16096
rect 18463 16065 18475 16068
rect 18417 16059 18475 16065
rect 18598 16056 18604 16068
rect 18656 16096 18662 16108
rect 18966 16096 18972 16108
rect 18656 16068 18972 16096
rect 18656 16056 18662 16068
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 19076 16105 19104 16204
rect 19518 16192 19524 16204
rect 19576 16192 19582 16244
rect 20806 16192 20812 16244
rect 20864 16192 20870 16244
rect 21818 16192 21824 16244
rect 21876 16232 21882 16244
rect 26602 16232 26608 16244
rect 21876 16204 26608 16232
rect 21876 16192 21882 16204
rect 26602 16192 26608 16204
rect 26660 16232 26666 16244
rect 28166 16232 28172 16244
rect 26660 16204 28172 16232
rect 26660 16192 26666 16204
rect 19334 16124 19340 16176
rect 19392 16124 19398 16176
rect 22646 16124 22652 16176
rect 22704 16124 22710 16176
rect 23934 16124 23940 16176
rect 23992 16164 23998 16176
rect 23992 16136 24518 16164
rect 23992 16124 23998 16136
rect 25958 16124 25964 16176
rect 26016 16124 26022 16176
rect 26988 16173 27016 16204
rect 28166 16192 28172 16204
rect 28224 16192 28230 16244
rect 29086 16192 29092 16244
rect 29144 16232 29150 16244
rect 30377 16235 30435 16241
rect 30377 16232 30389 16235
rect 29144 16204 30389 16232
rect 29144 16192 29150 16204
rect 30377 16201 30389 16204
rect 30423 16232 30435 16235
rect 32677 16235 32735 16241
rect 32677 16232 32689 16235
rect 30423 16204 32689 16232
rect 30423 16201 30435 16204
rect 30377 16195 30435 16201
rect 32677 16201 32689 16204
rect 32723 16201 32735 16235
rect 32677 16195 32735 16201
rect 33502 16192 33508 16244
rect 33560 16192 33566 16244
rect 33965 16235 34023 16241
rect 33965 16201 33977 16235
rect 34011 16232 34023 16235
rect 34238 16232 34244 16244
rect 34011 16204 34244 16232
rect 34011 16201 34023 16204
rect 33965 16195 34023 16201
rect 34238 16192 34244 16204
rect 34296 16192 34302 16244
rect 26145 16167 26203 16173
rect 26145 16133 26157 16167
rect 26191 16133 26203 16167
rect 26145 16127 26203 16133
rect 26973 16167 27031 16173
rect 26973 16133 26985 16167
rect 27019 16133 27031 16167
rect 26973 16127 27031 16133
rect 19061 16099 19119 16105
rect 19061 16065 19073 16099
rect 19107 16065 19119 16099
rect 21637 16099 21695 16105
rect 19061 16059 19119 16065
rect 4062 16028 4068 16040
rect 3804 16000 4068 16028
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 16028 7527 16031
rect 7650 16028 7656 16040
rect 7515 16000 7656 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 14366 15988 14372 16040
rect 14424 16028 14430 16040
rect 14737 16031 14795 16037
rect 14737 16028 14749 16031
rect 14424 16000 14749 16028
rect 14424 15988 14430 16000
rect 14737 15997 14749 16000
rect 14783 15997 14795 16031
rect 14737 15991 14795 15997
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 18141 16031 18199 16037
rect 18141 15997 18153 16031
rect 18187 16028 18199 16031
rect 18782 16028 18788 16040
rect 18187 16000 18788 16028
rect 18187 15997 18199 16000
rect 18141 15991 18199 15997
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 19978 15988 19984 16040
rect 20036 16028 20042 16040
rect 20456 16028 20484 16082
rect 21637 16065 21649 16099
rect 21683 16096 21695 16099
rect 21818 16096 21824 16108
rect 21683 16068 21824 16096
rect 21683 16065 21695 16068
rect 21637 16059 21695 16065
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 23106 16056 23112 16108
rect 23164 16056 23170 16108
rect 23290 16056 23296 16108
rect 23348 16056 23354 16108
rect 20898 16028 20904 16040
rect 20036 16000 20904 16028
rect 20036 15988 20042 16000
rect 20898 15988 20904 16000
rect 20956 15988 20962 16040
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 3142 15920 3148 15972
rect 3200 15960 3206 15972
rect 3513 15963 3571 15969
rect 3513 15960 3525 15963
rect 3200 15932 3525 15960
rect 3200 15920 3206 15932
rect 3513 15929 3525 15932
rect 3559 15929 3571 15963
rect 3513 15923 3571 15929
rect 7101 15963 7159 15969
rect 7101 15929 7113 15963
rect 7147 15960 7159 15963
rect 7742 15960 7748 15972
rect 7147 15932 7748 15960
rect 7147 15929 7159 15932
rect 7101 15923 7159 15929
rect 7742 15920 7748 15932
rect 7800 15920 7806 15972
rect 10781 15963 10839 15969
rect 10781 15929 10793 15963
rect 10827 15960 10839 15963
rect 11054 15960 11060 15972
rect 10827 15932 11060 15960
rect 10827 15929 10839 15932
rect 10781 15923 10839 15929
rect 11054 15920 11060 15932
rect 11112 15920 11118 15972
rect 1670 15852 1676 15904
rect 1728 15892 1734 15904
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 1728 15864 2421 15892
rect 1728 15852 1734 15864
rect 2409 15861 2421 15864
rect 2455 15861 2467 15895
rect 2409 15855 2467 15861
rect 7009 15895 7067 15901
rect 7009 15861 7021 15895
rect 7055 15892 7067 15895
rect 7190 15892 7196 15904
rect 7055 15864 7196 15892
rect 7055 15861 7067 15864
rect 7009 15855 7067 15861
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 10928 15864 10977 15892
rect 10928 15852 10934 15864
rect 10965 15861 10977 15864
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 16669 15895 16727 15901
rect 16669 15861 16681 15895
rect 16715 15892 16727 15895
rect 18414 15892 18420 15904
rect 16715 15864 18420 15892
rect 16715 15861 16727 15864
rect 16669 15855 16727 15861
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 23400 15892 23428 15991
rect 23750 15988 23756 16040
rect 23808 15988 23814 16040
rect 24029 16031 24087 16037
rect 24029 15997 24041 16031
rect 24075 16028 24087 16031
rect 24394 16028 24400 16040
rect 24075 16000 24400 16028
rect 24075 15997 24087 16000
rect 24029 15991 24087 15997
rect 24394 15988 24400 16000
rect 24452 15988 24458 16040
rect 25498 15988 25504 16040
rect 25556 16028 25562 16040
rect 26160 16028 26188 16127
rect 27522 16124 27528 16176
rect 27580 16164 27586 16176
rect 27709 16167 27767 16173
rect 27709 16164 27721 16167
rect 27580 16136 27721 16164
rect 27580 16124 27586 16136
rect 27709 16133 27721 16136
rect 27755 16133 27767 16167
rect 28994 16164 29000 16176
rect 27709 16127 27767 16133
rect 28644 16136 29000 16164
rect 27724 16096 27752 16127
rect 28644 16105 28672 16136
rect 28994 16124 29000 16136
rect 29052 16124 29058 16176
rect 30650 16164 30656 16176
rect 30130 16136 30656 16164
rect 30650 16124 30656 16136
rect 30708 16124 30714 16176
rect 33597 16167 33655 16173
rect 33597 16133 33609 16167
rect 33643 16164 33655 16167
rect 34054 16164 34060 16176
rect 33643 16136 34060 16164
rect 33643 16133 33655 16136
rect 33597 16127 33655 16133
rect 34054 16124 34060 16136
rect 34112 16124 34118 16176
rect 28629 16099 28687 16105
rect 28629 16096 28641 16099
rect 27724 16068 28641 16096
rect 28629 16065 28641 16068
rect 28675 16065 28687 16099
rect 28629 16059 28687 16065
rect 30469 16099 30527 16105
rect 30469 16065 30481 16099
rect 30515 16065 30527 16099
rect 30469 16059 30527 16065
rect 25556 16000 26188 16028
rect 26237 16031 26295 16037
rect 25556 15988 25562 16000
rect 26237 15997 26249 16031
rect 26283 16028 26295 16031
rect 26326 16028 26332 16040
rect 26283 16000 26332 16028
rect 26283 15997 26295 16000
rect 26237 15991 26295 15997
rect 26326 15988 26332 16000
rect 26384 16028 26390 16040
rect 28534 16028 28540 16040
rect 26384 16000 28540 16028
rect 26384 15988 26390 16000
rect 28534 15988 28540 16000
rect 28592 15988 28598 16040
rect 28902 15988 28908 16040
rect 28960 15988 28966 16040
rect 29270 15988 29276 16040
rect 29328 16028 29334 16040
rect 30484 16028 30512 16059
rect 31754 16056 31760 16108
rect 31812 16056 31818 16108
rect 29328 16000 30512 16028
rect 29328 15988 29334 16000
rect 30834 15988 30840 16040
rect 30892 15988 30898 16040
rect 31938 15988 31944 16040
rect 31996 16028 32002 16040
rect 32585 16031 32643 16037
rect 32585 16028 32597 16031
rect 31996 16000 32597 16028
rect 31996 15988 32002 16000
rect 32585 15997 32597 16000
rect 32631 15997 32643 16031
rect 32585 15991 32643 15997
rect 32766 15988 32772 16040
rect 32824 15988 32830 16040
rect 33134 15988 33140 16040
rect 33192 16028 33198 16040
rect 33321 16031 33379 16037
rect 33321 16028 33333 16031
rect 33192 16000 33333 16028
rect 33192 15988 33198 16000
rect 33321 15997 33333 16000
rect 33367 15997 33379 16031
rect 33321 15991 33379 15997
rect 25682 15920 25688 15972
rect 25740 15920 25746 15972
rect 25038 15892 25044 15904
rect 23400 15864 25044 15892
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 28166 15852 28172 15904
rect 28224 15892 28230 15904
rect 29914 15892 29920 15904
rect 28224 15864 29920 15892
rect 28224 15852 28230 15864
rect 29914 15852 29920 15864
rect 29972 15852 29978 15904
rect 32214 15852 32220 15904
rect 32272 15852 32278 15904
rect 1104 15802 37076 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 37076 15802
rect 1104 15728 37076 15750
rect 3418 15648 3424 15700
rect 3476 15648 3482 15700
rect 3878 15648 3884 15700
rect 3936 15688 3942 15700
rect 4341 15691 4399 15697
rect 4341 15688 4353 15691
rect 3936 15660 4353 15688
rect 3936 15648 3942 15660
rect 4341 15657 4353 15660
rect 4387 15657 4399 15691
rect 4341 15651 4399 15657
rect 10502 15648 10508 15700
rect 10560 15648 10566 15700
rect 15470 15648 15476 15700
rect 15528 15688 15534 15700
rect 15654 15688 15660 15700
rect 15528 15660 15660 15688
rect 15528 15648 15534 15660
rect 15654 15648 15660 15660
rect 15712 15688 15718 15700
rect 15841 15691 15899 15697
rect 15841 15688 15853 15691
rect 15712 15660 15853 15688
rect 15712 15648 15718 15660
rect 15841 15657 15853 15660
rect 15887 15657 15899 15691
rect 15841 15651 15899 15657
rect 15930 15648 15936 15700
rect 15988 15648 15994 15700
rect 23290 15648 23296 15700
rect 23348 15688 23354 15700
rect 23569 15691 23627 15697
rect 23569 15688 23581 15691
rect 23348 15660 23581 15688
rect 23348 15648 23354 15660
rect 23569 15657 23581 15660
rect 23615 15657 23627 15691
rect 23569 15651 23627 15657
rect 28721 15691 28779 15697
rect 28721 15657 28733 15691
rect 28767 15688 28779 15691
rect 28902 15688 28908 15700
rect 28767 15660 28908 15688
rect 28767 15657 28779 15660
rect 28721 15651 28779 15657
rect 28902 15648 28908 15660
rect 28960 15648 28966 15700
rect 31297 15623 31355 15629
rect 17144 15592 18552 15620
rect 1670 15512 1676 15564
rect 1728 15512 1734 15564
rect 3145 15555 3203 15561
rect 3145 15521 3157 15555
rect 3191 15552 3203 15555
rect 3191 15524 4108 15552
rect 3191 15521 3203 15524
rect 3145 15515 3203 15521
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 3252 15493 3280 15524
rect 4080 15496 4108 15524
rect 7190 15512 7196 15564
rect 7248 15512 7254 15564
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 7708 15524 9812 15552
rect 7708 15512 7714 15524
rect 3237 15487 3295 15493
rect 3237 15453 3249 15487
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15484 3479 15487
rect 3510 15484 3516 15496
rect 3467 15456 3516 15484
rect 3467 15453 3479 15456
rect 3421 15447 3479 15453
rect 3510 15444 3516 15456
rect 3568 15444 3574 15496
rect 4062 15444 4068 15496
rect 4120 15444 4126 15496
rect 6914 15444 6920 15496
rect 6972 15444 6978 15496
rect 3050 15416 3056 15428
rect 2898 15388 3056 15416
rect 3050 15376 3056 15388
rect 3108 15376 3114 15428
rect 3142 15376 3148 15428
rect 3200 15416 3206 15428
rect 3789 15419 3847 15425
rect 3789 15416 3801 15419
rect 3200 15388 3801 15416
rect 3200 15376 3206 15388
rect 3789 15385 3801 15388
rect 3835 15385 3847 15419
rect 3789 15379 3847 15385
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 9232 15416 9260 15524
rect 9784 15493 9812 15524
rect 10594 15512 10600 15564
rect 10652 15512 10658 15564
rect 10870 15512 10876 15564
rect 10928 15512 10934 15564
rect 14366 15512 14372 15564
rect 14424 15512 14430 15564
rect 15562 15552 15568 15564
rect 15488 15524 15568 15552
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9585 15487 9643 15493
rect 9585 15484 9597 15487
rect 9355 15456 9597 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 9585 15453 9597 15456
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15484 9827 15487
rect 10318 15484 10324 15496
rect 9815 15456 10324 15484
rect 9815 15453 9827 15456
rect 9769 15447 9827 15453
rect 9493 15419 9551 15425
rect 9493 15416 9505 15419
rect 5592 15388 7682 15416
rect 9232 15388 9505 15416
rect 5592 15376 5598 15388
rect 9493 15385 9505 15388
rect 9539 15385 9551 15419
rect 9600 15416 9628 15447
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15453 14151 15487
rect 15488 15470 15516 15524
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 16390 15512 16396 15564
rect 16448 15512 16454 15564
rect 16482 15512 16488 15564
rect 16540 15512 16546 15564
rect 16850 15512 16856 15564
rect 16908 15512 16914 15564
rect 14093 15447 14151 15453
rect 9953 15419 10011 15425
rect 9953 15416 9965 15419
rect 9600 15388 9965 15416
rect 9493 15379 9551 15385
rect 9953 15385 9965 15388
rect 9999 15416 10011 15419
rect 10042 15416 10048 15428
rect 9999 15388 10048 15416
rect 9999 15385 10011 15388
rect 9953 15379 10011 15385
rect 10042 15376 10048 15388
rect 10100 15376 10106 15428
rect 10229 15419 10287 15425
rect 10229 15385 10241 15419
rect 10275 15416 10287 15419
rect 10275 15388 10640 15416
rect 10275 15385 10287 15388
rect 10229 15379 10287 15385
rect 10612 15360 10640 15388
rect 11330 15376 11336 15428
rect 11388 15376 11394 15428
rect 14108 15416 14136 15447
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 16301 15487 16359 15493
rect 16301 15484 16313 15487
rect 15896 15456 16313 15484
rect 15896 15444 15902 15456
rect 16301 15453 16313 15456
rect 16347 15453 16359 15487
rect 16301 15447 16359 15453
rect 14274 15416 14280 15428
rect 14108 15388 14280 15416
rect 14274 15376 14280 15388
rect 14332 15376 14338 15428
rect 15930 15376 15936 15428
rect 15988 15416 15994 15428
rect 16206 15416 16212 15428
rect 15988 15388 16212 15416
rect 15988 15376 15994 15388
rect 16206 15376 16212 15388
rect 16264 15416 16270 15428
rect 17144 15416 17172 15592
rect 18049 15555 18107 15561
rect 18049 15521 18061 15555
rect 18095 15552 18107 15555
rect 18414 15552 18420 15564
rect 18095 15524 18420 15552
rect 18095 15521 18107 15524
rect 18049 15515 18107 15521
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15484 18383 15487
rect 18524 15484 18552 15592
rect 31297 15589 31309 15623
rect 31343 15620 31355 15623
rect 31938 15620 31944 15632
rect 31343 15592 31944 15620
rect 31343 15589 31355 15592
rect 31297 15583 31355 15589
rect 31938 15580 31944 15592
rect 31996 15580 32002 15632
rect 32030 15580 32036 15632
rect 32088 15620 32094 15632
rect 32585 15623 32643 15629
rect 32585 15620 32597 15623
rect 32088 15592 32597 15620
rect 32088 15580 32094 15592
rect 32585 15589 32597 15592
rect 32631 15589 32643 15623
rect 32585 15583 32643 15589
rect 18782 15512 18788 15564
rect 18840 15512 18846 15564
rect 20165 15555 20223 15561
rect 20165 15521 20177 15555
rect 20211 15552 20223 15555
rect 20714 15552 20720 15564
rect 20211 15524 20720 15552
rect 20211 15521 20223 15524
rect 20165 15515 20223 15521
rect 20180 15484 20208 15515
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 20864 15524 21404 15552
rect 20864 15512 20870 15524
rect 18371 15456 20208 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 16264 15388 17172 15416
rect 16264 15376 16270 15388
rect 17310 15376 17316 15428
rect 17368 15416 17374 15428
rect 17681 15419 17739 15425
rect 17681 15416 17693 15419
rect 17368 15388 17693 15416
rect 17368 15376 17374 15388
rect 17681 15385 17693 15388
rect 17727 15385 17739 15419
rect 17681 15379 17739 15385
rect 3326 15308 3332 15360
rect 3384 15348 3390 15360
rect 3694 15348 3700 15360
rect 3384 15320 3700 15348
rect 3384 15308 3390 15320
rect 3694 15308 3700 15320
rect 3752 15348 3758 15360
rect 3973 15351 4031 15357
rect 3973 15348 3985 15351
rect 3752 15320 3985 15348
rect 3752 15308 3758 15320
rect 3973 15317 3985 15320
rect 4019 15317 4031 15351
rect 3973 15311 4031 15317
rect 4062 15308 4068 15360
rect 4120 15348 4126 15360
rect 4157 15351 4215 15357
rect 4157 15348 4169 15351
rect 4120 15320 4169 15348
rect 4120 15308 4126 15320
rect 4157 15317 4169 15320
rect 4203 15317 4215 15351
rect 4157 15311 4215 15317
rect 7282 15308 7288 15360
rect 7340 15348 7346 15360
rect 8018 15348 8024 15360
rect 7340 15320 8024 15348
rect 7340 15308 7346 15320
rect 8018 15308 8024 15320
rect 8076 15308 8082 15360
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 8665 15351 8723 15357
rect 8665 15348 8677 15351
rect 8536 15320 8677 15348
rect 8536 15308 8542 15320
rect 8665 15317 8677 15320
rect 8711 15317 8723 15351
rect 8665 15311 8723 15317
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 9214 15348 9220 15360
rect 9171 15320 9220 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9214 15308 9220 15320
rect 9272 15308 9278 15360
rect 9674 15308 9680 15360
rect 9732 15308 9738 15360
rect 10134 15308 10140 15360
rect 10192 15308 10198 15360
rect 10594 15308 10600 15360
rect 10652 15348 10658 15360
rect 12345 15351 12403 15357
rect 12345 15348 12357 15351
rect 10652 15320 12357 15348
rect 10652 15308 10658 15320
rect 12345 15317 12357 15320
rect 12391 15317 12403 15351
rect 17696 15348 17724 15379
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 18156 15416 18184 15447
rect 20622 15444 20628 15496
rect 20680 15444 20686 15496
rect 20732 15484 20760 15512
rect 21376 15493 21404 15524
rect 23106 15512 23112 15564
rect 23164 15552 23170 15564
rect 23164 15524 23336 15552
rect 23164 15512 23170 15524
rect 21177 15487 21235 15493
rect 21177 15484 21189 15487
rect 20732 15456 21189 15484
rect 21177 15453 21189 15456
rect 21223 15453 21235 15487
rect 21177 15447 21235 15453
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 18012 15388 18184 15416
rect 18012 15376 18018 15388
rect 20714 15376 20720 15428
rect 20772 15376 20778 15428
rect 21192 15416 21220 15447
rect 21450 15444 21456 15496
rect 21508 15444 21514 15496
rect 21818 15444 21824 15496
rect 21876 15444 21882 15496
rect 23308 15484 23336 15524
rect 24394 15512 24400 15564
rect 24452 15512 24458 15564
rect 25133 15555 25191 15561
rect 25133 15521 25145 15555
rect 25179 15552 25191 15555
rect 25498 15552 25504 15564
rect 25179 15524 25504 15552
rect 25179 15521 25191 15524
rect 25133 15515 25191 15521
rect 25498 15512 25504 15524
rect 25556 15512 25562 15564
rect 27890 15512 27896 15564
rect 27948 15552 27954 15564
rect 28169 15555 28227 15561
rect 28169 15552 28181 15555
rect 27948 15524 28181 15552
rect 27948 15512 27954 15524
rect 28169 15521 28181 15524
rect 28215 15521 28227 15555
rect 28169 15515 28227 15521
rect 28718 15512 28724 15564
rect 28776 15552 28782 15564
rect 28776 15524 28948 15552
rect 28776 15512 28782 15524
rect 24857 15487 24915 15493
rect 24857 15484 24869 15487
rect 23308 15456 24869 15484
rect 24857 15453 24869 15456
rect 24903 15453 24915 15487
rect 24857 15447 24915 15453
rect 21192 15388 22048 15416
rect 21910 15348 21916 15360
rect 17696 15320 21916 15348
rect 12345 15311 12403 15317
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 22020 15348 22048 15388
rect 22094 15376 22100 15428
rect 22152 15376 22158 15428
rect 23842 15416 23848 15428
rect 23322 15388 23848 15416
rect 23842 15376 23848 15388
rect 23900 15376 23906 15428
rect 24872 15416 24900 15447
rect 25038 15444 25044 15496
rect 25096 15444 25102 15496
rect 27985 15487 28043 15493
rect 27985 15453 27997 15487
rect 28031 15484 28043 15487
rect 28810 15484 28816 15496
rect 28031 15456 28816 15484
rect 28031 15453 28043 15456
rect 27985 15447 28043 15453
rect 28810 15444 28816 15456
rect 28868 15444 28874 15496
rect 28920 15484 28948 15524
rect 28994 15512 29000 15564
rect 29052 15552 29058 15564
rect 29549 15555 29607 15561
rect 29549 15552 29561 15555
rect 29052 15524 29561 15552
rect 29052 15512 29058 15524
rect 29549 15521 29561 15524
rect 29595 15521 29607 15555
rect 29549 15515 29607 15521
rect 29825 15555 29883 15561
rect 29825 15521 29837 15555
rect 29871 15552 29883 15555
rect 32214 15552 32220 15564
rect 29871 15524 32220 15552
rect 29871 15521 29883 15524
rect 29825 15515 29883 15521
rect 32214 15512 32220 15524
rect 32272 15512 32278 15564
rect 33045 15555 33103 15561
rect 33045 15521 33057 15555
rect 33091 15552 33103 15555
rect 33502 15552 33508 15564
rect 33091 15524 33508 15552
rect 33091 15521 33103 15524
rect 33045 15515 33103 15521
rect 33502 15512 33508 15524
rect 33560 15512 33566 15564
rect 31849 15487 31907 15493
rect 28920 15456 29316 15484
rect 27062 15416 27068 15428
rect 24872 15388 27068 15416
rect 27062 15376 27068 15388
rect 27120 15376 27126 15428
rect 28997 15419 29055 15425
rect 28997 15385 29009 15419
rect 29043 15416 29055 15419
rect 29086 15416 29092 15428
rect 29043 15388 29092 15416
rect 29043 15385 29055 15388
rect 28997 15379 29055 15385
rect 29086 15376 29092 15388
rect 29144 15376 29150 15428
rect 29288 15425 29316 15456
rect 31849 15453 31861 15487
rect 31895 15453 31907 15487
rect 31849 15447 31907 15453
rect 29273 15419 29331 15425
rect 29273 15385 29285 15419
rect 29319 15416 29331 15419
rect 29319 15388 29684 15416
rect 29319 15385 29331 15388
rect 29273 15379 29331 15385
rect 22278 15348 22284 15360
rect 22020 15320 22284 15348
rect 22278 15308 22284 15320
rect 22336 15308 22342 15360
rect 27614 15308 27620 15360
rect 27672 15308 27678 15360
rect 28074 15308 28080 15360
rect 28132 15308 28138 15360
rect 29181 15351 29239 15357
rect 29181 15317 29193 15351
rect 29227 15348 29239 15351
rect 29546 15348 29552 15360
rect 29227 15320 29552 15348
rect 29227 15317 29239 15320
rect 29181 15311 29239 15317
rect 29546 15308 29552 15320
rect 29604 15308 29610 15360
rect 29656 15348 29684 15388
rect 30558 15376 30564 15428
rect 30616 15376 30622 15428
rect 31386 15376 31392 15428
rect 31444 15376 31450 15428
rect 30466 15348 30472 15360
rect 29656 15320 30472 15348
rect 30466 15308 30472 15320
rect 30524 15308 30530 15360
rect 30834 15308 30840 15360
rect 30892 15348 30898 15360
rect 31570 15348 31576 15360
rect 30892 15320 31576 15348
rect 30892 15308 30898 15320
rect 31570 15308 31576 15320
rect 31628 15348 31634 15360
rect 31864 15348 31892 15447
rect 31938 15444 31944 15496
rect 31996 15484 32002 15496
rect 32033 15487 32091 15493
rect 32033 15484 32045 15487
rect 31996 15456 32045 15484
rect 31996 15444 32002 15456
rect 32033 15453 32045 15456
rect 32079 15453 32091 15487
rect 32033 15447 32091 15453
rect 32122 15444 32128 15496
rect 32180 15444 32186 15496
rect 33137 15487 33195 15493
rect 33137 15453 33149 15487
rect 33183 15484 33195 15487
rect 33410 15484 33416 15496
rect 33183 15456 33416 15484
rect 33183 15453 33195 15456
rect 33137 15447 33195 15453
rect 33410 15444 33416 15456
rect 33468 15444 33474 15496
rect 32140 15416 32168 15444
rect 33045 15419 33103 15425
rect 33045 15416 33057 15419
rect 32140 15388 33057 15416
rect 33045 15385 33057 15388
rect 33091 15385 33103 15419
rect 33045 15379 33103 15385
rect 34514 15348 34520 15360
rect 31628 15320 34520 15348
rect 31628 15308 31634 15320
rect 34514 15308 34520 15320
rect 34572 15308 34578 15360
rect 1104 15258 37076 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 37076 15258
rect 1104 15184 37076 15206
rect 3510 15104 3516 15156
rect 3568 15104 3574 15156
rect 7282 15104 7288 15156
rect 7340 15104 7346 15156
rect 7650 15104 7656 15156
rect 7708 15104 7714 15156
rect 7742 15104 7748 15156
rect 7800 15104 7806 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 10376 15116 10916 15144
rect 10376 15104 10382 15116
rect 3142 15036 3148 15088
rect 3200 15036 3206 15088
rect 3234 15036 3240 15088
rect 3292 15076 3298 15088
rect 3345 15079 3403 15085
rect 3345 15076 3357 15079
rect 3292 15048 3357 15076
rect 3292 15036 3298 15048
rect 3345 15045 3357 15048
rect 3391 15076 3403 15079
rect 4062 15076 4068 15088
rect 3391 15048 4068 15076
rect 3391 15045 3403 15048
rect 3345 15039 3403 15045
rect 4062 15036 4068 15048
rect 4120 15076 4126 15088
rect 4120 15048 5672 15076
rect 4120 15036 4126 15048
rect 5261 15011 5319 15017
rect 5261 14977 5273 15011
rect 5307 15008 5319 15011
rect 5537 15011 5595 15017
rect 5537 15008 5549 15011
rect 5307 14980 5549 15008
rect 5307 14977 5319 14980
rect 5261 14971 5319 14977
rect 5537 14977 5549 14980
rect 5583 14977 5595 15011
rect 5644 15008 5672 15048
rect 5718 15036 5724 15088
rect 5776 15036 5782 15088
rect 5920 15048 6868 15076
rect 5920 15017 5948 15048
rect 6196 15017 6224 15048
rect 5905 15011 5963 15017
rect 5905 15008 5917 15011
rect 5644 14980 5917 15008
rect 5537 14971 5595 14977
rect 5905 14977 5917 14980
rect 5951 14977 5963 15011
rect 6181 15011 6239 15017
rect 5905 14971 5963 14977
rect 5997 15001 6055 15007
rect 5997 14967 6009 15001
rect 6043 14967 6055 15001
rect 6181 14977 6193 15011
rect 6227 14977 6239 15011
rect 6840 15008 6868 15048
rect 7300 15008 7328 15104
rect 7377 15079 7435 15085
rect 7377 15045 7389 15079
rect 7423 15076 7435 15079
rect 7926 15076 7932 15088
rect 7423 15048 7932 15076
rect 7423 15045 7435 15048
rect 7377 15039 7435 15045
rect 7926 15036 7932 15048
rect 7984 15036 7990 15088
rect 10134 15036 10140 15088
rect 10192 15076 10198 15088
rect 10192 15048 10824 15076
rect 10192 15036 10198 15048
rect 6840 14980 7328 15008
rect 7469 15011 7527 15017
rect 6181 14971 6239 14977
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7515 14980 8217 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 8205 14977 8217 14980
rect 8251 15008 8263 15011
rect 8478 15008 8484 15020
rect 8251 14980 8484 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 5997 14961 6055 14967
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14940 5503 14943
rect 5491 14912 5672 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 5644 14816 5672 14912
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 6012 14872 6040 14961
rect 7926 14900 7932 14952
rect 7984 14900 7990 14952
rect 8018 14900 8024 14952
rect 8076 14900 8082 14952
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14909 8171 14943
rect 8113 14903 8171 14909
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 6730 14872 6736 14884
rect 5776 14844 6736 14872
rect 5776 14832 5782 14844
rect 6730 14832 6736 14844
rect 6788 14872 6794 14884
rect 7101 14875 7159 14881
rect 7101 14872 7113 14875
rect 6788 14844 7113 14872
rect 6788 14832 6794 14844
rect 7101 14841 7113 14844
rect 7147 14872 7159 14875
rect 7147 14844 7788 14872
rect 7147 14841 7159 14844
rect 7101 14835 7159 14841
rect 3326 14764 3332 14816
rect 3384 14764 3390 14816
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5258 14804 5264 14816
rect 5123 14776 5264 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 6089 14807 6147 14813
rect 6089 14804 6101 14807
rect 5684 14776 6101 14804
rect 5684 14764 5690 14776
rect 6089 14773 6101 14776
rect 6135 14773 6147 14807
rect 7760 14804 7788 14844
rect 8128 14804 8156 14903
rect 7760 14776 8156 14804
rect 8588 14804 8616 14903
rect 8846 14900 8852 14952
rect 8904 14900 8910 14952
rect 9968 14872 9996 14994
rect 10594 14968 10600 15020
rect 10652 14968 10658 15020
rect 10796 14952 10824 15048
rect 10888 15017 10916 15116
rect 11054 15104 11060 15156
rect 11112 15104 11118 15156
rect 19058 15144 19064 15156
rect 15488 15116 19064 15144
rect 15488 15017 15516 15116
rect 19058 15104 19064 15116
rect 19116 15104 19122 15156
rect 20714 15144 20720 15156
rect 19168 15116 20116 15144
rect 19168 15076 19196 15116
rect 18170 15048 19196 15076
rect 19978 15036 19984 15088
rect 20036 15076 20042 15088
rect 20088 15076 20116 15116
rect 20456 15116 20720 15144
rect 20456 15085 20484 15116
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22152 15116 22937 15144
rect 22152 15104 22158 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 22925 15107 22983 15113
rect 23290 15104 23296 15156
rect 23348 15104 23354 15156
rect 27724 15116 28672 15144
rect 20036 15048 20116 15076
rect 20441 15079 20499 15085
rect 20036 15036 20042 15048
rect 20441 15045 20453 15079
rect 20487 15045 20499 15079
rect 21818 15076 21824 15088
rect 20441 15039 20499 15045
rect 20732 15048 21824 15076
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 20732 15017 20760 15048
rect 21818 15036 21824 15048
rect 21876 15076 21882 15088
rect 22741 15079 22799 15085
rect 22741 15076 22753 15079
rect 21876 15048 22753 15076
rect 21876 15036 21882 15048
rect 22741 15045 22753 15048
rect 22787 15076 22799 15079
rect 23750 15076 23756 15088
rect 22787 15048 23756 15076
rect 22787 15045 22799 15048
rect 22741 15039 22799 15045
rect 23750 15036 23756 15048
rect 23808 15076 23814 15088
rect 24394 15076 24400 15088
rect 23808 15048 24400 15076
rect 23808 15036 23814 15048
rect 24394 15036 24400 15048
rect 24452 15036 24458 15088
rect 25961 15079 26019 15085
rect 25961 15045 25973 15079
rect 26007 15076 26019 15079
rect 26142 15076 26148 15088
rect 26007 15048 26148 15076
rect 26007 15045 26019 15048
rect 25961 15039 26019 15045
rect 26142 15036 26148 15048
rect 26200 15036 26206 15088
rect 27341 15079 27399 15085
rect 27341 15045 27353 15079
rect 27387 15076 27399 15079
rect 27614 15076 27620 15088
rect 27387 15048 27620 15076
rect 27387 15045 27399 15048
rect 27341 15039 27399 15045
rect 27614 15036 27620 15048
rect 27672 15036 27678 15088
rect 27724 15076 27752 15116
rect 27798 15076 27804 15088
rect 27724 15048 27804 15076
rect 27798 15036 27804 15048
rect 27856 15036 27862 15088
rect 28644 15076 28672 15116
rect 28810 15104 28816 15156
rect 28868 15104 28874 15156
rect 30193 15147 30251 15153
rect 30193 15113 30205 15147
rect 30239 15144 30251 15147
rect 30466 15144 30472 15156
rect 30239 15116 30472 15144
rect 30239 15113 30251 15116
rect 30193 15107 30251 15113
rect 30466 15104 30472 15116
rect 30524 15144 30530 15156
rect 32766 15144 32772 15156
rect 30524 15116 32772 15144
rect 30524 15104 30530 15116
rect 32766 15104 32772 15116
rect 32824 15144 32830 15156
rect 34606 15144 34612 15156
rect 32824 15116 34612 15144
rect 32824 15104 32830 15116
rect 34606 15104 34612 15116
rect 34664 15104 34670 15156
rect 30650 15076 30656 15088
rect 28644 15048 30656 15076
rect 30650 15036 30656 15048
rect 30708 15036 30714 15088
rect 33594 15036 33600 15088
rect 33652 15036 33658 15088
rect 34164 15048 35190 15076
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 21910 14968 21916 15020
rect 21968 14968 21974 15020
rect 26053 15011 26111 15017
rect 26053 14977 26065 15011
rect 26099 15008 26111 15011
rect 26326 15008 26332 15020
rect 26099 14980 26332 15008
rect 26099 14977 26111 14980
rect 26053 14971 26111 14977
rect 26326 14968 26332 14980
rect 26384 14968 26390 15020
rect 31294 14968 31300 15020
rect 31352 15008 31358 15020
rect 31481 15011 31539 15017
rect 31481 15008 31493 15011
rect 31352 14980 31493 15008
rect 31352 14968 31358 14980
rect 31481 14977 31493 14980
rect 31527 14977 31539 15011
rect 31481 14971 31539 14977
rect 10042 14900 10048 14952
rect 10100 14940 10106 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 10100 14912 10333 14940
rect 10100 14900 10106 14912
rect 10321 14909 10333 14912
rect 10367 14940 10379 14943
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 10367 14912 10701 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 10778 14900 10784 14952
rect 10836 14900 10842 14952
rect 15013 14943 15071 14949
rect 15013 14909 15025 14943
rect 15059 14940 15071 14943
rect 15562 14940 15568 14952
rect 15059 14912 15568 14940
rect 15059 14909 15071 14912
rect 15013 14903 15071 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 15746 14900 15752 14952
rect 15804 14900 15810 14952
rect 16666 14900 16672 14952
rect 16724 14900 16730 14952
rect 16945 14943 17003 14949
rect 16945 14909 16957 14943
rect 16991 14940 17003 14943
rect 17586 14940 17592 14952
rect 16991 14912 17592 14940
rect 16991 14909 17003 14912
rect 16945 14903 17003 14909
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14940 19027 14943
rect 21450 14940 21456 14952
rect 19015 14912 21456 14940
rect 19015 14909 19027 14912
rect 18969 14903 19027 14909
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 23385 14943 23443 14949
rect 23385 14909 23397 14943
rect 23431 14909 23443 14943
rect 23385 14903 23443 14909
rect 23569 14943 23627 14949
rect 23569 14909 23581 14943
rect 23615 14940 23627 14943
rect 23658 14940 23664 14952
rect 23615 14912 23664 14940
rect 23615 14909 23627 14912
rect 23569 14903 23627 14909
rect 11330 14872 11336 14884
rect 9968 14844 11336 14872
rect 11330 14832 11336 14844
rect 11388 14832 11394 14884
rect 23400 14872 23428 14903
rect 23658 14900 23664 14912
rect 23716 14900 23722 14952
rect 25958 14900 25964 14952
rect 26016 14900 26022 14952
rect 26234 14900 26240 14952
rect 26292 14940 26298 14952
rect 27065 14943 27123 14949
rect 27065 14940 27077 14943
rect 26292 14912 27077 14940
rect 26292 14900 26298 14912
rect 27065 14909 27077 14912
rect 27111 14909 27123 14943
rect 30834 14940 30840 14952
rect 27065 14903 27123 14909
rect 27172 14912 30840 14940
rect 23934 14872 23940 14884
rect 23400 14844 23940 14872
rect 23934 14832 23940 14844
rect 23992 14832 23998 14884
rect 24854 14832 24860 14884
rect 24912 14872 24918 14884
rect 27172 14872 27200 14912
rect 30834 14900 30840 14912
rect 30892 14900 30898 14952
rect 32585 14943 32643 14949
rect 32585 14909 32597 14943
rect 32631 14909 32643 14943
rect 32585 14903 32643 14909
rect 24912 14844 27200 14872
rect 24912 14832 24918 14844
rect 9858 14804 9864 14816
rect 8588 14776 9864 14804
rect 6089 14767 6147 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18417 14807 18475 14813
rect 18417 14804 18429 14807
rect 18012 14776 18429 14804
rect 18012 14764 18018 14776
rect 18417 14773 18429 14776
rect 18463 14773 18475 14807
rect 18417 14767 18475 14773
rect 25498 14764 25504 14816
rect 25556 14764 25562 14816
rect 31754 14764 31760 14816
rect 31812 14804 31818 14816
rect 32600 14804 32628 14903
rect 32858 14900 32864 14952
rect 32916 14900 32922 14952
rect 33594 14900 33600 14952
rect 33652 14940 33658 14952
rect 34164 14940 34192 15048
rect 33652 14912 34192 14940
rect 33652 14900 33658 14912
rect 34422 14900 34428 14952
rect 34480 14900 34486 14952
rect 34698 14900 34704 14952
rect 34756 14900 34762 14952
rect 34440 14872 34468 14900
rect 33888 14844 34468 14872
rect 33888 14804 33916 14844
rect 31812 14776 33916 14804
rect 31812 14764 31818 14776
rect 34330 14764 34336 14816
rect 34388 14764 34394 14816
rect 35434 14764 35440 14816
rect 35492 14804 35498 14816
rect 36173 14807 36231 14813
rect 36173 14804 36185 14807
rect 35492 14776 36185 14804
rect 35492 14764 35498 14776
rect 36173 14773 36185 14776
rect 36219 14773 36231 14807
rect 36173 14767 36231 14773
rect 1104 14714 37076 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 37076 14714
rect 1104 14640 37076 14662
rect 6730 14560 6736 14612
rect 6788 14560 6794 14612
rect 10778 14600 10784 14612
rect 9416 14572 10784 14600
rect 3421 14535 3479 14541
rect 3421 14501 3433 14535
rect 3467 14501 3479 14535
rect 3421 14495 3479 14501
rect 1670 14424 1676 14476
rect 1728 14424 1734 14476
rect 1854 14424 1860 14476
rect 1912 14464 1918 14476
rect 1949 14467 2007 14473
rect 1949 14464 1961 14467
rect 1912 14436 1961 14464
rect 1912 14424 1918 14436
rect 1949 14433 1961 14436
rect 1995 14433 2007 14467
rect 3436 14464 3464 14495
rect 3436 14436 4016 14464
rect 1949 14427 2007 14433
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14365 1639 14399
rect 1688 14396 1716 14424
rect 3145 14399 3203 14405
rect 3145 14396 3157 14399
rect 1688 14368 3157 14396
rect 1581 14359 1639 14365
rect 3145 14365 3157 14368
rect 3191 14396 3203 14399
rect 3234 14396 3240 14408
rect 3191 14368 3240 14396
rect 3191 14365 3203 14368
rect 3145 14359 3203 14365
rect 1596 14260 1624 14359
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3510 14356 3516 14408
rect 3568 14396 3574 14408
rect 3988 14405 4016 14436
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 4985 14467 5043 14473
rect 4985 14464 4997 14467
rect 4672 14436 4997 14464
rect 4672 14424 4678 14436
rect 4985 14433 4997 14436
rect 5031 14433 5043 14467
rect 4985 14427 5043 14433
rect 5258 14424 5264 14476
rect 5316 14424 5322 14476
rect 9416 14405 9444 14572
rect 10778 14560 10784 14572
rect 10836 14600 10842 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 10836 14572 11621 14600
rect 10836 14560 10842 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 11609 14563 11667 14569
rect 14093 14603 14151 14609
rect 14093 14569 14105 14603
rect 14139 14600 14151 14603
rect 15746 14600 15752 14612
rect 14139 14572 15752 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 23934 14560 23940 14612
rect 23992 14560 23998 14612
rect 27985 14603 28043 14609
rect 27985 14569 27997 14603
rect 28031 14600 28043 14603
rect 28074 14600 28080 14612
rect 28031 14572 28080 14600
rect 28031 14569 28043 14572
rect 27985 14563 28043 14569
rect 28074 14560 28080 14572
rect 28132 14560 28138 14612
rect 29917 14603 29975 14609
rect 29917 14569 29929 14603
rect 29963 14600 29975 14603
rect 32122 14600 32128 14612
rect 29963 14572 32128 14600
rect 29963 14569 29975 14572
rect 29917 14563 29975 14569
rect 32122 14560 32128 14572
rect 32180 14560 32186 14612
rect 33502 14560 33508 14612
rect 33560 14560 33566 14612
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14464 9551 14467
rect 9674 14464 9680 14476
rect 9539 14436 9680 14464
rect 9539 14433 9551 14436
rect 9493 14427 9551 14433
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 9858 14424 9864 14476
rect 9916 14424 9922 14476
rect 11330 14424 11336 14476
rect 11388 14424 11394 14476
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 15841 14467 15899 14473
rect 15841 14464 15853 14467
rect 14332 14436 15853 14464
rect 14332 14424 14338 14436
rect 15841 14433 15853 14436
rect 15887 14464 15899 14467
rect 16666 14464 16672 14476
rect 15887 14436 16672 14464
rect 15887 14433 15899 14436
rect 15841 14427 15899 14433
rect 16666 14424 16672 14436
rect 16724 14464 16730 14476
rect 18598 14464 18604 14476
rect 16724 14436 18604 14464
rect 16724 14424 16730 14436
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 21818 14424 21824 14476
rect 21876 14464 21882 14476
rect 22189 14467 22247 14473
rect 22189 14464 22201 14467
rect 21876 14436 22201 14464
rect 21876 14424 21882 14436
rect 22189 14433 22201 14436
rect 22235 14433 22247 14467
rect 22189 14427 22247 14433
rect 24394 14424 24400 14476
rect 24452 14424 24458 14476
rect 31386 14424 31392 14476
rect 31444 14424 31450 14476
rect 31665 14467 31723 14473
rect 31665 14433 31677 14467
rect 31711 14464 31723 14467
rect 31754 14464 31760 14476
rect 31711 14436 31760 14464
rect 31711 14433 31723 14436
rect 31665 14427 31723 14433
rect 31754 14424 31760 14436
rect 31812 14424 31818 14476
rect 32030 14424 32036 14476
rect 32088 14424 32094 14476
rect 34698 14424 34704 14476
rect 34756 14424 34762 14476
rect 35434 14424 35440 14476
rect 35492 14424 35498 14476
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3568 14368 3801 14396
rect 3568 14356 3574 14368
rect 3789 14365 3801 14368
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14365 9459 14399
rect 9876 14396 9904 14424
rect 11348 14396 11376 14424
rect 9401 14359 9459 14365
rect 9508 14368 9904 14396
rect 11270 14368 11376 14396
rect 2958 14288 2964 14340
rect 3016 14328 3022 14340
rect 3326 14328 3332 14340
rect 3016 14300 3332 14328
rect 3016 14288 3022 14300
rect 3326 14288 3332 14300
rect 3384 14328 3390 14340
rect 3421 14331 3479 14337
rect 3421 14328 3433 14331
rect 3384 14300 3433 14328
rect 3384 14288 3390 14300
rect 3421 14297 3433 14300
rect 3467 14297 3479 14331
rect 3421 14291 3479 14297
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 5592 14300 5750 14328
rect 5592 14288 5598 14300
rect 6914 14288 6920 14340
rect 6972 14328 6978 14340
rect 9508 14328 9536 14368
rect 26234 14356 26240 14408
rect 26292 14356 26298 14408
rect 34514 14356 34520 14408
rect 34572 14396 34578 14408
rect 35161 14399 35219 14405
rect 35161 14396 35173 14399
rect 34572 14368 35173 14396
rect 34572 14356 34578 14368
rect 35161 14365 35173 14368
rect 35207 14365 35219 14399
rect 35161 14359 35219 14365
rect 35345 14399 35403 14405
rect 35345 14365 35357 14399
rect 35391 14365 35403 14399
rect 35345 14359 35403 14365
rect 10137 14331 10195 14337
rect 10137 14328 10149 14331
rect 6972 14300 9536 14328
rect 9784 14300 10149 14328
rect 6972 14288 6978 14300
rect 3142 14260 3148 14272
rect 1596 14232 3148 14260
rect 3142 14220 3148 14232
rect 3200 14260 3206 14272
rect 3237 14263 3295 14269
rect 3237 14260 3249 14263
rect 3200 14232 3249 14260
rect 3200 14220 3206 14232
rect 3237 14229 3249 14232
rect 3283 14229 3295 14263
rect 3237 14223 3295 14229
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 4430 14260 4436 14272
rect 3927 14232 4436 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 9784 14269 9812 14300
rect 10137 14297 10149 14300
rect 10183 14297 10195 14331
rect 15470 14328 15476 14340
rect 15134 14300 15476 14328
rect 10137 14291 10195 14297
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 15562 14288 15568 14340
rect 15620 14288 15626 14340
rect 18325 14331 18383 14337
rect 16546 14300 17158 14328
rect 9769 14263 9827 14269
rect 9769 14229 9781 14263
rect 9815 14229 9827 14263
rect 15488 14260 15516 14288
rect 16390 14260 16396 14272
rect 15488 14232 16396 14260
rect 9769 14223 9827 14229
rect 16390 14220 16396 14232
rect 16448 14260 16454 14272
rect 16546 14260 16574 14300
rect 18325 14297 18337 14331
rect 18371 14328 18383 14331
rect 18414 14328 18420 14340
rect 18371 14300 18420 14328
rect 18371 14297 18383 14300
rect 18325 14291 18383 14297
rect 18414 14288 18420 14300
rect 18472 14288 18478 14340
rect 20349 14331 20407 14337
rect 20349 14297 20361 14331
rect 20395 14328 20407 14331
rect 20622 14328 20628 14340
rect 20395 14300 20628 14328
rect 20395 14297 20407 14300
rect 20349 14291 20407 14297
rect 20622 14288 20628 14300
rect 20680 14328 20686 14340
rect 21266 14328 21272 14340
rect 20680 14300 21272 14328
rect 20680 14288 20686 14300
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 22465 14331 22523 14337
rect 22465 14297 22477 14331
rect 22511 14328 22523 14331
rect 22738 14328 22744 14340
rect 22511 14300 22744 14328
rect 22511 14297 22523 14300
rect 22465 14291 22523 14297
rect 22738 14288 22744 14300
rect 22796 14288 22802 14340
rect 23842 14328 23848 14340
rect 23690 14300 23848 14328
rect 23842 14288 23848 14300
rect 23900 14328 23906 14340
rect 23900 14300 24624 14328
rect 23900 14288 23906 14300
rect 16448 14232 16574 14260
rect 16853 14263 16911 14269
rect 16448 14220 16454 14232
rect 16853 14229 16865 14263
rect 16899 14260 16911 14263
rect 18046 14260 18052 14272
rect 16899 14232 18052 14260
rect 16899 14229 16911 14232
rect 16853 14223 16911 14229
rect 18046 14220 18052 14232
rect 18104 14220 18110 14272
rect 21634 14220 21640 14272
rect 21692 14260 21698 14272
rect 21821 14263 21879 14269
rect 21821 14260 21833 14263
rect 21692 14232 21833 14260
rect 21692 14220 21698 14232
rect 21821 14229 21833 14232
rect 21867 14260 21879 14263
rect 22830 14260 22836 14272
rect 21867 14232 22836 14260
rect 21867 14229 21879 14232
rect 21821 14223 21879 14229
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 24596 14260 24624 14300
rect 24670 14288 24676 14340
rect 24728 14288 24734 14340
rect 25898 14300 26372 14328
rect 25976 14260 26004 14300
rect 26344 14272 26372 14300
rect 26510 14288 26516 14340
rect 26568 14288 26574 14340
rect 27798 14328 27804 14340
rect 27738 14300 27804 14328
rect 27798 14288 27804 14300
rect 27856 14288 27862 14340
rect 30650 14288 30656 14340
rect 30708 14288 30714 14340
rect 33318 14328 33324 14340
rect 33258 14300 33324 14328
rect 33318 14288 33324 14300
rect 33376 14328 33382 14340
rect 33594 14328 33600 14340
rect 33376 14300 33600 14328
rect 33376 14288 33382 14300
rect 33594 14288 33600 14300
rect 33652 14288 33658 14340
rect 34330 14288 34336 14340
rect 34388 14328 34394 14340
rect 35360 14328 35388 14359
rect 34388 14300 35388 14328
rect 34388 14288 34394 14300
rect 24596 14232 26004 14260
rect 26142 14220 26148 14272
rect 26200 14220 26206 14272
rect 26326 14220 26332 14272
rect 26384 14220 26390 14272
rect 1104 14170 37076 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 37076 14170
rect 1104 14096 37076 14118
rect 1302 14016 1308 14068
rect 1360 14056 1366 14068
rect 1397 14059 1455 14065
rect 1397 14056 1409 14059
rect 1360 14028 1409 14056
rect 1360 14016 1366 14028
rect 1397 14025 1409 14028
rect 1443 14025 1455 14059
rect 1397 14019 1455 14025
rect 2958 14016 2964 14068
rect 3016 14016 3022 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5592 14028 7052 14056
rect 5592 14016 5598 14028
rect 3050 13948 3056 14000
rect 3108 13988 3114 14000
rect 3108 13960 3266 13988
rect 3108 13948 3114 13960
rect 4430 13948 4436 14000
rect 4488 13948 4494 14000
rect 6914 13988 6920 14000
rect 6380 13960 6920 13988
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 1670 13920 1676 13932
rect 1627 13892 1676 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 4706 13880 4712 13932
rect 4764 13880 4770 13932
rect 6380 13929 6408 13960
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 7024 13988 7052 14028
rect 17586 14016 17592 14068
rect 17644 14016 17650 14068
rect 17954 14016 17960 14068
rect 18012 14016 18018 14068
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 19613 14059 19671 14065
rect 18104 14028 19196 14056
rect 18104 14016 18110 14028
rect 7024 13960 7130 13988
rect 8846 13948 8852 14000
rect 8904 13988 8910 14000
rect 9033 13991 9091 13997
rect 9033 13988 9045 13991
rect 8904 13960 9045 13988
rect 8904 13948 8910 13960
rect 9033 13957 9045 13960
rect 9079 13957 9091 13991
rect 9033 13951 9091 13957
rect 15562 13948 15568 14000
rect 15620 13948 15626 14000
rect 18414 13948 18420 14000
rect 18472 13948 18478 14000
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 5626 13812 5632 13864
rect 5684 13812 5690 13864
rect 5736 13852 5764 13883
rect 9214 13880 9220 13932
rect 9272 13880 9278 13932
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9674 13920 9680 13932
rect 9447 13892 9680 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13920 18935 13923
rect 18966 13920 18972 13932
rect 18923 13892 18972 13920
rect 18923 13889 18935 13892
rect 18877 13883 18935 13889
rect 18966 13880 18972 13892
rect 19024 13880 19030 13932
rect 19168 13929 19196 14028
rect 19613 14025 19625 14059
rect 19659 14056 19671 14059
rect 19659 14028 21404 14056
rect 19659 14025 19671 14028
rect 19613 14019 19671 14025
rect 21376 13988 21404 14028
rect 21450 14016 21456 14068
rect 21508 14056 21514 14068
rect 26234 14056 26240 14068
rect 21508 14028 22094 14056
rect 21508 14016 21514 14028
rect 22066 13988 22094 14028
rect 24964 14028 26240 14056
rect 21376 13960 21956 13988
rect 22066 13960 22508 13988
rect 19061 13923 19119 13929
rect 19061 13889 19073 13923
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 19153 13923 19211 13929
rect 19153 13889 19165 13923
rect 19199 13889 19211 13923
rect 19153 13883 19211 13889
rect 7926 13852 7932 13864
rect 5736 13824 7932 13852
rect 7926 13812 7932 13824
rect 7984 13852 7990 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 7984 13824 8125 13852
rect 7984 13812 7990 13824
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 8113 13815 8171 13821
rect 14274 13812 14280 13864
rect 14332 13812 14338 13864
rect 14550 13812 14556 13864
rect 14608 13812 14614 13864
rect 18141 13855 18199 13861
rect 18141 13821 18153 13855
rect 18187 13821 18199 13855
rect 18141 13815 18199 13821
rect 18156 13784 18184 13815
rect 18506 13812 18512 13864
rect 18564 13852 18570 13864
rect 19076 13852 19104 13883
rect 19978 13880 19984 13932
rect 20036 13880 20042 13932
rect 21361 13923 21419 13929
rect 21361 13889 21373 13923
rect 21407 13920 21419 13923
rect 21726 13920 21732 13932
rect 21407 13892 21732 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 21726 13880 21732 13892
rect 21784 13880 21790 13932
rect 18564 13824 19104 13852
rect 21085 13855 21143 13861
rect 18564 13812 18570 13824
rect 21085 13821 21097 13855
rect 21131 13852 21143 13855
rect 21821 13855 21879 13861
rect 21821 13852 21833 13855
rect 21131 13824 21833 13852
rect 21131 13821 21143 13824
rect 21085 13815 21143 13821
rect 21821 13821 21833 13824
rect 21867 13821 21879 13855
rect 21928 13852 21956 13960
rect 22002 13880 22008 13932
rect 22060 13920 22066 13932
rect 22480 13929 22508 13960
rect 22738 13948 22744 14000
rect 22796 13988 22802 14000
rect 22925 13991 22983 13997
rect 22925 13988 22937 13991
rect 22796 13960 22937 13988
rect 22796 13948 22802 13960
rect 22925 13957 22937 13960
rect 22971 13957 22983 13991
rect 22925 13951 22983 13957
rect 22281 13923 22339 13929
rect 22281 13920 22293 13923
rect 22060 13892 22293 13920
rect 22060 13880 22066 13892
rect 22281 13889 22293 13892
rect 22327 13889 22339 13923
rect 22281 13883 22339 13889
rect 22465 13923 22523 13929
rect 22465 13889 22477 13923
rect 22511 13889 22523 13923
rect 22465 13883 22523 13889
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13920 23443 13923
rect 23431 13892 23520 13920
rect 23431 13889 23443 13892
rect 23385 13883 23443 13889
rect 22557 13855 22615 13861
rect 22557 13852 22569 13855
rect 21928 13824 22569 13852
rect 21821 13815 21879 13821
rect 22557 13821 22569 13824
rect 22603 13852 22615 13855
rect 23014 13852 23020 13864
rect 22603 13824 23020 13852
rect 22603 13821 22615 13824
rect 22557 13815 22615 13821
rect 23014 13812 23020 13824
rect 23072 13812 23078 13864
rect 23492 13852 23520 13892
rect 23566 13880 23572 13932
rect 23624 13880 23630 13932
rect 23661 13923 23719 13929
rect 23661 13889 23673 13923
rect 23707 13920 23719 13923
rect 23934 13920 23940 13932
rect 23707 13892 23940 13920
rect 23707 13889 23719 13892
rect 23661 13883 23719 13889
rect 23934 13880 23940 13892
rect 23992 13880 23998 13932
rect 24964 13929 24992 14028
rect 26234 14016 26240 14028
rect 26292 14016 26298 14068
rect 26510 14016 26516 14068
rect 26568 14056 26574 14068
rect 26973 14059 27031 14065
rect 26973 14056 26985 14059
rect 26568 14028 26985 14056
rect 26568 14016 26574 14028
rect 26973 14025 26985 14028
rect 27019 14025 27031 14059
rect 26973 14019 27031 14025
rect 27341 14059 27399 14065
rect 27341 14025 27353 14059
rect 27387 14056 27399 14059
rect 28074 14056 28080 14068
rect 27387 14028 28080 14056
rect 27387 14025 27399 14028
rect 27341 14019 27399 14025
rect 28074 14016 28080 14028
rect 28132 14016 28138 14068
rect 31662 14016 31668 14068
rect 31720 14056 31726 14068
rect 32582 14056 32588 14068
rect 31720 14028 32588 14056
rect 31720 14016 31726 14028
rect 32582 14016 32588 14028
rect 32640 14056 32646 14068
rect 32640 14028 33548 14056
rect 32640 14016 32646 14028
rect 25225 13991 25283 13997
rect 25225 13957 25237 13991
rect 25271 13988 25283 13991
rect 25498 13988 25504 14000
rect 25271 13960 25504 13988
rect 25271 13957 25283 13960
rect 25225 13951 25283 13957
rect 25498 13948 25504 13960
rect 25556 13948 25562 14000
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13889 25007 13923
rect 24949 13883 25007 13889
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 26292 13892 26358 13920
rect 26292 13880 26298 13892
rect 29638 13880 29644 13932
rect 29696 13880 29702 13932
rect 29825 13923 29883 13929
rect 29825 13889 29837 13923
rect 29871 13920 29883 13923
rect 31680 13920 31708 14016
rect 32309 13991 32367 13997
rect 32309 13957 32321 13991
rect 32355 13988 32367 13991
rect 32766 13988 32772 14000
rect 32355 13960 32772 13988
rect 32355 13957 32367 13960
rect 32309 13951 32367 13957
rect 32766 13948 32772 13960
rect 32824 13948 32830 14000
rect 32858 13948 32864 14000
rect 32916 13988 32922 14000
rect 33045 13991 33103 13997
rect 33045 13988 33057 13991
rect 32916 13960 33057 13988
rect 32916 13948 32922 13960
rect 33045 13957 33057 13960
rect 33091 13957 33103 13991
rect 33045 13951 33103 13957
rect 29871 13892 31708 13920
rect 29871 13889 29883 13892
rect 29825 13883 29883 13889
rect 32030 13880 32036 13932
rect 32088 13920 32094 13932
rect 32217 13923 32275 13929
rect 32217 13920 32229 13923
rect 32088 13892 32229 13920
rect 32088 13880 32094 13892
rect 32217 13889 32229 13892
rect 32263 13920 32275 13923
rect 33410 13920 33416 13932
rect 32263 13892 33416 13920
rect 32263 13889 32275 13892
rect 32217 13883 32275 13889
rect 33410 13880 33416 13892
rect 33468 13880 33474 13932
rect 33520 13929 33548 14028
rect 33505 13923 33563 13929
rect 33505 13889 33517 13923
rect 33551 13889 33563 13923
rect 33505 13883 33563 13889
rect 33594 13880 33600 13932
rect 33652 13920 33658 13932
rect 33689 13923 33747 13929
rect 33689 13920 33701 13923
rect 33652 13892 33701 13920
rect 33652 13880 33658 13892
rect 33689 13889 33701 13892
rect 33735 13889 33747 13923
rect 33689 13883 33747 13889
rect 33781 13923 33839 13929
rect 33781 13889 33793 13923
rect 33827 13920 33839 13923
rect 34330 13920 34336 13932
rect 33827 13892 34336 13920
rect 33827 13889 33839 13892
rect 33781 13883 33839 13889
rect 34330 13880 34336 13892
rect 34388 13880 34394 13932
rect 24854 13852 24860 13864
rect 23492 13824 24860 13852
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 25958 13812 25964 13864
rect 26016 13852 26022 13864
rect 26697 13855 26755 13861
rect 26697 13852 26709 13855
rect 26016 13824 26709 13852
rect 26016 13812 26022 13824
rect 26697 13821 26709 13824
rect 26743 13852 26755 13855
rect 27433 13855 27491 13861
rect 27433 13852 27445 13855
rect 26743 13824 27445 13852
rect 26743 13821 26755 13824
rect 26697 13815 26755 13821
rect 27433 13821 27445 13824
rect 27479 13821 27491 13855
rect 27433 13815 27491 13821
rect 27617 13855 27675 13861
rect 27617 13821 27629 13855
rect 27663 13821 27675 13855
rect 27617 13815 27675 13821
rect 18230 13784 18236 13796
rect 18156 13756 18236 13784
rect 18230 13744 18236 13756
rect 18288 13744 18294 13796
rect 27632 13784 27660 13815
rect 28902 13812 28908 13864
rect 28960 13812 28966 13864
rect 29181 13855 29239 13861
rect 29181 13821 29193 13855
rect 29227 13852 29239 13855
rect 29270 13852 29276 13864
rect 29227 13824 29276 13852
rect 29227 13821 29239 13824
rect 29181 13815 29239 13821
rect 29270 13812 29276 13824
rect 29328 13812 29334 13864
rect 29546 13812 29552 13864
rect 29604 13812 29610 13864
rect 30282 13812 30288 13864
rect 30340 13812 30346 13864
rect 32398 13812 32404 13864
rect 32456 13812 32462 13864
rect 27890 13784 27896 13796
rect 27632 13756 27896 13784
rect 27890 13744 27896 13756
rect 27948 13744 27954 13796
rect 5997 13719 6055 13725
rect 5997 13685 6009 13719
rect 6043 13716 6055 13719
rect 6622 13719 6680 13725
rect 6622 13716 6634 13719
rect 6043 13688 6634 13716
rect 6043 13685 6055 13688
rect 5997 13679 6055 13685
rect 6622 13685 6634 13688
rect 6668 13685 6680 13719
rect 6622 13679 6680 13685
rect 16022 13676 16028 13728
rect 16080 13676 16086 13728
rect 32769 13719 32827 13725
rect 32769 13685 32781 13719
rect 32815 13716 32827 13719
rect 33870 13716 33876 13728
rect 32815 13688 33876 13716
rect 32815 13685 32827 13688
rect 32769 13679 32827 13685
rect 33870 13676 33876 13688
rect 33928 13676 33934 13728
rect 1104 13626 37076 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 37076 13626
rect 1104 13552 37076 13574
rect 3142 13472 3148 13524
rect 3200 13512 3206 13524
rect 3329 13515 3387 13521
rect 3329 13512 3341 13515
rect 3200 13484 3341 13512
rect 3200 13472 3206 13484
rect 3329 13481 3341 13484
rect 3375 13481 3387 13515
rect 3329 13475 3387 13481
rect 22554 13472 22560 13524
rect 22612 13512 22618 13524
rect 23566 13512 23572 13524
rect 22612 13484 23572 13512
rect 22612 13472 22618 13484
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 32398 13472 32404 13524
rect 32456 13472 32462 13524
rect 28074 13404 28080 13456
rect 28132 13404 28138 13456
rect 1394 13336 1400 13388
rect 1452 13376 1458 13388
rect 1581 13379 1639 13385
rect 1581 13376 1593 13379
rect 1452 13348 1593 13376
rect 1452 13336 1458 13348
rect 1581 13345 1593 13348
rect 1627 13345 1639 13379
rect 1581 13339 1639 13345
rect 1854 13336 1860 13388
rect 1912 13336 1918 13388
rect 3050 13336 3056 13388
rect 3108 13336 3114 13388
rect 14550 13336 14556 13388
rect 14608 13376 14614 13388
rect 15105 13379 15163 13385
rect 15105 13376 15117 13379
rect 14608 13348 15117 13376
rect 14608 13336 14614 13348
rect 15105 13345 15117 13348
rect 15151 13345 15163 13379
rect 15105 13339 15163 13345
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 16022 13376 16028 13388
rect 15887 13348 16028 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 18598 13376 18604 13388
rect 16807 13348 18604 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 18598 13336 18604 13348
rect 18656 13336 18662 13388
rect 20809 13379 20867 13385
rect 20809 13345 20821 13379
rect 20855 13376 20867 13379
rect 21726 13376 21732 13388
rect 20855 13348 21732 13376
rect 20855 13345 20867 13348
rect 20809 13339 20867 13345
rect 21726 13336 21732 13348
rect 21784 13336 21790 13388
rect 24397 13379 24455 13385
rect 24397 13345 24409 13379
rect 24443 13376 24455 13379
rect 24670 13376 24676 13388
rect 24443 13348 24676 13376
rect 24443 13345 24455 13348
rect 24397 13339 24455 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 25133 13379 25191 13385
rect 25133 13345 25145 13379
rect 25179 13376 25191 13379
rect 26142 13376 26148 13388
rect 25179 13348 26148 13376
rect 25179 13345 25191 13348
rect 25133 13339 25191 13345
rect 26142 13336 26148 13348
rect 26200 13336 26206 13388
rect 28629 13379 28687 13385
rect 28629 13345 28641 13379
rect 28675 13376 28687 13379
rect 28902 13376 28908 13388
rect 28675 13348 28908 13376
rect 28675 13345 28687 13348
rect 28629 13339 28687 13345
rect 28902 13336 28908 13348
rect 28960 13336 28966 13388
rect 32309 13379 32367 13385
rect 32309 13345 32321 13379
rect 32355 13376 32367 13379
rect 34149 13379 34207 13385
rect 34149 13376 34161 13379
rect 32355 13348 34161 13376
rect 32355 13345 32367 13348
rect 32309 13339 32367 13345
rect 34149 13345 34161 13348
rect 34195 13376 34207 13379
rect 34422 13376 34428 13388
rect 34195 13348 34428 13376
rect 34195 13345 34207 13348
rect 34149 13339 34207 13345
rect 34422 13336 34428 13348
rect 34480 13336 34486 13388
rect 35253 13379 35311 13385
rect 35253 13345 35265 13379
rect 35299 13376 35311 13379
rect 35342 13376 35348 13388
rect 35299 13348 35348 13376
rect 35299 13345 35311 13348
rect 35253 13339 35311 13345
rect 35342 13336 35348 13348
rect 35400 13336 35406 13388
rect 3068 13308 3096 13336
rect 2990 13280 3096 13308
rect 15562 13268 15568 13320
rect 15620 13268 15626 13320
rect 15746 13268 15752 13320
rect 15804 13268 15810 13320
rect 24854 13268 24860 13320
rect 24912 13268 24918 13320
rect 24946 13268 24952 13320
rect 25004 13308 25010 13320
rect 25041 13311 25099 13317
rect 25041 13308 25053 13311
rect 25004 13280 25053 13308
rect 25004 13268 25010 13280
rect 25041 13277 25053 13280
rect 25087 13277 25099 13311
rect 25041 13271 25099 13277
rect 30098 13268 30104 13320
rect 30156 13308 30162 13320
rect 30650 13308 30656 13320
rect 30156 13280 30656 13308
rect 30156 13268 30162 13280
rect 30650 13268 30656 13280
rect 30708 13308 30714 13320
rect 30708 13294 30958 13308
rect 30708 13280 30972 13294
rect 30708 13268 30714 13280
rect 17034 13200 17040 13252
rect 17092 13200 17098 13252
rect 19978 13240 19984 13252
rect 18262 13212 19984 13240
rect 16390 13132 16396 13184
rect 16448 13172 16454 13184
rect 18340 13172 18368 13212
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 21082 13200 21088 13252
rect 21140 13200 21146 13252
rect 21542 13240 21548 13252
rect 21192 13212 21548 13240
rect 16448 13144 18368 13172
rect 16448 13132 16454 13144
rect 18506 13132 18512 13184
rect 18564 13132 18570 13184
rect 19996 13172 20024 13200
rect 21192 13172 21220 13212
rect 21542 13200 21548 13212
rect 21600 13200 21606 13252
rect 27706 13200 27712 13252
rect 27764 13240 27770 13252
rect 28353 13243 28411 13249
rect 28353 13240 28365 13243
rect 27764 13212 28365 13240
rect 27764 13200 27770 13212
rect 28353 13209 28365 13212
rect 28399 13209 28411 13243
rect 28353 13203 28411 13209
rect 28537 13243 28595 13249
rect 28537 13209 28549 13243
rect 28583 13240 28595 13243
rect 28994 13240 29000 13252
rect 28583 13212 29000 13240
rect 28583 13209 28595 13212
rect 28537 13203 28595 13209
rect 28994 13200 29000 13212
rect 29052 13240 29058 13252
rect 29546 13240 29552 13252
rect 29052 13212 29552 13240
rect 29052 13200 29058 13212
rect 29546 13200 29552 13212
rect 29604 13200 29610 13252
rect 19996 13144 21220 13172
rect 30561 13175 30619 13181
rect 30561 13141 30573 13175
rect 30607 13172 30619 13175
rect 30742 13172 30748 13184
rect 30607 13144 30748 13172
rect 30607 13141 30619 13144
rect 30561 13135 30619 13141
rect 30742 13132 30748 13144
rect 30800 13132 30806 13184
rect 30944 13172 30972 13280
rect 32033 13243 32091 13249
rect 32033 13209 32045 13243
rect 32079 13240 32091 13243
rect 32122 13240 32128 13252
rect 32079 13212 32128 13240
rect 32079 13209 32091 13212
rect 32033 13203 32091 13209
rect 32122 13200 32128 13212
rect 32180 13200 32186 13252
rect 33318 13200 33324 13252
rect 33376 13200 33382 13252
rect 33870 13200 33876 13252
rect 33928 13200 33934 13252
rect 34606 13200 34612 13252
rect 34664 13240 34670 13252
rect 35345 13243 35403 13249
rect 35345 13240 35357 13243
rect 34664 13212 35357 13240
rect 34664 13200 34670 13212
rect 35345 13209 35357 13212
rect 35391 13209 35403 13243
rect 35345 13203 35403 13209
rect 33594 13172 33600 13184
rect 30944 13144 33600 13172
rect 33594 13132 33600 13144
rect 33652 13132 33658 13184
rect 33686 13132 33692 13184
rect 33744 13172 33750 13184
rect 34775 13175 34833 13181
rect 34775 13172 34787 13175
rect 33744 13144 34787 13172
rect 33744 13132 33750 13144
rect 34775 13141 34787 13144
rect 34821 13141 34833 13175
rect 34775 13135 34833 13141
rect 35253 13175 35311 13181
rect 35253 13141 35265 13175
rect 35299 13172 35311 13175
rect 35434 13172 35440 13184
rect 35299 13144 35440 13172
rect 35299 13141 35311 13144
rect 35253 13135 35311 13141
rect 35434 13132 35440 13144
rect 35492 13132 35498 13184
rect 1104 13082 37076 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 37076 13082
rect 1104 13008 37076 13030
rect 22002 12968 22008 12980
rect 18892 12940 22008 12968
rect 16390 12900 16396 12912
rect 15870 12872 16396 12900
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 18892 12900 18920 12940
rect 22002 12928 22008 12940
rect 22060 12928 22066 12980
rect 24596 12940 24900 12968
rect 18432 12872 18920 12900
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 14332 12804 14381 12832
rect 14332 12792 14338 12804
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 14645 12767 14703 12773
rect 14645 12733 14657 12767
rect 14691 12764 14703 12767
rect 15194 12764 15200 12776
rect 14691 12736 15200 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15654 12724 15660 12776
rect 15712 12764 15718 12776
rect 18046 12764 18052 12776
rect 15712 12736 18052 12764
rect 15712 12724 15718 12736
rect 18046 12724 18052 12736
rect 18104 12764 18110 12776
rect 18432 12773 18460 12872
rect 19978 12860 19984 12912
rect 20036 12860 20042 12912
rect 21726 12860 21732 12912
rect 21784 12900 21790 12912
rect 21784 12872 23244 12900
rect 21784 12860 21790 12872
rect 18874 12792 18880 12844
rect 18932 12792 18938 12844
rect 21082 12792 21088 12844
rect 21140 12832 21146 12844
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 21140 12804 21833 12832
rect 21140 12792 21146 12804
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 22278 12792 22284 12844
rect 22336 12792 22342 12844
rect 22465 12835 22523 12841
rect 22465 12801 22477 12835
rect 22511 12801 22523 12835
rect 22465 12795 22523 12801
rect 18417 12767 18475 12773
rect 18417 12764 18429 12767
rect 18104 12736 18429 12764
rect 18104 12724 18110 12736
rect 18417 12733 18429 12736
rect 18463 12733 18475 12767
rect 18417 12727 18475 12733
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 18656 12736 18981 12764
rect 18656 12724 18662 12736
rect 18969 12733 18981 12736
rect 19015 12733 19027 12767
rect 18969 12727 19027 12733
rect 19245 12767 19303 12773
rect 19245 12733 19257 12767
rect 19291 12764 19303 12767
rect 19610 12764 19616 12776
rect 19291 12736 19616 12764
rect 19291 12733 19303 12736
rect 19245 12727 19303 12733
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 20714 12724 20720 12776
rect 20772 12764 20778 12776
rect 22480 12764 22508 12795
rect 22554 12792 22560 12844
rect 22612 12792 22618 12844
rect 23216 12841 23244 12872
rect 24596 12844 24624 12940
rect 24872 12900 24900 12940
rect 24946 12928 24952 12980
rect 25004 12968 25010 12980
rect 25409 12971 25467 12977
rect 25409 12968 25421 12971
rect 25004 12940 25421 12968
rect 25004 12928 25010 12940
rect 25409 12937 25421 12940
rect 25455 12937 25467 12971
rect 25409 12931 25467 12937
rect 28537 12971 28595 12977
rect 28537 12937 28549 12971
rect 28583 12968 28595 12971
rect 28994 12968 29000 12980
rect 28583 12940 29000 12968
rect 28583 12937 28595 12940
rect 28537 12931 28595 12937
rect 28994 12928 29000 12940
rect 29052 12928 29058 12980
rect 29638 12928 29644 12980
rect 29696 12968 29702 12980
rect 34606 12968 34612 12980
rect 29696 12940 30696 12968
rect 29696 12928 29702 12940
rect 26234 12900 26240 12912
rect 24872 12872 26240 12900
rect 26234 12860 26240 12872
rect 26292 12860 26298 12912
rect 29914 12900 29920 12912
rect 29578 12872 29920 12900
rect 29914 12860 29920 12872
rect 29972 12860 29978 12912
rect 30009 12903 30067 12909
rect 30009 12869 30021 12903
rect 30055 12900 30067 12903
rect 30282 12900 30288 12912
rect 30055 12872 30288 12900
rect 30055 12869 30067 12872
rect 30009 12863 30067 12869
rect 30282 12860 30288 12872
rect 30340 12860 30346 12912
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 24578 12792 24584 12844
rect 24636 12792 24642 12844
rect 27338 12792 27344 12844
rect 27396 12792 27402 12844
rect 30668 12841 30696 12940
rect 31726 12940 34612 12968
rect 30653 12835 30711 12841
rect 30653 12801 30665 12835
rect 30699 12801 30711 12835
rect 30653 12795 30711 12801
rect 30742 12792 30748 12844
rect 30800 12792 30806 12844
rect 30929 12835 30987 12841
rect 30929 12801 30941 12835
rect 30975 12832 30987 12835
rect 31110 12832 31116 12844
rect 30975 12804 31116 12832
rect 30975 12801 30987 12804
rect 30929 12795 30987 12801
rect 31110 12792 31116 12804
rect 31168 12832 31174 12844
rect 31726 12832 31754 12940
rect 34606 12928 34612 12940
rect 34664 12928 34670 12980
rect 32122 12860 32128 12912
rect 32180 12860 32186 12912
rect 32398 12860 32404 12912
rect 32456 12900 32462 12912
rect 32456 12872 32812 12900
rect 32456 12860 32462 12872
rect 31168 12804 31754 12832
rect 31168 12792 31174 12804
rect 32582 12792 32588 12844
rect 32640 12792 32646 12844
rect 32784 12841 32812 12872
rect 33686 12860 33692 12912
rect 33744 12860 33750 12912
rect 33778 12860 33784 12912
rect 33836 12900 33842 12912
rect 33836 12872 34178 12900
rect 33836 12860 33842 12872
rect 32769 12835 32827 12841
rect 32769 12801 32781 12835
rect 32815 12801 32827 12835
rect 32769 12795 32827 12801
rect 20772 12736 22508 12764
rect 23477 12767 23535 12773
rect 20772 12724 20778 12736
rect 23477 12733 23489 12767
rect 23523 12764 23535 12767
rect 23523 12736 25084 12764
rect 23523 12733 23535 12736
rect 23477 12727 23535 12733
rect 25056 12705 25084 12736
rect 25498 12724 25504 12776
rect 25556 12724 25562 12776
rect 25685 12767 25743 12773
rect 25685 12733 25697 12767
rect 25731 12733 25743 12767
rect 25685 12727 25743 12733
rect 25041 12699 25099 12705
rect 25041 12665 25053 12699
rect 25087 12665 25099 12699
rect 25700 12696 25728 12727
rect 26970 12724 26976 12776
rect 27028 12764 27034 12776
rect 27433 12767 27491 12773
rect 27433 12764 27445 12767
rect 27028 12736 27445 12764
rect 27028 12724 27034 12736
rect 27433 12733 27445 12736
rect 27479 12733 27491 12767
rect 27433 12727 27491 12733
rect 27525 12767 27583 12773
rect 27525 12733 27537 12767
rect 27571 12733 27583 12767
rect 27525 12727 27583 12733
rect 30285 12767 30343 12773
rect 30285 12733 30297 12767
rect 30331 12764 30343 12767
rect 30558 12764 30564 12776
rect 30331 12736 30564 12764
rect 30331 12733 30343 12736
rect 30285 12727 30343 12733
rect 26050 12696 26056 12708
rect 25700 12668 26056 12696
rect 25041 12659 25099 12665
rect 26050 12656 26056 12668
rect 26108 12696 26114 12708
rect 27540 12696 27568 12727
rect 30558 12724 30564 12736
rect 30616 12724 30622 12776
rect 26108 12668 27568 12696
rect 30760 12696 30788 12792
rect 31018 12724 31024 12776
rect 31076 12764 31082 12776
rect 31389 12767 31447 12773
rect 31389 12764 31401 12767
rect 31076 12736 31401 12764
rect 31076 12724 31082 12736
rect 31389 12733 31401 12736
rect 31435 12733 31447 12767
rect 32861 12767 32919 12773
rect 32861 12764 32873 12767
rect 31389 12727 31447 12733
rect 31726 12736 32873 12764
rect 31726 12696 31754 12736
rect 32861 12733 32873 12736
rect 32907 12733 32919 12767
rect 32861 12727 32919 12733
rect 33042 12724 33048 12776
rect 33100 12764 33106 12776
rect 33413 12767 33471 12773
rect 33413 12764 33425 12767
rect 33100 12736 33425 12764
rect 33100 12724 33106 12736
rect 33413 12733 33425 12736
rect 33459 12733 33471 12767
rect 33413 12727 33471 12733
rect 30760 12668 31754 12696
rect 26108 12656 26114 12668
rect 15838 12588 15844 12640
rect 15896 12628 15902 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15896 12600 16129 12628
rect 15896 12588 15902 12600
rect 16117 12597 16129 12600
rect 16163 12597 16175 12631
rect 16117 12591 16175 12597
rect 26973 12631 27031 12637
rect 26973 12597 26985 12631
rect 27019 12628 27031 12631
rect 28350 12628 28356 12640
rect 27019 12600 28356 12628
rect 27019 12597 27031 12600
rect 26973 12591 27031 12597
rect 28350 12588 28356 12600
rect 28408 12588 28414 12640
rect 35161 12631 35219 12637
rect 35161 12597 35173 12631
rect 35207 12628 35219 12631
rect 35342 12628 35348 12640
rect 35207 12600 35348 12628
rect 35207 12597 35219 12600
rect 35161 12591 35219 12597
rect 35342 12588 35348 12600
rect 35400 12588 35406 12640
rect 1104 12538 37076 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 37076 12538
rect 1104 12464 37076 12486
rect 20980 12427 21038 12433
rect 20980 12393 20992 12427
rect 21026 12424 21038 12427
rect 22557 12427 22615 12433
rect 22557 12424 22569 12427
rect 21026 12396 22569 12424
rect 21026 12393 21038 12396
rect 20980 12387 21038 12393
rect 22557 12393 22569 12396
rect 22603 12393 22615 12427
rect 22557 12387 22615 12393
rect 29549 12427 29607 12433
rect 29549 12393 29561 12427
rect 29595 12424 29607 12427
rect 29638 12424 29644 12436
rect 29595 12396 29644 12424
rect 29595 12393 29607 12396
rect 29549 12387 29607 12393
rect 29638 12384 29644 12396
rect 29696 12384 29702 12436
rect 32766 12384 32772 12436
rect 32824 12424 32830 12436
rect 32824 12396 35480 12424
rect 32824 12384 32830 12396
rect 10318 12248 10324 12300
rect 10376 12288 10382 12300
rect 10376 12260 22232 12288
rect 10376 12248 10382 12260
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12220 15163 12223
rect 15194 12220 15200 12232
rect 15151 12192 15200 12220
rect 15151 12189 15163 12192
rect 15105 12183 15163 12189
rect 15194 12180 15200 12192
rect 15252 12180 15258 12232
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 15764 12152 15792 12183
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 16206 12220 16212 12232
rect 15896 12192 16212 12220
rect 15896 12180 15902 12192
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12220 18291 12223
rect 18598 12220 18604 12232
rect 18279 12192 18604 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 19610 12180 19616 12232
rect 19668 12180 19674 12232
rect 19794 12180 19800 12232
rect 19852 12220 19858 12232
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19852 12192 20085 12220
rect 19852 12180 19858 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20254 12180 20260 12232
rect 20312 12180 20318 12232
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12220 20407 12223
rect 20622 12220 20628 12232
rect 20395 12192 20628 12220
rect 20395 12189 20407 12192
rect 20349 12183 20407 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 20714 12180 20720 12232
rect 20772 12180 20778 12232
rect 22204 12220 22232 12260
rect 23014 12248 23020 12300
rect 23072 12248 23078 12300
rect 23201 12291 23259 12297
rect 23201 12257 23213 12291
rect 23247 12288 23259 12291
rect 23290 12288 23296 12300
rect 23247 12260 23296 12288
rect 23247 12257 23259 12260
rect 23201 12251 23259 12257
rect 23290 12248 23296 12260
rect 23348 12248 23354 12300
rect 24121 12291 24179 12297
rect 24121 12257 24133 12291
rect 24167 12288 24179 12291
rect 26050 12288 26056 12300
rect 24167 12260 26056 12288
rect 24167 12257 24179 12260
rect 24121 12251 24179 12257
rect 26050 12248 26056 12260
rect 26108 12248 26114 12300
rect 28350 12248 28356 12300
rect 28408 12248 28414 12300
rect 30558 12248 30564 12300
rect 30616 12288 30622 12300
rect 31297 12291 31355 12297
rect 31297 12288 31309 12291
rect 30616 12260 31309 12288
rect 30616 12248 30622 12260
rect 31297 12257 31309 12260
rect 31343 12288 31355 12291
rect 31386 12288 31392 12300
rect 31343 12260 31392 12288
rect 31343 12257 31355 12260
rect 31297 12251 31355 12257
rect 31386 12248 31392 12260
rect 31444 12248 31450 12300
rect 35452 12297 35480 12396
rect 35437 12291 35495 12297
rect 35437 12257 35449 12291
rect 35483 12257 35495 12291
rect 35437 12251 35495 12257
rect 25041 12223 25099 12229
rect 25041 12220 25053 12223
rect 22204 12192 25053 12220
rect 25041 12189 25053 12192
rect 25087 12189 25099 12223
rect 25041 12183 25099 12189
rect 28629 12223 28687 12229
rect 28629 12189 28641 12223
rect 28675 12189 28687 12223
rect 28629 12183 28687 12189
rect 16022 12152 16028 12164
rect 15764 12124 16028 12152
rect 16022 12112 16028 12124
rect 16080 12112 16086 12164
rect 16390 12112 16396 12164
rect 16448 12152 16454 12164
rect 16448 12124 16790 12152
rect 16448 12112 16454 12124
rect 17954 12112 17960 12164
rect 18012 12112 18018 12164
rect 21542 12112 21548 12164
rect 21600 12112 21606 12164
rect 26602 12112 26608 12164
rect 26660 12112 26666 12164
rect 27922 12124 28028 12152
rect 16485 12087 16543 12093
rect 16485 12053 16497 12087
rect 16531 12084 16543 12087
rect 17862 12084 17868 12096
rect 16531 12056 17868 12084
rect 16531 12053 16543 12056
rect 16485 12047 16543 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 22465 12087 22523 12093
rect 22465 12053 22477 12087
rect 22511 12084 22523 12087
rect 22922 12084 22928 12096
rect 22511 12056 22928 12084
rect 22511 12053 22523 12056
rect 22465 12047 22523 12053
rect 22922 12044 22928 12056
rect 22980 12044 22986 12096
rect 23106 12044 23112 12096
rect 23164 12084 23170 12096
rect 23477 12087 23535 12093
rect 23477 12084 23489 12087
rect 23164 12056 23489 12084
rect 23164 12044 23170 12056
rect 23477 12053 23489 12056
rect 23523 12053 23535 12087
rect 23477 12047 23535 12053
rect 23842 12044 23848 12096
rect 23900 12044 23906 12096
rect 23937 12087 23995 12093
rect 23937 12053 23949 12087
rect 23983 12084 23995 12087
rect 25038 12084 25044 12096
rect 23983 12056 25044 12084
rect 23983 12053 23995 12056
rect 23937 12047 23995 12053
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 26326 12044 26332 12096
rect 26384 12084 26390 12096
rect 26881 12087 26939 12093
rect 26881 12084 26893 12087
rect 26384 12056 26893 12084
rect 26384 12044 26390 12056
rect 26881 12053 26893 12056
rect 26927 12084 26939 12087
rect 27338 12084 27344 12096
rect 26927 12056 27344 12084
rect 26927 12053 26939 12056
rect 26881 12047 26939 12053
rect 27338 12044 27344 12056
rect 27396 12044 27402 12096
rect 27430 12044 27436 12096
rect 27488 12084 27494 12096
rect 28000 12084 28028 12124
rect 28442 12112 28448 12164
rect 28500 12152 28506 12164
rect 28644 12152 28672 12183
rect 34514 12180 34520 12232
rect 34572 12180 34578 12232
rect 34606 12180 34612 12232
rect 34664 12220 34670 12232
rect 35161 12223 35219 12229
rect 35161 12220 35173 12223
rect 34664 12192 35173 12220
rect 34664 12180 34670 12192
rect 35161 12189 35173 12192
rect 35207 12189 35219 12223
rect 35161 12183 35219 12189
rect 35342 12180 35348 12232
rect 35400 12180 35406 12232
rect 28500 12124 28672 12152
rect 28500 12112 28506 12124
rect 30006 12112 30012 12164
rect 30064 12112 30070 12164
rect 31018 12112 31024 12164
rect 31076 12112 31082 12164
rect 33594 12112 33600 12164
rect 33652 12112 33658 12164
rect 34241 12155 34299 12161
rect 34241 12121 34253 12155
rect 34287 12152 34299 12155
rect 34701 12155 34759 12161
rect 34701 12152 34713 12155
rect 34287 12124 34713 12152
rect 34287 12121 34299 12124
rect 34241 12115 34299 12121
rect 34701 12121 34713 12124
rect 34747 12121 34759 12155
rect 34701 12115 34759 12121
rect 28994 12084 29000 12096
rect 27488 12056 29000 12084
rect 27488 12044 27494 12056
rect 28994 12044 29000 12056
rect 29052 12044 29058 12096
rect 1104 11994 37076 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 37076 11994
rect 1104 11920 37076 11942
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 16022 11880 16028 11892
rect 15703 11852 16028 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 16022 11840 16028 11852
rect 16080 11880 16086 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 16080 11852 16129 11880
rect 16080 11840 16086 11852
rect 16117 11849 16129 11852
rect 16163 11849 16175 11883
rect 16117 11843 16175 11849
rect 16206 11840 16212 11892
rect 16264 11840 16270 11892
rect 23842 11840 23848 11892
rect 23900 11880 23906 11892
rect 24305 11883 24363 11889
rect 24305 11880 24317 11883
rect 23900 11852 24317 11880
rect 23900 11840 23906 11852
rect 24305 11849 24317 11852
rect 24351 11880 24363 11883
rect 25498 11880 25504 11892
rect 24351 11852 25504 11880
rect 24351 11849 24363 11852
rect 24305 11843 24363 11849
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 27249 11883 27307 11889
rect 27249 11849 27261 11883
rect 27295 11880 27307 11883
rect 27706 11880 27712 11892
rect 27295 11852 27712 11880
rect 27295 11849 27307 11852
rect 27249 11843 27307 11849
rect 27706 11840 27712 11852
rect 27764 11840 27770 11892
rect 28994 11880 29000 11892
rect 28368 11852 29000 11880
rect 16390 11812 16396 11824
rect 15410 11784 16396 11812
rect 16390 11772 16396 11784
rect 16448 11772 16454 11824
rect 17034 11772 17040 11824
rect 17092 11812 17098 11824
rect 17497 11815 17555 11821
rect 17497 11812 17509 11815
rect 17092 11784 17509 11812
rect 17092 11772 17098 11784
rect 17497 11781 17509 11784
rect 17543 11781 17555 11815
rect 17497 11775 17555 11781
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 22833 11815 22891 11821
rect 17920 11784 18184 11812
rect 17920 11772 17926 11784
rect 17957 11747 18015 11753
rect 17957 11713 17969 11747
rect 18003 11744 18015 11747
rect 18046 11744 18052 11756
rect 18003 11716 18052 11744
rect 18003 11713 18015 11716
rect 17957 11707 18015 11713
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18156 11753 18184 11784
rect 22833 11781 22845 11815
rect 22879 11812 22891 11815
rect 23106 11812 23112 11824
rect 22879 11784 23112 11812
rect 22879 11781 22891 11784
rect 22833 11775 22891 11781
rect 23106 11772 23112 11784
rect 23164 11772 23170 11824
rect 24578 11812 24584 11824
rect 24058 11784 24584 11812
rect 24578 11772 24584 11784
rect 24636 11772 24642 11824
rect 25958 11812 25964 11824
rect 25898 11784 25964 11812
rect 25958 11772 25964 11784
rect 26016 11812 26022 11824
rect 26234 11812 26240 11824
rect 26016 11784 26240 11812
rect 26016 11772 26022 11784
rect 26234 11772 26240 11784
rect 26292 11812 26298 11824
rect 27430 11812 27436 11824
rect 26292 11784 27436 11812
rect 26292 11772 26298 11784
rect 27430 11772 27436 11784
rect 27488 11772 27494 11824
rect 28368 11812 28396 11852
rect 28994 11840 29000 11852
rect 29052 11880 29058 11892
rect 30006 11880 30012 11892
rect 29052 11852 30012 11880
rect 29052 11840 29058 11852
rect 30006 11840 30012 11852
rect 30064 11840 30070 11892
rect 28290 11784 28396 11812
rect 28442 11772 28448 11824
rect 28500 11812 28506 11824
rect 28500 11784 29040 11812
rect 28500 11772 28506 11784
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 18233 11747 18291 11753
rect 18233 11713 18245 11747
rect 18279 11744 18291 11747
rect 18506 11744 18512 11756
rect 18279 11716 18512 11744
rect 18279 11713 18291 11716
rect 18233 11707 18291 11713
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 19978 11704 19984 11756
rect 20036 11704 20042 11756
rect 29012 11753 29040 11784
rect 28997 11747 29055 11753
rect 28997 11713 29009 11747
rect 29043 11713 29055 11747
rect 28997 11707 29055 11713
rect 30653 11747 30711 11753
rect 30653 11713 30665 11747
rect 30699 11713 30711 11747
rect 30653 11707 30711 11713
rect 31205 11747 31263 11753
rect 31205 11713 31217 11747
rect 31251 11713 31263 11747
rect 31205 11707 31263 11713
rect 31573 11747 31631 11753
rect 31573 11713 31585 11747
rect 31619 11744 31631 11747
rect 32122 11744 32128 11756
rect 31619 11716 32128 11744
rect 31619 11713 31631 11716
rect 31573 11707 31631 11713
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13780 11648 13921 11676
rect 13780 11636 13786 11648
rect 13909 11645 13921 11648
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14231 11648 15792 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 15764 11617 15792 11648
rect 16206 11636 16212 11688
rect 16264 11676 16270 11688
rect 16301 11679 16359 11685
rect 16301 11676 16313 11679
rect 16264 11648 16313 11676
rect 16264 11636 16270 11648
rect 16301 11645 16313 11648
rect 16347 11676 16359 11679
rect 16482 11676 16488 11688
rect 16347 11648 16488 11676
rect 16347 11645 16359 11648
rect 16301 11639 16359 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 18598 11636 18604 11688
rect 18656 11636 18662 11688
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 19334 11676 19340 11688
rect 18923 11648 19340 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 19334 11636 19340 11648
rect 19392 11636 19398 11688
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 21910 11676 21916 11688
rect 20772 11648 21916 11676
rect 20772 11636 20778 11648
rect 21910 11636 21916 11648
rect 21968 11676 21974 11688
rect 22557 11679 22615 11685
rect 22557 11676 22569 11679
rect 21968 11648 22569 11676
rect 21968 11636 21974 11648
rect 22557 11645 22569 11648
rect 22603 11645 22615 11679
rect 22557 11639 22615 11645
rect 24394 11636 24400 11688
rect 24452 11636 24458 11688
rect 24670 11636 24676 11688
rect 24728 11636 24734 11688
rect 28074 11636 28080 11688
rect 28132 11676 28138 11688
rect 28721 11679 28779 11685
rect 28721 11676 28733 11679
rect 28132 11648 28733 11676
rect 28132 11636 28138 11648
rect 28721 11645 28733 11648
rect 28767 11645 28779 11679
rect 28721 11639 28779 11645
rect 15749 11611 15807 11617
rect 15749 11577 15761 11611
rect 15795 11577 15807 11611
rect 30668 11608 30696 11707
rect 31220 11676 31248 11707
rect 32122 11704 32128 11716
rect 32180 11704 32186 11756
rect 31297 11679 31355 11685
rect 31297 11676 31309 11679
rect 31220 11648 31309 11676
rect 31297 11645 31309 11648
rect 31343 11645 31355 11679
rect 31297 11639 31355 11645
rect 31481 11679 31539 11685
rect 31481 11645 31493 11679
rect 31527 11645 31539 11679
rect 31481 11639 31539 11645
rect 31202 11608 31208 11620
rect 30668 11580 31208 11608
rect 15749 11571 15807 11577
rect 31202 11568 31208 11580
rect 31260 11608 31266 11620
rect 31496 11608 31524 11639
rect 31662 11636 31668 11688
rect 31720 11636 31726 11688
rect 31754 11636 31760 11688
rect 31812 11636 31818 11688
rect 31260 11580 31524 11608
rect 31260 11568 31266 11580
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 20254 11540 20260 11552
rect 20128 11512 20260 11540
rect 20128 11500 20134 11512
rect 20254 11500 20260 11512
rect 20312 11540 20318 11552
rect 20349 11543 20407 11549
rect 20349 11540 20361 11543
rect 20312 11512 20361 11540
rect 20312 11500 20318 11512
rect 20349 11509 20361 11512
rect 20395 11509 20407 11543
rect 20349 11503 20407 11509
rect 25038 11500 25044 11552
rect 25096 11540 25102 11552
rect 26145 11543 26203 11549
rect 26145 11540 26157 11543
rect 25096 11512 26157 11540
rect 25096 11500 25102 11512
rect 26145 11509 26157 11512
rect 26191 11509 26203 11543
rect 26145 11503 26203 11509
rect 30834 11500 30840 11552
rect 30892 11500 30898 11552
rect 31110 11500 31116 11552
rect 31168 11500 31174 11552
rect 1104 11450 37076 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 37076 11450
rect 1104 11376 37076 11398
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 21358 11336 21364 11348
rect 16264 11308 21364 11336
rect 16264 11296 16270 11308
rect 16301 11271 16359 11277
rect 16301 11237 16313 11271
rect 16347 11268 16359 11271
rect 16758 11268 16764 11280
rect 16347 11240 16764 11268
rect 16347 11237 16359 11240
rect 16301 11231 16359 11237
rect 16758 11228 16764 11240
rect 16816 11228 16822 11280
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 16172 11172 18061 11200
rect 16172 11160 16178 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 18892 11200 18920 11308
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 24670 11296 24676 11348
rect 24728 11296 24734 11348
rect 26237 11339 26295 11345
rect 26237 11305 26249 11339
rect 26283 11336 26295 11339
rect 28457 11339 28515 11345
rect 28457 11336 28469 11339
rect 26283 11308 28469 11336
rect 26283 11305 26295 11308
rect 26237 11299 26295 11305
rect 28457 11305 28469 11308
rect 28503 11305 28515 11339
rect 28457 11299 28515 11305
rect 31110 11296 31116 11348
rect 31168 11336 31174 11348
rect 31646 11339 31704 11345
rect 31646 11336 31658 11339
rect 31168 11308 31658 11336
rect 31168 11296 31174 11308
rect 31646 11305 31658 11308
rect 31692 11305 31704 11339
rect 31646 11299 31704 11305
rect 32122 11296 32128 11348
rect 32180 11336 32186 11348
rect 33137 11339 33195 11345
rect 33137 11336 33149 11339
rect 32180 11308 33149 11336
rect 32180 11296 32186 11308
rect 33137 11305 33149 11308
rect 33183 11305 33195 11339
rect 33137 11299 33195 11305
rect 23290 11228 23296 11280
rect 23348 11268 23354 11280
rect 26970 11268 26976 11280
rect 23348 11240 23888 11268
rect 23348 11228 23354 11240
rect 18831 11172 18920 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 18064 11132 18092 11163
rect 20162 11160 20168 11212
rect 20220 11200 20226 11212
rect 20993 11203 21051 11209
rect 20993 11200 21005 11203
rect 20220 11172 21005 11200
rect 20220 11160 20226 11172
rect 20993 11169 21005 11172
rect 21039 11169 21051 11203
rect 20993 11163 21051 11169
rect 21266 11160 21272 11212
rect 21324 11160 21330 11212
rect 22572 11172 22876 11200
rect 22572 11144 22600 11172
rect 18598 11132 18604 11144
rect 18064 11104 18604 11132
rect 18598 11092 18604 11104
rect 18656 11132 18662 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18656 11104 19257 11132
rect 18656 11092 18662 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 22005 11135 22063 11141
rect 22005 11101 22017 11135
rect 22051 11132 22063 11135
rect 22094 11132 22100 11144
rect 22051 11104 22100 11132
rect 22051 11101 22063 11104
rect 22005 11095 22063 11101
rect 22094 11092 22100 11104
rect 22152 11092 22158 11144
rect 22278 11092 22284 11144
rect 22336 11132 22342 11144
rect 22465 11135 22523 11141
rect 22465 11132 22477 11135
rect 22336 11104 22477 11132
rect 22336 11092 22342 11104
rect 22465 11101 22477 11104
rect 22511 11101 22523 11135
rect 22465 11095 22523 11101
rect 22554 11092 22560 11144
rect 22612 11092 22618 11144
rect 22741 11135 22799 11141
rect 22741 11101 22753 11135
rect 22787 11101 22799 11135
rect 22848 11132 22876 11172
rect 22922 11160 22928 11212
rect 22980 11200 22986 11212
rect 23860 11209 23888 11240
rect 26712 11240 26976 11268
rect 23753 11203 23811 11209
rect 23753 11200 23765 11203
rect 22980 11172 23765 11200
rect 22980 11160 22986 11172
rect 23753 11169 23765 11172
rect 23799 11169 23811 11203
rect 23753 11163 23811 11169
rect 23845 11203 23903 11209
rect 23845 11169 23857 11203
rect 23891 11169 23903 11203
rect 23845 11163 23903 11169
rect 25314 11160 25320 11212
rect 25372 11160 25378 11212
rect 26712 11209 26740 11240
rect 26970 11228 26976 11240
rect 27028 11228 27034 11280
rect 34698 11268 34704 11280
rect 33704 11240 34704 11268
rect 26697 11203 26755 11209
rect 26697 11169 26709 11203
rect 26743 11169 26755 11203
rect 27706 11200 27712 11212
rect 26697 11163 26755 11169
rect 27172 11172 27712 11200
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 22848 11104 23673 11132
rect 22741 11095 22799 11101
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 16390 11024 16396 11076
rect 16448 11064 16454 11076
rect 17773 11067 17831 11073
rect 17773 11064 17785 11067
rect 16448 11036 16606 11064
rect 17604 11036 17785 11064
rect 16448 11024 16454 11036
rect 17604 11008 17632 11036
rect 17773 11033 17785 11036
rect 17819 11033 17831 11067
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 17773 11027 17831 11033
rect 18064 11036 18521 11064
rect 17586 10956 17592 11008
rect 17644 10956 17650 11008
rect 17862 10956 17868 11008
rect 17920 10996 17926 11008
rect 18064 10996 18092 11036
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 18509 11027 18567 11033
rect 19518 11024 19524 11076
rect 19576 11024 19582 11076
rect 19978 11024 19984 11076
rect 20036 11024 20042 11076
rect 22756 11064 22784 11095
rect 25038 11092 25044 11144
rect 25096 11092 25102 11144
rect 26234 11092 26240 11144
rect 26292 11132 26298 11144
rect 26789 11135 26847 11141
rect 26789 11132 26801 11135
rect 26292 11104 26801 11132
rect 26292 11092 26298 11104
rect 26789 11101 26801 11104
rect 26835 11101 26847 11135
rect 26789 11095 26847 11101
rect 22830 11064 22836 11076
rect 22756 11036 22836 11064
rect 22830 11024 22836 11036
rect 22888 11024 22894 11076
rect 23198 11024 23204 11076
rect 23256 11024 23262 11076
rect 23382 11024 23388 11076
rect 23440 11064 23446 11076
rect 26697 11067 26755 11073
rect 23440 11036 26234 11064
rect 23440 11024 23446 11036
rect 17920 10968 18092 10996
rect 17920 10956 17926 10968
rect 18138 10956 18144 11008
rect 18196 10956 18202 11008
rect 18601 10999 18659 11005
rect 18601 10965 18613 10999
rect 18647 10996 18659 10999
rect 18690 10996 18696 11008
rect 18647 10968 18696 10996
rect 18647 10965 18659 10968
rect 18601 10959 18659 10965
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 22186 10956 22192 11008
rect 22244 10996 22250 11008
rect 23293 10999 23351 11005
rect 23293 10996 23305 10999
rect 22244 10968 23305 10996
rect 22244 10956 22250 10968
rect 23293 10965 23305 10968
rect 23339 10965 23351 10999
rect 23293 10959 23351 10965
rect 25130 10956 25136 11008
rect 25188 10956 25194 11008
rect 26206 10996 26234 11036
rect 26697 11033 26709 11067
rect 26743 11064 26755 11067
rect 27172 11064 27200 11172
rect 27706 11160 27712 11172
rect 27764 11160 27770 11212
rect 28442 11160 28448 11212
rect 28500 11200 28506 11212
rect 28721 11203 28779 11209
rect 28721 11200 28733 11203
rect 28500 11172 28733 11200
rect 28500 11160 28506 11172
rect 28721 11169 28733 11172
rect 28767 11200 28779 11203
rect 29549 11203 29607 11209
rect 29549 11200 29561 11203
rect 28767 11172 29561 11200
rect 28767 11169 28779 11172
rect 28721 11163 28779 11169
rect 29549 11169 29561 11172
rect 29595 11169 29607 11203
rect 29549 11163 29607 11169
rect 29825 11203 29883 11209
rect 29825 11169 29837 11203
rect 29871 11200 29883 11203
rect 30374 11200 30380 11212
rect 29871 11172 30380 11200
rect 29871 11169 29883 11172
rect 29825 11163 29883 11169
rect 30374 11160 30380 11172
rect 30432 11160 30438 11212
rect 31386 11160 31392 11212
rect 31444 11200 31450 11212
rect 32674 11200 32680 11212
rect 31444 11172 32680 11200
rect 31444 11160 31450 11172
rect 32674 11160 32680 11172
rect 32732 11200 32738 11212
rect 33042 11200 33048 11212
rect 32732 11172 33048 11200
rect 32732 11160 32738 11172
rect 33042 11160 33048 11172
rect 33100 11160 33106 11212
rect 33704 11141 33732 11240
rect 34698 11228 34704 11240
rect 34756 11228 34762 11280
rect 35434 11200 35440 11212
rect 33888 11172 35440 11200
rect 33888 11141 33916 11172
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 33689 11135 33747 11141
rect 33689 11101 33701 11135
rect 33735 11101 33747 11135
rect 33689 11095 33747 11101
rect 33873 11135 33931 11141
rect 33873 11101 33885 11135
rect 33919 11101 33931 11135
rect 33873 11095 33931 11101
rect 33962 11092 33968 11144
rect 34020 11092 34026 11144
rect 34333 11135 34391 11141
rect 34333 11101 34345 11135
rect 34379 11101 34391 11135
rect 34333 11095 34391 11101
rect 28994 11064 29000 11076
rect 26743 11036 27200 11064
rect 28014 11036 29000 11064
rect 26743 11033 26755 11036
rect 26697 11027 26755 11033
rect 28994 11024 29000 11036
rect 29052 11024 29058 11076
rect 33229 11067 33287 11073
rect 31050 11036 32076 11064
rect 32890 11036 33180 11064
rect 26602 10996 26608 11008
rect 26206 10968 26608 10996
rect 26602 10956 26608 10968
rect 26660 10956 26666 11008
rect 31297 10999 31355 11005
rect 31297 10965 31309 10999
rect 31343 10996 31355 10999
rect 31662 10996 31668 11008
rect 31343 10968 31668 10996
rect 31343 10965 31355 10968
rect 31297 10959 31355 10965
rect 31662 10956 31668 10968
rect 31720 10996 31726 11008
rect 31846 10996 31852 11008
rect 31720 10968 31852 10996
rect 31720 10956 31726 10968
rect 31846 10956 31852 10968
rect 31904 10956 31910 11008
rect 32048 10996 32076 11036
rect 32968 10996 32996 11036
rect 32048 10968 32996 10996
rect 33152 10996 33180 11036
rect 33229 11033 33241 11067
rect 33275 11064 33287 11067
rect 34348 11064 34376 11095
rect 33275 11036 34376 11064
rect 33275 11033 33287 11036
rect 33229 11027 33287 11033
rect 33594 10996 33600 11008
rect 33152 10968 33600 10996
rect 33594 10956 33600 10968
rect 33652 10996 33658 11008
rect 34238 10996 34244 11008
rect 33652 10968 34244 10996
rect 33652 10956 33658 10968
rect 34238 10956 34244 10968
rect 34296 10956 34302 11008
rect 34422 10956 34428 11008
rect 34480 10956 34486 11008
rect 1104 10906 37076 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 37076 10906
rect 1104 10832 37076 10854
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15473 10795 15531 10801
rect 15473 10792 15485 10795
rect 15436 10764 15485 10792
rect 15436 10752 15442 10764
rect 15473 10761 15485 10764
rect 15519 10792 15531 10795
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15519 10764 15945 10792
rect 15519 10761 15531 10764
rect 15473 10755 15531 10761
rect 15933 10761 15945 10764
rect 15979 10761 15991 10795
rect 15933 10755 15991 10761
rect 16022 10752 16028 10804
rect 16080 10752 16086 10804
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 18046 10792 18052 10804
rect 17644 10764 18052 10792
rect 17644 10752 17650 10764
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 19058 10752 19064 10804
rect 19116 10792 19122 10804
rect 23842 10792 23848 10804
rect 19116 10764 23848 10792
rect 19116 10752 19122 10764
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 26326 10752 26332 10804
rect 26384 10752 26390 10804
rect 30374 10752 30380 10804
rect 30432 10801 30438 10804
rect 30432 10792 30441 10801
rect 34422 10792 34428 10804
rect 30432 10764 30477 10792
rect 30760 10764 31892 10792
rect 30432 10755 30441 10764
rect 30432 10752 30438 10755
rect 16390 10724 16396 10736
rect 15226 10696 16396 10724
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 17954 10684 17960 10736
rect 18012 10724 18018 10736
rect 18233 10727 18291 10733
rect 18233 10724 18245 10727
rect 18012 10696 18245 10724
rect 18012 10684 18018 10696
rect 18233 10693 18245 10696
rect 18279 10693 18291 10727
rect 18233 10687 18291 10693
rect 18414 10684 18420 10736
rect 18472 10724 18478 10736
rect 21085 10727 21143 10733
rect 21085 10724 21097 10727
rect 18472 10696 21097 10724
rect 18472 10684 18478 10696
rect 21085 10693 21097 10696
rect 21131 10693 21143 10727
rect 21085 10687 21143 10693
rect 22094 10684 22100 10736
rect 22152 10724 22158 10736
rect 26421 10727 26479 10733
rect 22152 10696 23796 10724
rect 22152 10684 22158 10696
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 17402 10656 17408 10668
rect 16816 10628 17408 10656
rect 16816 10616 16822 10628
rect 17402 10616 17408 10628
rect 17460 10656 17466 10668
rect 17589 10659 17647 10665
rect 17589 10656 17601 10659
rect 17460 10628 17601 10656
rect 17460 10616 17466 10628
rect 17589 10625 17601 10628
rect 17635 10625 17647 10659
rect 17589 10619 17647 10625
rect 17773 10659 17831 10665
rect 17773 10625 17785 10659
rect 17819 10625 17831 10659
rect 17773 10619 17831 10625
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10588 14059 10591
rect 14047 10560 15608 10588
rect 14047 10557 14059 10560
rect 14001 10551 14059 10557
rect 15580 10529 15608 10560
rect 16206 10548 16212 10600
rect 16264 10548 16270 10600
rect 17497 10591 17555 10597
rect 17497 10557 17509 10591
rect 17543 10588 17555 10591
rect 17678 10588 17684 10600
rect 17543 10560 17684 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 17678 10548 17684 10560
rect 17736 10548 17742 10600
rect 17788 10588 17816 10619
rect 18874 10616 18880 10668
rect 18932 10656 18938 10668
rect 21266 10656 21272 10668
rect 18932 10628 21272 10656
rect 18932 10616 18938 10628
rect 21266 10616 21272 10628
rect 21324 10656 21330 10668
rect 22848 10665 22876 10696
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21324 10628 22017 10656
rect 21324 10616 21330 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10625 22891 10659
rect 22833 10619 22891 10625
rect 23293 10659 23351 10665
rect 23293 10625 23305 10659
rect 23339 10656 23351 10659
rect 23658 10656 23664 10668
rect 23339 10628 23664 10656
rect 23339 10625 23351 10628
rect 23293 10619 23351 10625
rect 23658 10616 23664 10628
rect 23716 10616 23722 10668
rect 18230 10588 18236 10600
rect 17788 10560 18236 10588
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 20806 10548 20812 10600
rect 20864 10588 20870 10600
rect 21177 10591 21235 10597
rect 21177 10588 21189 10591
rect 20864 10560 21189 10588
rect 20864 10548 20870 10560
rect 21177 10557 21189 10560
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21358 10548 21364 10600
rect 21416 10548 21422 10600
rect 22278 10548 22284 10600
rect 22336 10588 22342 10600
rect 23385 10591 23443 10597
rect 23385 10588 23397 10591
rect 22336 10560 23397 10588
rect 22336 10548 22342 10560
rect 23385 10557 23397 10560
rect 23431 10557 23443 10591
rect 23385 10551 23443 10557
rect 23477 10591 23535 10597
rect 23477 10557 23489 10591
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 15565 10523 15623 10529
rect 15565 10489 15577 10523
rect 15611 10489 15623 10523
rect 21376 10520 21404 10548
rect 23290 10520 23296 10532
rect 21376 10492 23296 10520
rect 15565 10483 15623 10489
rect 23290 10480 23296 10492
rect 23348 10520 23354 10532
rect 23492 10520 23520 10551
rect 23348 10492 23520 10520
rect 23768 10520 23796 10696
rect 26421 10693 26433 10727
rect 26467 10724 26479 10727
rect 28626 10724 28632 10736
rect 26467 10696 28632 10724
rect 26467 10693 26479 10696
rect 26421 10687 26479 10693
rect 28626 10684 28632 10696
rect 28684 10684 28690 10736
rect 30006 10724 30012 10736
rect 29946 10696 30012 10724
rect 30006 10684 30012 10696
rect 30064 10684 30070 10736
rect 30469 10727 30527 10733
rect 30469 10693 30481 10727
rect 30515 10724 30527 10727
rect 30760 10724 30788 10764
rect 31864 10736 31892 10764
rect 32968 10764 34428 10792
rect 30515 10696 30788 10724
rect 30515 10693 30527 10696
rect 30469 10687 30527 10693
rect 30834 10684 30840 10736
rect 30892 10724 30898 10736
rect 31665 10727 31723 10733
rect 31665 10724 31677 10727
rect 30892 10696 31677 10724
rect 30892 10684 30898 10696
rect 31665 10693 31677 10696
rect 31711 10693 31723 10727
rect 31665 10687 31723 10693
rect 31846 10684 31852 10736
rect 31904 10684 31910 10736
rect 32968 10733 32996 10764
rect 34422 10752 34428 10764
rect 34480 10752 34486 10804
rect 32953 10727 33011 10733
rect 32953 10693 32965 10727
rect 32999 10693 33011 10727
rect 32953 10687 33011 10693
rect 33594 10684 33600 10736
rect 33652 10684 33658 10736
rect 34238 10684 34244 10736
rect 34296 10724 34302 10736
rect 34296 10696 35282 10724
rect 34296 10684 34302 10696
rect 25130 10616 25136 10668
rect 25188 10616 25194 10668
rect 25225 10659 25283 10665
rect 25225 10625 25237 10659
rect 25271 10656 25283 10659
rect 26142 10656 26148 10668
rect 25271 10628 26148 10656
rect 25271 10625 25283 10628
rect 25225 10619 25283 10625
rect 26142 10616 26148 10628
rect 26200 10616 26206 10668
rect 26602 10616 26608 10668
rect 26660 10656 26666 10668
rect 27433 10659 27491 10665
rect 27433 10656 27445 10659
rect 26660 10628 27445 10656
rect 26660 10616 26666 10628
rect 27433 10625 27445 10628
rect 27479 10656 27491 10659
rect 27982 10656 27988 10668
rect 27479 10628 27988 10656
rect 27479 10625 27491 10628
rect 27433 10619 27491 10625
rect 27982 10616 27988 10628
rect 28040 10616 28046 10668
rect 30285 10659 30343 10665
rect 30285 10625 30297 10659
rect 30331 10625 30343 10659
rect 30285 10619 30343 10625
rect 30561 10659 30619 10665
rect 30561 10625 30573 10659
rect 30607 10625 30619 10659
rect 30561 10619 30619 10625
rect 25314 10548 25320 10600
rect 25372 10588 25378 10600
rect 25409 10591 25467 10597
rect 25409 10588 25421 10591
rect 25372 10560 25421 10588
rect 25372 10548 25378 10560
rect 25409 10557 25421 10560
rect 25455 10588 25467 10591
rect 26050 10588 26056 10600
rect 25455 10560 26056 10588
rect 25455 10557 25467 10560
rect 25409 10551 25467 10557
rect 26050 10548 26056 10560
rect 26108 10548 26114 10600
rect 26234 10548 26240 10600
rect 26292 10548 26298 10600
rect 26970 10548 26976 10600
rect 27028 10588 27034 10600
rect 28169 10591 28227 10597
rect 28169 10588 28181 10591
rect 27028 10560 28181 10588
rect 27028 10548 27034 10560
rect 28169 10557 28181 10560
rect 28215 10588 28227 10591
rect 28442 10588 28448 10600
rect 28215 10560 28448 10588
rect 28215 10557 28227 10560
rect 28169 10551 28227 10557
rect 28442 10548 28448 10560
rect 28500 10548 28506 10600
rect 28718 10548 28724 10600
rect 28776 10548 28782 10600
rect 26694 10520 26700 10532
rect 23768 10492 26700 10520
rect 23348 10480 23354 10492
rect 17954 10412 17960 10464
rect 18012 10452 18018 10464
rect 19058 10452 19064 10464
rect 18012 10424 19064 10452
rect 18012 10412 18018 10424
rect 19058 10412 19064 10424
rect 19116 10452 19122 10464
rect 20165 10455 20223 10461
rect 20165 10452 20177 10455
rect 19116 10424 20177 10452
rect 19116 10412 19122 10424
rect 20165 10421 20177 10424
rect 20211 10421 20223 10455
rect 20165 10415 20223 10421
rect 20714 10412 20720 10464
rect 20772 10412 20778 10464
rect 22922 10412 22928 10464
rect 22980 10412 22986 10464
rect 23492 10452 23520 10492
rect 26694 10480 26700 10492
rect 26752 10480 26758 10532
rect 30300 10520 30328 10619
rect 30576 10588 30604 10619
rect 31478 10616 31484 10668
rect 31536 10656 31542 10668
rect 31941 10659 31999 10665
rect 31536 10628 31800 10656
rect 31536 10616 31542 10628
rect 31202 10588 31208 10600
rect 30576 10560 31208 10588
rect 31202 10548 31208 10560
rect 31260 10548 31266 10600
rect 31665 10523 31723 10529
rect 31665 10520 31677 10523
rect 30300 10492 31677 10520
rect 31665 10489 31677 10492
rect 31711 10489 31723 10523
rect 31772 10520 31800 10628
rect 31941 10625 31953 10659
rect 31987 10656 31999 10659
rect 32490 10656 32496 10668
rect 31987 10628 32496 10656
rect 31987 10625 31999 10628
rect 31941 10619 31999 10625
rect 32490 10616 32496 10628
rect 32548 10616 32554 10668
rect 32674 10616 32680 10668
rect 32732 10616 32738 10668
rect 33410 10548 33416 10600
rect 33468 10588 33474 10600
rect 34514 10588 34520 10600
rect 33468 10560 34520 10588
rect 33468 10548 33474 10560
rect 34514 10548 34520 10560
rect 34572 10548 34578 10600
rect 34790 10548 34796 10600
rect 34848 10548 34854 10600
rect 32398 10520 32404 10532
rect 31772 10492 32404 10520
rect 31665 10483 31723 10489
rect 32398 10480 32404 10492
rect 32456 10480 32462 10532
rect 23934 10452 23940 10464
rect 23492 10424 23940 10452
rect 23934 10412 23940 10424
rect 23992 10412 23998 10464
rect 24670 10412 24676 10464
rect 24728 10452 24734 10464
rect 24765 10455 24823 10461
rect 24765 10452 24777 10455
rect 24728 10424 24777 10452
rect 24728 10412 24734 10424
rect 24765 10421 24777 10424
rect 24811 10421 24823 10455
rect 24765 10415 24823 10421
rect 26786 10412 26792 10464
rect 26844 10412 26850 10464
rect 30193 10455 30251 10461
rect 30193 10421 30205 10455
rect 30239 10452 30251 10455
rect 30374 10452 30380 10464
rect 30239 10424 30380 10452
rect 30239 10421 30251 10424
rect 30193 10415 30251 10421
rect 30374 10412 30380 10424
rect 30432 10412 30438 10464
rect 33962 10412 33968 10464
rect 34020 10452 34026 10464
rect 34422 10452 34428 10464
rect 34020 10424 34428 10452
rect 34020 10412 34026 10424
rect 34422 10412 34428 10424
rect 34480 10412 34486 10464
rect 35342 10412 35348 10464
rect 35400 10452 35406 10464
rect 36265 10455 36323 10461
rect 36265 10452 36277 10455
rect 35400 10424 36277 10452
rect 35400 10412 35406 10424
rect 36265 10421 36277 10424
rect 36311 10421 36323 10455
rect 36265 10415 36323 10421
rect 1104 10362 37076 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 37076 10362
rect 1104 10288 37076 10310
rect 17862 10208 17868 10260
rect 17920 10208 17926 10260
rect 20888 10251 20946 10257
rect 20888 10217 20900 10251
rect 20934 10248 20946 10251
rect 22186 10248 22192 10260
rect 20934 10220 22192 10248
rect 20934 10217 20946 10220
rect 20888 10211 20946 10217
rect 22186 10208 22192 10220
rect 22244 10208 22250 10260
rect 22373 10251 22431 10257
rect 22373 10217 22385 10251
rect 22419 10248 22431 10251
rect 22554 10248 22560 10260
rect 22419 10220 22560 10248
rect 22419 10217 22431 10220
rect 22373 10211 22431 10217
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 25130 10208 25136 10260
rect 25188 10248 25194 10260
rect 26145 10251 26203 10257
rect 26145 10248 26157 10251
rect 25188 10220 26157 10248
rect 25188 10208 25194 10220
rect 26145 10217 26157 10220
rect 26191 10217 26203 10251
rect 26145 10211 26203 10217
rect 28718 10208 28724 10260
rect 28776 10248 28782 10260
rect 30285 10251 30343 10257
rect 30285 10248 30297 10251
rect 28776 10220 30297 10248
rect 28776 10208 28782 10220
rect 30285 10217 30297 10220
rect 30331 10217 30343 10251
rect 30285 10211 30343 10217
rect 31754 10208 31760 10260
rect 31812 10208 31818 10260
rect 31846 10208 31852 10260
rect 31904 10248 31910 10260
rect 31904 10220 32352 10248
rect 31904 10208 31910 10220
rect 29917 10183 29975 10189
rect 29917 10149 29929 10183
rect 29963 10149 29975 10183
rect 29917 10143 29975 10149
rect 15930 10112 15936 10124
rect 15212 10084 15936 10112
rect 15212 10053 15240 10084
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 18138 10112 18144 10124
rect 16439 10084 18144 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 19061 10115 19119 10121
rect 18288 10084 18644 10112
rect 18288 10072 18294 10084
rect 15197 10047 15255 10053
rect 15197 10013 15209 10047
rect 15243 10013 15255 10047
rect 15197 10007 15255 10013
rect 15378 10004 15384 10056
rect 15436 10004 15442 10056
rect 15470 10004 15476 10056
rect 15528 10004 15534 10056
rect 16114 10004 16120 10056
rect 16172 10004 16178 10056
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 14737 9979 14795 9985
rect 14737 9976 14749 9979
rect 13964 9948 14749 9976
rect 13964 9936 13970 9948
rect 14737 9945 14749 9948
rect 14783 9945 14795 9979
rect 14737 9939 14795 9945
rect 16390 9936 16396 9988
rect 16448 9976 16454 9988
rect 18340 9976 18368 10007
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 18616 10053 18644 10084
rect 19061 10081 19073 10115
rect 19107 10112 19119 10115
rect 19518 10112 19524 10124
rect 19107 10084 19524 10112
rect 19107 10081 19119 10084
rect 19061 10075 19119 10081
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 20070 10072 20076 10124
rect 20128 10072 20134 10124
rect 20625 10115 20683 10121
rect 20625 10081 20637 10115
rect 20671 10112 20683 10115
rect 21910 10112 21916 10124
rect 20671 10084 21916 10112
rect 20671 10081 20683 10084
rect 20625 10075 20683 10081
rect 21910 10072 21916 10084
rect 21968 10112 21974 10124
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 21968 10084 23305 10112
rect 21968 10072 21974 10084
rect 23293 10081 23305 10084
rect 23339 10112 23351 10115
rect 23566 10112 23572 10124
rect 23339 10084 23572 10112
rect 23339 10081 23351 10084
rect 23293 10075 23351 10081
rect 23566 10072 23572 10084
rect 23624 10112 23630 10124
rect 24394 10112 24400 10124
rect 23624 10084 24400 10112
rect 23624 10072 23630 10084
rect 24394 10072 24400 10084
rect 24452 10072 24458 10124
rect 24670 10072 24676 10124
rect 24728 10072 24734 10124
rect 29932 10112 29960 10143
rect 29932 10084 30328 10112
rect 18601 10047 18659 10053
rect 18601 10013 18613 10047
rect 18647 10013 18659 10047
rect 18601 10007 18659 10013
rect 19334 10004 19340 10056
rect 19392 10004 19398 10056
rect 19794 10004 19800 10056
rect 19852 10004 19858 10056
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20162 10044 20168 10056
rect 20027 10016 20168 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 19996 9976 20024 10007
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10044 22615 10047
rect 23014 10044 23020 10056
rect 22603 10016 23020 10044
rect 22603 10013 22615 10016
rect 22557 10007 22615 10013
rect 23014 10004 23020 10016
rect 23072 10044 23078 10056
rect 23382 10044 23388 10056
rect 23072 10016 23388 10044
rect 23072 10004 23078 10016
rect 23382 10004 23388 10016
rect 23440 10004 23446 10056
rect 26970 10004 26976 10056
rect 27028 10044 27034 10056
rect 27249 10047 27307 10053
rect 27249 10044 27261 10047
rect 27028 10016 27261 10044
rect 27028 10004 27034 10016
rect 27249 10013 27261 10016
rect 27295 10013 27307 10047
rect 27249 10007 27307 10013
rect 29638 10004 29644 10056
rect 29696 10044 29702 10056
rect 29917 10047 29975 10053
rect 29917 10044 29929 10047
rect 29696 10016 29929 10044
rect 29696 10004 29702 10016
rect 29917 10013 29929 10016
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 30190 10004 30196 10056
rect 30248 10004 30254 10056
rect 30300 10053 30328 10084
rect 31202 10072 31208 10124
rect 31260 10112 31266 10124
rect 31389 10115 31447 10121
rect 31389 10112 31401 10115
rect 31260 10084 31401 10112
rect 31260 10072 31266 10084
rect 31389 10081 31401 10084
rect 31435 10112 31447 10115
rect 32324 10112 32352 10220
rect 32490 10208 32496 10260
rect 32548 10248 32554 10260
rect 33686 10248 33692 10260
rect 32548 10220 33692 10248
rect 32548 10208 32554 10220
rect 33686 10208 33692 10220
rect 33744 10248 33750 10260
rect 34606 10248 34612 10260
rect 33744 10220 34612 10248
rect 33744 10208 33750 10220
rect 34606 10208 34612 10220
rect 34664 10208 34670 10260
rect 34790 10208 34796 10260
rect 34848 10248 34854 10260
rect 34977 10251 35035 10257
rect 34977 10248 34989 10251
rect 34848 10220 34989 10248
rect 34848 10208 34854 10220
rect 34977 10217 34989 10220
rect 35023 10217 35035 10251
rect 34977 10211 35035 10217
rect 35434 10208 35440 10260
rect 35492 10208 35498 10260
rect 32398 10140 32404 10192
rect 32456 10180 32462 10192
rect 32456 10152 34008 10180
rect 32456 10140 32462 10152
rect 33689 10115 33747 10121
rect 33689 10112 33701 10115
rect 31435 10084 32076 10112
rect 32324 10084 33701 10112
rect 31435 10081 31447 10084
rect 31389 10075 31447 10081
rect 30285 10047 30343 10053
rect 30285 10013 30297 10047
rect 30331 10013 30343 10047
rect 30285 10007 30343 10013
rect 30469 10047 30527 10053
rect 30469 10013 30481 10047
rect 30515 10044 30527 10047
rect 30745 10047 30803 10053
rect 30745 10044 30757 10047
rect 30515 10016 30757 10044
rect 30515 10013 30527 10016
rect 30469 10007 30527 10013
rect 30745 10013 30757 10016
rect 30791 10013 30803 10047
rect 30745 10007 30803 10013
rect 31665 10047 31723 10053
rect 31665 10013 31677 10047
rect 31711 10013 31723 10047
rect 31665 10007 31723 10013
rect 16448 9948 16882 9976
rect 18340 9948 20024 9976
rect 16448 9936 16454 9948
rect 21542 9936 21548 9988
rect 21600 9936 21606 9988
rect 25958 9976 25964 9988
rect 25898 9948 25964 9976
rect 25958 9936 25964 9948
rect 26016 9936 26022 9988
rect 30101 9979 30159 9985
rect 30101 9945 30113 9979
rect 30147 9976 30159 9979
rect 30374 9976 30380 9988
rect 30147 9948 30380 9976
rect 30147 9945 30159 9948
rect 30101 9939 30159 9945
rect 30374 9936 30380 9948
rect 30432 9936 30438 9988
rect 31680 9976 31708 10007
rect 31846 10004 31852 10056
rect 31904 10004 31910 10056
rect 32048 10053 32076 10084
rect 33689 10081 33701 10084
rect 33735 10081 33747 10115
rect 33689 10075 33747 10081
rect 32033 10047 32091 10053
rect 32033 10013 32045 10047
rect 32079 10013 32091 10047
rect 32033 10007 32091 10013
rect 32122 10004 32128 10056
rect 32180 10046 32186 10056
rect 32217 10047 32275 10053
rect 32217 10046 32229 10047
rect 32180 10018 32229 10046
rect 32180 10004 32186 10018
rect 32217 10013 32229 10018
rect 32263 10044 32275 10047
rect 32263 10016 32444 10044
rect 32263 10013 32275 10016
rect 32217 10007 32275 10013
rect 32306 9976 32312 9988
rect 31680 9948 32312 9976
rect 32306 9936 32312 9948
rect 32364 9936 32370 9988
rect 32416 9976 32444 10016
rect 32490 10004 32496 10056
rect 32548 10004 32554 10056
rect 32674 10004 32680 10056
rect 32732 10004 32738 10056
rect 33980 10053 34008 10152
rect 34422 10072 34428 10124
rect 34480 10112 34486 10124
rect 34480 10084 35388 10112
rect 34480 10072 34486 10084
rect 33965 10047 34023 10053
rect 33965 10013 33977 10047
rect 34011 10013 34023 10047
rect 33965 10007 34023 10013
rect 34698 10004 34704 10056
rect 34756 10004 34762 10056
rect 34790 10004 34796 10056
rect 34848 10004 34854 10056
rect 35360 10053 35388 10084
rect 35345 10047 35403 10053
rect 35345 10013 35357 10047
rect 35391 10013 35403 10047
rect 35345 10007 35403 10013
rect 35529 10047 35587 10053
rect 35529 10013 35541 10047
rect 35575 10013 35587 10047
rect 35529 10007 35587 10013
rect 33873 9979 33931 9985
rect 33873 9976 33885 9979
rect 32416 9948 33885 9976
rect 33873 9945 33885 9948
rect 33919 9945 33931 9979
rect 33873 9939 33931 9945
rect 34606 9936 34612 9988
rect 34664 9976 34670 9988
rect 35544 9976 35572 10007
rect 34664 9948 35572 9976
rect 34664 9936 34670 9948
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 25976 9908 26004 9936
rect 25004 9880 26004 9908
rect 25004 9868 25010 9880
rect 29822 9868 29828 9920
rect 29880 9868 29886 9920
rect 31573 9911 31631 9917
rect 31573 9877 31585 9911
rect 31619 9908 31631 9911
rect 33778 9908 33784 9920
rect 31619 9880 33784 9908
rect 31619 9877 31631 9880
rect 31573 9871 31631 9877
rect 33778 9868 33784 9880
rect 33836 9868 33842 9920
rect 34054 9868 34060 9920
rect 34112 9868 34118 9920
rect 34238 9868 34244 9920
rect 34296 9868 34302 9920
rect 1104 9818 37076 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 37076 9818
rect 1104 9744 37076 9766
rect 15381 9707 15439 9713
rect 15381 9673 15393 9707
rect 15427 9704 15439 9707
rect 15470 9704 15476 9716
rect 15427 9676 15476 9704
rect 15427 9673 15439 9676
rect 15381 9667 15439 9673
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 18233 9707 18291 9713
rect 18233 9673 18245 9707
rect 18279 9704 18291 9707
rect 18414 9704 18420 9716
rect 18279 9676 18420 9704
rect 18279 9673 18291 9676
rect 18233 9667 18291 9673
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 19978 9704 19984 9716
rect 19628 9676 19984 9704
rect 13906 9596 13912 9648
rect 13964 9596 13970 9648
rect 16390 9636 16396 9648
rect 15134 9608 16396 9636
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 17862 9636 17868 9648
rect 17512 9608 17868 9636
rect 13630 9528 13636 9580
rect 13688 9528 13694 9580
rect 16482 9528 16488 9580
rect 16540 9528 16546 9580
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 17512 9577 17540 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 18141 9639 18199 9645
rect 18141 9636 18153 9639
rect 18104 9608 18153 9636
rect 18104 9596 18110 9608
rect 18141 9605 18153 9608
rect 18187 9605 18199 9639
rect 19628 9636 19656 9676
rect 19978 9664 19984 9676
rect 20036 9704 20042 9716
rect 20622 9704 20628 9716
rect 20036 9676 20628 9704
rect 20036 9664 20042 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 23124 9676 23428 9704
rect 19274 9608 19656 9636
rect 19705 9639 19763 9645
rect 18141 9599 18199 9605
rect 19705 9605 19717 9639
rect 19751 9636 19763 9639
rect 20714 9636 20720 9648
rect 19751 9608 20720 9636
rect 19751 9605 19763 9608
rect 19705 9599 19763 9605
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 23124 9636 23152 9676
rect 23400 9648 23428 9676
rect 26142 9664 26148 9716
rect 26200 9664 26206 9716
rect 28626 9664 28632 9716
rect 28684 9704 28690 9716
rect 28721 9707 28779 9713
rect 28721 9704 28733 9707
rect 28684 9676 28733 9704
rect 28684 9664 28690 9676
rect 28721 9673 28733 9676
rect 28767 9673 28779 9707
rect 28721 9667 28779 9673
rect 22862 9608 23152 9636
rect 23198 9596 23204 9648
rect 23256 9636 23262 9648
rect 23293 9639 23351 9645
rect 23293 9636 23305 9639
rect 23256 9608 23305 9636
rect 23256 9596 23262 9608
rect 23293 9605 23305 9608
rect 23339 9605 23351 9639
rect 23293 9599 23351 9605
rect 23382 9596 23388 9648
rect 23440 9636 23446 9648
rect 24946 9636 24952 9648
rect 23440 9608 24952 9636
rect 23440 9596 23446 9608
rect 24946 9596 24952 9608
rect 25004 9636 25010 9648
rect 25130 9636 25136 9648
rect 25004 9608 25136 9636
rect 25004 9596 25010 9608
rect 25130 9596 25136 9608
rect 25188 9596 25194 9648
rect 26234 9596 26240 9648
rect 26292 9636 26298 9648
rect 26513 9639 26571 9645
rect 26513 9636 26525 9639
rect 26292 9608 26525 9636
rect 26292 9596 26298 9608
rect 26513 9605 26525 9608
rect 26559 9605 26571 9639
rect 26513 9599 26571 9605
rect 26694 9596 26700 9648
rect 26752 9596 26758 9648
rect 26786 9596 26792 9648
rect 26844 9636 26850 9648
rect 27249 9639 27307 9645
rect 27249 9636 27261 9639
rect 26844 9608 27261 9636
rect 26844 9596 26850 9608
rect 27249 9605 27261 9608
rect 27295 9605 27307 9639
rect 28736 9636 28764 9667
rect 30190 9664 30196 9716
rect 30248 9704 30254 9716
rect 32490 9704 32496 9716
rect 30248 9676 32496 9704
rect 30248 9664 30254 9676
rect 32490 9664 32496 9676
rect 32548 9664 32554 9716
rect 32674 9664 32680 9716
rect 32732 9704 32738 9716
rect 33781 9707 33839 9713
rect 32732 9676 33456 9704
rect 32732 9664 32738 9676
rect 33428 9648 33456 9676
rect 33781 9673 33793 9707
rect 33827 9704 33839 9707
rect 33827 9676 35020 9704
rect 33827 9673 33839 9676
rect 33781 9667 33839 9673
rect 29273 9639 29331 9645
rect 29273 9636 29285 9639
rect 28736 9608 29285 9636
rect 27249 9599 27307 9605
rect 29273 9605 29285 9608
rect 29319 9605 29331 9639
rect 29273 9599 29331 9605
rect 31757 9639 31815 9645
rect 31757 9605 31769 9639
rect 31803 9636 31815 9639
rect 32030 9636 32036 9648
rect 31803 9608 32036 9636
rect 31803 9605 31815 9608
rect 31757 9599 31815 9605
rect 32030 9596 32036 9608
rect 32088 9596 32094 9648
rect 32306 9596 32312 9648
rect 32364 9596 32370 9648
rect 33410 9596 33416 9648
rect 33468 9596 33474 9648
rect 34393 9639 34451 9645
rect 34393 9636 34405 9639
rect 33520 9608 34405 9636
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9537 17555 9571
rect 17497 9531 17555 9537
rect 17681 9571 17739 9577
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 13648 9500 13676 9528
rect 15657 9503 15715 9509
rect 15657 9500 15669 9503
rect 13648 9472 15669 9500
rect 15657 9469 15669 9472
rect 15703 9500 15715 9503
rect 16114 9500 16120 9512
rect 15703 9472 16120 9500
rect 15703 9469 15715 9472
rect 15657 9463 15715 9469
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 17696 9500 17724 9531
rect 21266 9528 21272 9580
rect 21324 9528 21330 9580
rect 23566 9528 23572 9580
rect 23624 9568 23630 9580
rect 23661 9571 23719 9577
rect 23661 9568 23673 9571
rect 23624 9540 23673 9568
rect 23624 9528 23630 9540
rect 23661 9537 23673 9540
rect 23707 9568 23719 9571
rect 24397 9571 24455 9577
rect 24397 9568 24409 9571
rect 23707 9540 24409 9568
rect 23707 9537 23719 9540
rect 23661 9531 23719 9537
rect 24397 9537 24409 9540
rect 24443 9537 24455 9571
rect 24397 9531 24455 9537
rect 28350 9528 28356 9580
rect 28408 9528 28414 9580
rect 28718 9528 28724 9580
rect 28776 9568 28782 9580
rect 29181 9571 29239 9577
rect 29181 9568 29193 9571
rect 28776 9540 29193 9568
rect 28776 9528 28782 9540
rect 29181 9537 29193 9540
rect 29227 9537 29239 9571
rect 29181 9531 29239 9537
rect 29822 9528 29828 9580
rect 29880 9528 29886 9580
rect 30009 9571 30067 9577
rect 30009 9537 30021 9571
rect 30055 9537 30067 9571
rect 30009 9531 30067 9537
rect 17862 9500 17868 9512
rect 17696 9472 17868 9500
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 19981 9503 20039 9509
rect 19981 9500 19993 9503
rect 19904 9472 19993 9500
rect 16132 9432 16160 9460
rect 17218 9432 17224 9444
rect 16132 9404 17224 9432
rect 17218 9392 17224 9404
rect 17276 9432 17282 9444
rect 17276 9404 18736 9432
rect 17276 9392 17282 9404
rect 18708 9364 18736 9404
rect 19904 9364 19932 9472
rect 19981 9469 19993 9472
rect 20027 9469 20039 9503
rect 19981 9463 20039 9469
rect 20070 9460 20076 9512
rect 20128 9500 20134 9512
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 20128 9472 20269 9500
rect 20128 9460 20134 9472
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 21821 9503 21879 9509
rect 21821 9469 21833 9503
rect 21867 9500 21879 9503
rect 22278 9500 22284 9512
rect 21867 9472 22284 9500
rect 21867 9469 21879 9472
rect 21821 9463 21879 9469
rect 22278 9460 22284 9472
rect 22336 9460 22342 9512
rect 24670 9460 24676 9512
rect 24728 9460 24734 9512
rect 26970 9460 26976 9512
rect 27028 9460 27034 9512
rect 29270 9460 29276 9512
rect 29328 9500 29334 9512
rect 29457 9503 29515 9509
rect 29457 9500 29469 9503
rect 29328 9472 29469 9500
rect 29328 9460 29334 9472
rect 29457 9469 29469 9472
rect 29503 9500 29515 9503
rect 29546 9500 29552 9512
rect 29503 9472 29552 9500
rect 29503 9469 29515 9472
rect 29457 9463 29515 9469
rect 29546 9460 29552 9472
rect 29604 9460 29610 9512
rect 29641 9503 29699 9509
rect 29641 9469 29653 9503
rect 29687 9500 29699 9503
rect 29730 9500 29736 9512
rect 29687 9472 29736 9500
rect 29687 9469 29699 9472
rect 29641 9463 29699 9469
rect 29730 9460 29736 9472
rect 29788 9460 29794 9512
rect 30024 9432 30052 9531
rect 30282 9528 30288 9580
rect 30340 9528 30346 9580
rect 30742 9528 30748 9580
rect 30800 9568 30806 9580
rect 30837 9571 30895 9577
rect 30837 9568 30849 9571
rect 30800 9540 30849 9568
rect 30800 9528 30806 9540
rect 30837 9537 30849 9540
rect 30883 9537 30895 9571
rect 30837 9531 30895 9537
rect 31113 9571 31171 9577
rect 31113 9537 31125 9571
rect 31159 9568 31171 9571
rect 31294 9568 31300 9580
rect 31159 9540 31300 9568
rect 31159 9537 31171 9540
rect 31113 9531 31171 9537
rect 30653 9503 30711 9509
rect 30653 9469 30665 9503
rect 30699 9500 30711 9503
rect 31128 9500 31156 9531
rect 31294 9528 31300 9540
rect 31352 9528 31358 9580
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9537 32551 9571
rect 32493 9531 32551 9537
rect 30699 9472 31156 9500
rect 32508 9500 32536 9531
rect 32674 9528 32680 9580
rect 32732 9528 32738 9580
rect 32766 9528 32772 9580
rect 32824 9568 32830 9580
rect 33520 9568 33548 9608
rect 34393 9605 34405 9608
rect 34439 9605 34451 9639
rect 34393 9599 34451 9605
rect 34606 9596 34612 9648
rect 34664 9596 34670 9648
rect 32824 9540 33548 9568
rect 32824 9528 32830 9540
rect 33686 9528 33692 9580
rect 33744 9528 33750 9580
rect 33965 9571 34023 9577
rect 33965 9537 33977 9571
rect 34011 9568 34023 9571
rect 34238 9568 34244 9580
rect 34011 9540 34244 9568
rect 34011 9537 34023 9540
rect 33965 9531 34023 9537
rect 33980 9500 34008 9531
rect 34238 9528 34244 9540
rect 34296 9568 34302 9580
rect 34992 9577 35020 9676
rect 34701 9571 34759 9577
rect 34701 9568 34713 9571
rect 34296 9540 34713 9568
rect 34296 9528 34302 9540
rect 34701 9537 34713 9540
rect 34747 9537 34759 9571
rect 34701 9531 34759 9537
rect 34977 9571 35035 9577
rect 34977 9537 34989 9571
rect 35023 9568 35035 9571
rect 35342 9568 35348 9580
rect 35023 9540 35348 9568
rect 35023 9537 35035 9540
rect 34977 9531 35035 9537
rect 35342 9528 35348 9540
rect 35400 9528 35406 9580
rect 32508 9472 34008 9500
rect 34149 9503 34207 9509
rect 30699 9469 30711 9472
rect 30653 9463 30711 9469
rect 34149 9469 34161 9503
rect 34195 9500 34207 9503
rect 34790 9500 34796 9512
rect 34195 9472 34796 9500
rect 34195 9469 34207 9472
rect 34149 9463 34207 9469
rect 34790 9460 34796 9472
rect 34848 9460 34854 9512
rect 33042 9432 33048 9444
rect 30024 9404 33048 9432
rect 33042 9392 33048 9404
rect 33100 9392 33106 9444
rect 33778 9392 33784 9444
rect 33836 9432 33842 9444
rect 33836 9404 34468 9432
rect 33836 9392 33842 9404
rect 18708 9336 19932 9364
rect 28810 9324 28816 9376
rect 28868 9324 28874 9376
rect 33134 9324 33140 9376
rect 33192 9364 33198 9376
rect 34054 9364 34060 9376
rect 33192 9336 34060 9364
rect 33192 9324 33198 9336
rect 34054 9324 34060 9336
rect 34112 9324 34118 9376
rect 34238 9324 34244 9376
rect 34296 9324 34302 9376
rect 34440 9373 34468 9404
rect 34425 9367 34483 9373
rect 34425 9333 34437 9367
rect 34471 9333 34483 9367
rect 34425 9327 34483 9333
rect 34698 9324 34704 9376
rect 34756 9364 34762 9376
rect 34793 9367 34851 9373
rect 34793 9364 34805 9367
rect 34756 9336 34805 9364
rect 34756 9324 34762 9336
rect 34793 9333 34805 9336
rect 34839 9333 34851 9367
rect 34793 9327 34851 9333
rect 1104 9274 37076 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 37076 9274
rect 1104 9200 37076 9222
rect 23658 9120 23664 9172
rect 23716 9120 23722 9172
rect 24670 9120 24676 9172
rect 24728 9160 24734 9172
rect 25501 9163 25559 9169
rect 25501 9160 25513 9163
rect 24728 9132 25513 9160
rect 24728 9120 24734 9132
rect 25501 9129 25513 9132
rect 25547 9129 25559 9163
rect 25501 9123 25559 9129
rect 26694 9120 26700 9172
rect 26752 9160 26758 9172
rect 26752 9132 28672 9160
rect 26752 9120 26758 9132
rect 28644 9092 28672 9132
rect 28718 9120 28724 9172
rect 28776 9120 28782 9172
rect 29181 9163 29239 9169
rect 29181 9129 29193 9163
rect 29227 9129 29239 9163
rect 29181 9123 29239 9129
rect 29365 9163 29423 9169
rect 29365 9129 29377 9163
rect 29411 9160 29423 9163
rect 29638 9160 29644 9172
rect 29411 9132 29644 9160
rect 29411 9129 29423 9132
rect 29365 9123 29423 9129
rect 29196 9092 29224 9123
rect 29638 9120 29644 9132
rect 29696 9120 29702 9172
rect 31205 9163 31263 9169
rect 31205 9129 31217 9163
rect 31251 9160 31263 9163
rect 31478 9160 31484 9172
rect 31251 9132 31484 9160
rect 31251 9129 31263 9132
rect 31205 9123 31263 9129
rect 31478 9120 31484 9132
rect 31536 9120 31542 9172
rect 31941 9163 31999 9169
rect 31941 9129 31953 9163
rect 31987 9160 31999 9163
rect 32766 9160 32772 9172
rect 31987 9132 32772 9160
rect 31987 9129 31999 9132
rect 31941 9123 31999 9129
rect 32766 9120 32772 9132
rect 32824 9120 32830 9172
rect 33523 9163 33581 9169
rect 33523 9129 33535 9163
rect 33569 9160 33581 9163
rect 34238 9160 34244 9172
rect 33569 9132 34244 9160
rect 33569 9129 33581 9132
rect 33523 9123 33581 9129
rect 34238 9120 34244 9132
rect 34296 9120 34302 9172
rect 30190 9092 30196 9104
rect 28644 9064 29132 9092
rect 29196 9064 30196 9092
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 16025 9027 16083 9033
rect 16025 9024 16037 9027
rect 14332 8996 16037 9024
rect 14332 8984 14338 8996
rect 16025 8993 16037 8996
rect 16071 9024 16083 9027
rect 16666 9024 16672 9036
rect 16071 8996 16672 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 19705 9027 19763 9033
rect 19705 9024 19717 9027
rect 18524 8996 19717 9024
rect 15197 8959 15255 8965
rect 15197 8925 15209 8959
rect 15243 8956 15255 8959
rect 15286 8956 15292 8968
rect 15243 8928 15292 8956
rect 15243 8925 15255 8928
rect 15197 8919 15255 8925
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 15378 8916 15384 8968
rect 15436 8916 15442 8968
rect 15470 8916 15476 8968
rect 15528 8916 15534 8968
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18524 8965 18552 8996
rect 19705 8993 19717 8996
rect 19751 9024 19763 9027
rect 20438 9024 20444 9036
rect 19751 8996 20444 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 20438 8984 20444 8996
rect 20496 8984 20502 9036
rect 21910 8984 21916 9036
rect 21968 8984 21974 9036
rect 22189 9027 22247 9033
rect 22189 8993 22201 9027
rect 22235 9024 22247 9027
rect 22922 9024 22928 9036
rect 22235 8996 22928 9024
rect 22235 8993 22247 8996
rect 22189 8987 22247 8993
rect 22922 8984 22928 8996
rect 22980 8984 22986 9036
rect 23382 8984 23388 9036
rect 23440 8984 23446 9036
rect 23566 8984 23572 9036
rect 23624 9024 23630 9036
rect 23624 8996 25084 9024
rect 23624 8984 23630 8996
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18288 8928 18337 8956
rect 18288 8916 18294 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 18601 8959 18659 8965
rect 18601 8925 18613 8959
rect 18647 8956 18659 8959
rect 18690 8956 18696 8968
rect 18647 8928 18696 8956
rect 18647 8925 18659 8928
rect 18601 8919 18659 8925
rect 14090 8848 14096 8900
rect 14148 8888 14154 8900
rect 14737 8891 14795 8897
rect 14737 8888 14749 8891
rect 14148 8860 14749 8888
rect 14148 8848 14154 8860
rect 14737 8857 14749 8860
rect 14783 8857 14795 8891
rect 15304 8888 15332 8916
rect 15930 8888 15936 8900
rect 15304 8860 15936 8888
rect 14737 8851 14795 8857
rect 15930 8848 15936 8860
rect 15988 8888 15994 8900
rect 16206 8888 16212 8900
rect 15988 8860 16212 8888
rect 15988 8848 15994 8860
rect 16206 8848 16212 8860
rect 16264 8848 16270 8900
rect 16301 8891 16359 8897
rect 16301 8857 16313 8891
rect 16347 8857 16359 8891
rect 16301 8851 16359 8857
rect 16316 8820 16344 8851
rect 16390 8848 16396 8900
rect 16448 8888 16454 8900
rect 17865 8891 17923 8897
rect 17865 8888 17877 8891
rect 16448 8860 16790 8888
rect 17604 8860 17877 8888
rect 16448 8848 16454 8860
rect 17604 8820 17632 8860
rect 17865 8857 17877 8860
rect 17911 8857 17923 8891
rect 17865 8851 17923 8857
rect 16316 8792 17632 8820
rect 17773 8823 17831 8829
rect 17773 8789 17785 8823
rect 17819 8820 17831 8823
rect 18616 8820 18644 8919
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 21450 8916 21456 8968
rect 21508 8916 21514 8968
rect 23400 8956 23428 8984
rect 23322 8928 23428 8956
rect 23842 8916 23848 8968
rect 23900 8956 23906 8968
rect 24854 8956 24860 8968
rect 23900 8928 24860 8956
rect 23900 8916 23906 8928
rect 24854 8916 24860 8928
rect 24912 8916 24918 8968
rect 25056 8965 25084 8996
rect 26050 8984 26056 9036
rect 26108 8984 26114 9036
rect 26970 8984 26976 9036
rect 27028 8984 27034 9036
rect 27249 9027 27307 9033
rect 27249 8993 27261 9027
rect 27295 9024 27307 9027
rect 28810 9024 28816 9036
rect 27295 8996 28816 9024
rect 27295 8993 27307 8996
rect 27249 8987 27307 8993
rect 28810 8984 28816 8996
rect 28868 8984 28874 9036
rect 25041 8959 25099 8965
rect 25041 8925 25053 8959
rect 25087 8925 25099 8959
rect 25041 8919 25099 8925
rect 25133 8959 25191 8965
rect 25133 8925 25145 8959
rect 25179 8956 25191 8959
rect 25590 8956 25596 8968
rect 25179 8928 25596 8956
rect 25179 8925 25191 8928
rect 25133 8919 25191 8925
rect 25590 8916 25596 8928
rect 25648 8916 25654 8968
rect 25869 8959 25927 8965
rect 25869 8925 25881 8959
rect 25915 8956 25927 8959
rect 26142 8956 26148 8968
rect 25915 8928 26148 8956
rect 25915 8925 25927 8928
rect 25869 8919 25927 8925
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 26881 8959 26939 8965
rect 26881 8925 26893 8959
rect 26927 8925 26939 8959
rect 26881 8919 26939 8925
rect 20622 8848 20628 8900
rect 20680 8848 20686 8900
rect 21174 8848 21180 8900
rect 21232 8848 21238 8900
rect 24397 8891 24455 8897
rect 24397 8857 24409 8891
rect 24443 8888 24455 8891
rect 24578 8888 24584 8900
rect 24443 8860 24584 8888
rect 24443 8857 24455 8860
rect 24397 8851 24455 8857
rect 24578 8848 24584 8860
rect 24636 8848 24642 8900
rect 17819 8792 18644 8820
rect 17819 8789 17831 8792
rect 17773 8783 17831 8789
rect 25958 8780 25964 8832
rect 26016 8780 26022 8832
rect 26896 8820 26924 8919
rect 28350 8916 28356 8968
rect 28408 8916 28414 8968
rect 29104 8956 29132 9064
rect 30190 9052 30196 9064
rect 30248 9052 30254 9104
rect 29546 8984 29552 9036
rect 29604 9024 29610 9036
rect 29733 9027 29791 9033
rect 29733 9024 29745 9027
rect 29604 8996 29745 9024
rect 29604 8984 29610 8996
rect 29733 8993 29745 8996
rect 29779 8993 29791 9027
rect 29733 8987 29791 8993
rect 31297 9027 31355 9033
rect 31297 8993 31309 9027
rect 31343 9024 31355 9027
rect 31386 9024 31392 9036
rect 31343 8996 31392 9024
rect 31343 8993 31355 8996
rect 31297 8987 31355 8993
rect 31386 8984 31392 8996
rect 31444 8984 31450 9036
rect 31662 8984 31668 9036
rect 31720 8984 31726 9036
rect 31757 9027 31815 9033
rect 31757 8993 31769 9027
rect 31803 9024 31815 9027
rect 32033 9027 32091 9033
rect 32033 9024 32045 9027
rect 31803 8996 32045 9024
rect 31803 8993 31815 8996
rect 31757 8987 31815 8993
rect 32033 8993 32045 8996
rect 32079 9024 32091 9027
rect 33134 9024 33140 9036
rect 32079 8996 33140 9024
rect 32079 8993 32091 8996
rect 32033 8987 32091 8993
rect 33134 8984 33140 8996
rect 33192 8984 33198 9036
rect 33410 8984 33416 9036
rect 33468 9024 33474 9036
rect 33781 9027 33839 9033
rect 33781 9024 33793 9027
rect 33468 8996 33793 9024
rect 33468 8984 33474 8996
rect 33781 8993 33793 8996
rect 33827 8993 33839 9027
rect 33781 8987 33839 8993
rect 34606 8984 34612 9036
rect 34664 9024 34670 9036
rect 34701 9027 34759 9033
rect 34701 9024 34713 9027
rect 34664 8996 34713 9024
rect 34664 8984 34670 8996
rect 34701 8993 34713 8996
rect 34747 8993 34759 9027
rect 34701 8987 34759 8993
rect 30377 8959 30435 8965
rect 30377 8956 30389 8959
rect 29104 8928 30389 8956
rect 30377 8925 30389 8928
rect 30423 8925 30435 8959
rect 30377 8919 30435 8925
rect 28997 8891 29055 8897
rect 28997 8857 29009 8891
rect 29043 8888 29055 8891
rect 29454 8888 29460 8900
rect 29043 8860 29460 8888
rect 29043 8857 29055 8860
rect 28997 8851 29055 8857
rect 29454 8848 29460 8860
rect 29512 8848 29518 8900
rect 30392 8888 30420 8919
rect 30466 8916 30472 8968
rect 30524 8956 30530 8968
rect 31021 8959 31079 8965
rect 31021 8956 31033 8959
rect 30524 8928 31033 8956
rect 30524 8916 30530 8928
rect 31021 8925 31033 8928
rect 31067 8956 31079 8959
rect 31202 8956 31208 8968
rect 31067 8928 31208 8956
rect 31067 8925 31079 8928
rect 31021 8919 31079 8925
rect 31202 8916 31208 8928
rect 31260 8916 31266 8968
rect 31527 8959 31585 8965
rect 31527 8925 31539 8959
rect 31573 8956 31585 8959
rect 32122 8956 32128 8968
rect 31573 8928 32128 8956
rect 31573 8925 31585 8928
rect 31527 8919 31585 8925
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 34054 8916 34060 8968
rect 34112 8956 34118 8968
rect 34241 8959 34299 8965
rect 34241 8956 34253 8959
rect 34112 8928 34253 8956
rect 34112 8916 34118 8928
rect 34241 8925 34253 8928
rect 34287 8925 34299 8959
rect 34241 8919 34299 8925
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 34885 8959 34943 8965
rect 34885 8956 34897 8959
rect 34848 8928 34897 8956
rect 34848 8916 34854 8928
rect 34885 8925 34897 8928
rect 34931 8925 34943 8959
rect 34885 8919 34943 8925
rect 34974 8916 34980 8968
rect 35032 8916 35038 8968
rect 30558 8888 30564 8900
rect 30392 8860 30564 8888
rect 30558 8848 30564 8860
rect 30616 8848 30622 8900
rect 30650 8848 30656 8900
rect 30708 8848 30714 8900
rect 30929 8891 30987 8897
rect 30929 8888 30941 8891
rect 30760 8860 30941 8888
rect 27614 8820 27620 8832
rect 26896 8792 27620 8820
rect 27614 8780 27620 8792
rect 27672 8780 27678 8832
rect 29207 8823 29265 8829
rect 29207 8789 29219 8823
rect 29253 8820 29265 8823
rect 30760 8820 30788 8860
rect 30929 8857 30941 8860
rect 30975 8888 30987 8891
rect 31294 8888 31300 8900
rect 30975 8860 31300 8888
rect 30975 8857 30987 8860
rect 30929 8851 30987 8857
rect 31294 8848 31300 8860
rect 31352 8848 31358 8900
rect 31389 8891 31447 8897
rect 31389 8857 31401 8891
rect 31435 8888 31447 8891
rect 33594 8888 33600 8900
rect 31435 8860 31708 8888
rect 33074 8860 33600 8888
rect 31435 8857 31447 8860
rect 31389 8851 31447 8857
rect 29253 8792 30788 8820
rect 29253 8789 29265 8792
rect 29207 8783 29265 8789
rect 30834 8780 30840 8832
rect 30892 8820 30898 8832
rect 31570 8820 31576 8832
rect 30892 8792 31576 8820
rect 30892 8780 30898 8792
rect 31570 8780 31576 8792
rect 31628 8780 31634 8832
rect 31680 8820 31708 8860
rect 33594 8848 33600 8860
rect 33652 8848 33658 8900
rect 33873 8891 33931 8897
rect 33873 8857 33885 8891
rect 33919 8857 33931 8891
rect 33873 8851 33931 8857
rect 34425 8891 34483 8897
rect 34425 8857 34437 8891
rect 34471 8888 34483 8891
rect 35986 8888 35992 8900
rect 34471 8860 35992 8888
rect 34471 8857 34483 8860
rect 34425 8851 34483 8857
rect 33410 8820 33416 8832
rect 31680 8792 33416 8820
rect 33410 8780 33416 8792
rect 33468 8820 33474 8832
rect 33888 8820 33916 8851
rect 35986 8848 35992 8860
rect 36044 8888 36050 8900
rect 36446 8888 36452 8900
rect 36044 8860 36452 8888
rect 36044 8848 36050 8860
rect 36446 8848 36452 8860
rect 36504 8848 36510 8900
rect 33468 8792 33916 8820
rect 33468 8780 33474 8792
rect 34238 8780 34244 8832
rect 34296 8820 34302 8832
rect 34701 8823 34759 8829
rect 34701 8820 34713 8823
rect 34296 8792 34713 8820
rect 34296 8780 34302 8792
rect 34701 8789 34713 8792
rect 34747 8789 34759 8823
rect 34701 8783 34759 8789
rect 1104 8730 37076 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 37076 8730
rect 1104 8656 37076 8678
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 15565 8619 15623 8625
rect 15565 8616 15577 8619
rect 15528 8588 15577 8616
rect 15528 8576 15534 8588
rect 15565 8585 15577 8588
rect 15611 8585 15623 8619
rect 15565 8579 15623 8585
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 18690 8616 18696 8628
rect 16264 8588 18696 8616
rect 16264 8576 16270 8588
rect 18690 8576 18696 8588
rect 18748 8616 18754 8628
rect 19794 8616 19800 8628
rect 18748 8588 19800 8616
rect 18748 8576 18754 8588
rect 19794 8576 19800 8588
rect 19852 8576 19858 8628
rect 27982 8576 27988 8628
rect 28040 8616 28046 8628
rect 28040 8588 32720 8616
rect 28040 8576 28046 8588
rect 14090 8508 14096 8560
rect 14148 8508 14154 8560
rect 15654 8548 15660 8560
rect 15318 8520 15660 8548
rect 15654 8508 15660 8520
rect 15712 8548 15718 8560
rect 16390 8548 16396 8560
rect 15712 8520 16396 8548
rect 15712 8508 15718 8520
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 17589 8551 17647 8557
rect 17589 8548 17601 8551
rect 16540 8520 17601 8548
rect 16540 8508 16546 8520
rect 17589 8517 17601 8520
rect 17635 8548 17647 8551
rect 23014 8548 23020 8560
rect 17635 8520 23020 8548
rect 17635 8517 17647 8520
rect 17589 8511 17647 8517
rect 23014 8508 23020 8520
rect 23072 8508 23078 8560
rect 24026 8508 24032 8560
rect 24084 8548 24090 8560
rect 25593 8551 25651 8557
rect 25593 8548 25605 8551
rect 24084 8520 25605 8548
rect 24084 8508 24090 8520
rect 25593 8517 25605 8520
rect 25639 8517 25651 8551
rect 25593 8511 25651 8517
rect 26694 8508 26700 8560
rect 26752 8548 26758 8560
rect 27157 8551 27215 8557
rect 27157 8548 27169 8551
rect 26752 8520 27169 8548
rect 26752 8508 26758 8520
rect 27157 8517 27169 8520
rect 27203 8517 27215 8551
rect 27157 8511 27215 8517
rect 27614 8508 27620 8560
rect 27672 8508 27678 8560
rect 28460 8557 28488 8588
rect 32692 8560 32720 8588
rect 33686 8576 33692 8628
rect 33744 8616 33750 8628
rect 33744 8588 34360 8616
rect 33744 8576 33750 8588
rect 28445 8551 28503 8557
rect 28445 8517 28457 8551
rect 28491 8517 28503 8551
rect 28445 8511 28503 8517
rect 28718 8508 28724 8560
rect 28776 8548 28782 8560
rect 28997 8551 29055 8557
rect 28997 8548 29009 8551
rect 28776 8520 29009 8548
rect 28776 8508 28782 8520
rect 28997 8517 29009 8520
rect 29043 8517 29055 8551
rect 28997 8511 29055 8517
rect 29730 8508 29736 8560
rect 29788 8548 29794 8560
rect 29825 8551 29883 8557
rect 29825 8548 29837 8551
rect 29788 8520 29837 8548
rect 29788 8508 29794 8520
rect 29825 8517 29837 8520
rect 29871 8517 29883 8551
rect 29825 8511 29883 8517
rect 31202 8508 31208 8560
rect 31260 8548 31266 8560
rect 31541 8551 31599 8557
rect 31541 8548 31553 8551
rect 31260 8520 31553 8548
rect 31260 8508 31266 8520
rect 31541 8517 31553 8520
rect 31587 8517 31599 8551
rect 31541 8511 31599 8517
rect 31662 8508 31668 8560
rect 31720 8548 31726 8560
rect 31757 8551 31815 8557
rect 31757 8548 31769 8551
rect 31720 8520 31769 8548
rect 31720 8508 31726 8520
rect 31757 8517 31769 8520
rect 31803 8517 31815 8551
rect 31757 8511 31815 8517
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18598 8480 18604 8492
rect 18555 8452 18604 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 18690 8440 18696 8492
rect 18748 8440 18754 8492
rect 20438 8440 20444 8492
rect 20496 8440 20502 8492
rect 20530 8440 20536 8492
rect 20588 8440 20594 8492
rect 20717 8483 20775 8489
rect 20717 8480 20729 8483
rect 20640 8452 20729 8480
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8412 13875 8415
rect 13863 8384 13952 8412
rect 13863 8381 13875 8384
rect 13817 8375 13875 8381
rect 13924 8276 13952 8384
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 16724 8384 16773 8412
rect 16724 8372 16730 8384
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 18408 8415 18466 8421
rect 18408 8412 18420 8415
rect 16761 8375 16819 8381
rect 18340 8384 18420 8412
rect 18340 8356 18368 8384
rect 18408 8381 18420 8384
rect 18454 8381 18466 8415
rect 18408 8375 18466 8381
rect 18782 8372 18788 8424
rect 18840 8412 18846 8424
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 18840 8384 19165 8412
rect 18840 8372 18846 8384
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19153 8375 19211 8381
rect 19794 8372 19800 8424
rect 19852 8412 19858 8424
rect 20640 8412 20668 8452
rect 20717 8449 20729 8452
rect 20763 8449 20775 8483
rect 20717 8443 20775 8449
rect 21174 8440 21180 8492
rect 21232 8440 21238 8492
rect 23750 8440 23756 8492
rect 23808 8440 23814 8492
rect 23842 8440 23848 8492
rect 23900 8480 23906 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23900 8452 23949 8480
rect 23900 8440 23906 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 26789 8483 26847 8489
rect 26789 8449 26801 8483
rect 26835 8480 26847 8483
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26835 8452 26985 8480
rect 26835 8449 26847 8452
rect 26789 8443 26847 8449
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27890 8440 27896 8492
rect 27948 8480 27954 8492
rect 28905 8483 28963 8489
rect 28905 8480 28917 8483
rect 27948 8452 28917 8480
rect 27948 8440 27954 8452
rect 28905 8449 28917 8452
rect 28951 8449 28963 8483
rect 31772 8480 31800 8511
rect 32674 8508 32680 8560
rect 32732 8548 32738 8560
rect 33045 8551 33103 8557
rect 33045 8548 33057 8551
rect 32732 8520 33057 8548
rect 32732 8508 32738 8520
rect 33045 8517 33057 8520
rect 33091 8517 33103 8551
rect 33045 8511 33103 8517
rect 33965 8551 34023 8557
rect 33965 8517 33977 8551
rect 34011 8548 34023 8551
rect 34238 8548 34244 8560
rect 34011 8520 34244 8548
rect 34011 8517 34023 8520
rect 33965 8511 34023 8517
rect 34238 8508 34244 8520
rect 34296 8508 34302 8560
rect 34332 8548 34360 8588
rect 34974 8576 34980 8628
rect 35032 8616 35038 8628
rect 35621 8619 35679 8625
rect 35621 8616 35633 8619
rect 35032 8588 35633 8616
rect 35032 8576 35038 8588
rect 35621 8585 35633 8588
rect 35667 8585 35679 8619
rect 35621 8579 35679 8585
rect 34332 8520 34454 8548
rect 30958 8452 31340 8480
rect 31772 8452 32352 8480
rect 28905 8443 28963 8449
rect 19852 8384 20668 8412
rect 19852 8372 19858 8384
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 22189 8415 22247 8421
rect 22189 8412 22201 8415
rect 22152 8384 22201 8412
rect 22152 8372 22158 8384
rect 22189 8381 22201 8384
rect 22235 8381 22247 8415
rect 22189 8375 22247 8381
rect 23566 8372 23572 8424
rect 23624 8412 23630 8424
rect 23661 8415 23719 8421
rect 23661 8412 23673 8415
rect 23624 8384 23673 8412
rect 23624 8372 23630 8384
rect 23661 8381 23673 8384
rect 23707 8381 23719 8415
rect 23661 8375 23719 8381
rect 24026 8372 24032 8424
rect 24084 8412 24090 8424
rect 24397 8415 24455 8421
rect 24397 8412 24409 8415
rect 24084 8384 24409 8412
rect 24084 8372 24090 8384
rect 24397 8381 24409 8384
rect 24443 8381 24455 8415
rect 24397 8375 24455 8381
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 28350 8412 28356 8424
rect 27580 8384 28356 8412
rect 27580 8372 27586 8384
rect 28350 8372 28356 8384
rect 28408 8372 28414 8424
rect 29181 8415 29239 8421
rect 29181 8381 29193 8415
rect 29227 8381 29239 8415
rect 29181 8375 29239 8381
rect 18322 8304 18328 8356
rect 18380 8344 18386 8356
rect 20806 8344 20812 8356
rect 18380 8316 20812 8344
rect 18380 8304 18386 8316
rect 20806 8304 20812 8316
rect 20864 8304 20870 8356
rect 26234 8304 26240 8356
rect 26292 8344 26298 8356
rect 27706 8344 27712 8356
rect 26292 8316 27712 8344
rect 26292 8304 26298 8316
rect 27706 8304 27712 8316
rect 27764 8304 27770 8356
rect 14274 8276 14280 8288
rect 13924 8248 14280 8276
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 27982 8236 27988 8288
rect 28040 8276 28046 8288
rect 28537 8279 28595 8285
rect 28537 8276 28549 8279
rect 28040 8248 28549 8276
rect 28040 8236 28046 8248
rect 28537 8245 28549 8248
rect 28583 8245 28595 8279
rect 29196 8276 29224 8375
rect 29454 8372 29460 8424
rect 29512 8412 29518 8424
rect 29549 8415 29607 8421
rect 29549 8412 29561 8415
rect 29512 8384 29561 8412
rect 29512 8372 29518 8384
rect 29549 8381 29561 8384
rect 29595 8381 29607 8415
rect 29549 8375 29607 8381
rect 30190 8372 30196 8424
rect 30248 8412 30254 8424
rect 30834 8412 30840 8424
rect 30248 8384 30840 8412
rect 30248 8372 30254 8384
rect 30834 8372 30840 8384
rect 30892 8372 30898 8424
rect 31312 8412 31340 8452
rect 31312 8384 31524 8412
rect 31294 8304 31300 8356
rect 31352 8304 31358 8356
rect 31386 8304 31392 8356
rect 31444 8304 31450 8356
rect 31496 8344 31524 8384
rect 32122 8372 32128 8424
rect 32180 8412 32186 8424
rect 32217 8415 32275 8421
rect 32217 8412 32229 8415
rect 32180 8384 32229 8412
rect 32180 8372 32186 8384
rect 32217 8381 32229 8384
rect 32263 8381 32275 8415
rect 32324 8412 32352 8452
rect 32490 8440 32496 8492
rect 32548 8480 32554 8492
rect 33137 8483 33195 8489
rect 33137 8480 33149 8483
rect 32548 8452 33149 8480
rect 32548 8440 32554 8452
rect 33137 8449 33149 8452
rect 33183 8449 33195 8483
rect 33137 8443 33195 8449
rect 33321 8483 33379 8489
rect 33321 8449 33333 8483
rect 33367 8449 33379 8483
rect 33321 8443 33379 8449
rect 33336 8412 33364 8443
rect 33410 8440 33416 8492
rect 33468 8440 33474 8492
rect 33502 8440 33508 8492
rect 33560 8480 33566 8492
rect 33689 8483 33747 8489
rect 33689 8480 33701 8483
rect 33560 8452 33701 8480
rect 33560 8440 33566 8452
rect 33689 8449 33701 8452
rect 33735 8449 33747 8483
rect 35529 8483 35587 8489
rect 35529 8480 35541 8483
rect 33689 8443 33747 8449
rect 35452 8452 35541 8480
rect 35452 8421 35480 8452
rect 35529 8449 35541 8452
rect 35575 8449 35587 8483
rect 35529 8443 35587 8449
rect 32324 8384 33364 8412
rect 35437 8415 35495 8421
rect 32217 8375 32275 8381
rect 35437 8381 35449 8415
rect 35483 8381 35495 8415
rect 35437 8375 35495 8381
rect 31496 8316 32996 8344
rect 29914 8276 29920 8288
rect 29196 8248 29920 8276
rect 28537 8239 28595 8245
rect 29914 8236 29920 8248
rect 29972 8236 29978 8288
rect 31312 8276 31340 8304
rect 31573 8279 31631 8285
rect 31573 8276 31585 8279
rect 31312 8248 31585 8276
rect 31573 8245 31585 8248
rect 31619 8276 31631 8279
rect 32490 8276 32496 8288
rect 31619 8248 32496 8276
rect 31619 8245 31631 8248
rect 31573 8239 31631 8245
rect 32490 8236 32496 8248
rect 32548 8236 32554 8288
rect 32968 8276 32996 8316
rect 33042 8304 33048 8356
rect 33100 8344 33106 8356
rect 33137 8347 33195 8353
rect 33137 8344 33149 8347
rect 33100 8316 33149 8344
rect 33100 8304 33106 8316
rect 33137 8313 33149 8316
rect 33183 8313 33195 8347
rect 33137 8307 33195 8313
rect 33686 8276 33692 8288
rect 32968 8248 33692 8276
rect 33686 8236 33692 8248
rect 33744 8236 33750 8288
rect 1104 8186 37076 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 37076 8186
rect 1104 8112 37076 8134
rect 17313 8075 17371 8081
rect 17313 8041 17325 8075
rect 17359 8072 17371 8075
rect 18322 8072 18328 8084
rect 17359 8044 18328 8072
rect 17359 8041 17371 8044
rect 17313 8035 17371 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 25958 8032 25964 8084
rect 26016 8072 26022 8084
rect 26145 8075 26203 8081
rect 26145 8072 26157 8075
rect 26016 8044 26157 8072
rect 26016 8032 26022 8044
rect 26145 8041 26157 8044
rect 26191 8041 26203 8075
rect 26145 8035 26203 8041
rect 34606 8032 34612 8084
rect 34664 8072 34670 8084
rect 34977 8075 35035 8081
rect 34977 8072 34989 8075
rect 34664 8044 34989 8072
rect 34664 8032 34670 8044
rect 34977 8041 34989 8044
rect 35023 8041 35035 8075
rect 34977 8035 35035 8041
rect 23385 8007 23443 8013
rect 23385 7973 23397 8007
rect 23431 7973 23443 8007
rect 23385 7967 23443 7973
rect 14274 7896 14280 7948
rect 14332 7896 14338 7948
rect 18782 7896 18788 7948
rect 18840 7896 18846 7948
rect 21450 7896 21456 7948
rect 21508 7936 21514 7948
rect 21545 7939 21603 7945
rect 21545 7936 21557 7939
rect 21508 7908 21557 7936
rect 21508 7896 21514 7908
rect 21545 7905 21557 7908
rect 21591 7905 21603 7939
rect 21545 7899 21603 7905
rect 21821 7939 21879 7945
rect 21821 7905 21833 7939
rect 21867 7936 21879 7939
rect 23400 7936 23428 7967
rect 21867 7908 23428 7936
rect 21867 7905 21879 7908
rect 21821 7899 21879 7905
rect 23658 7896 23664 7948
rect 23716 7936 23722 7948
rect 23845 7939 23903 7945
rect 23845 7936 23857 7939
rect 23716 7908 23857 7936
rect 23716 7896 23722 7908
rect 23845 7905 23857 7908
rect 23891 7905 23903 7939
rect 23845 7899 23903 7905
rect 23934 7896 23940 7948
rect 23992 7936 23998 7948
rect 24118 7936 24124 7948
rect 23992 7908 24124 7936
rect 23992 7896 23998 7908
rect 24118 7896 24124 7908
rect 24176 7896 24182 7948
rect 25130 7896 25136 7948
rect 25188 7936 25194 7948
rect 25682 7936 25688 7948
rect 25188 7908 25688 7936
rect 25188 7896 25194 7908
rect 25682 7896 25688 7908
rect 25740 7936 25746 7948
rect 27522 7936 27528 7948
rect 25740 7908 27528 7936
rect 25740 7896 25746 7908
rect 27522 7896 27528 7908
rect 27580 7896 27586 7948
rect 27614 7896 27620 7948
rect 27672 7936 27678 7948
rect 28261 7939 28319 7945
rect 28261 7936 28273 7939
rect 27672 7908 28273 7936
rect 27672 7896 27678 7908
rect 28261 7905 28273 7908
rect 28307 7905 28319 7939
rect 28261 7899 28319 7905
rect 30190 7896 30196 7948
rect 30248 7896 30254 7948
rect 30650 7896 30656 7948
rect 30708 7896 30714 7948
rect 35986 7936 35992 7948
rect 35360 7908 35992 7936
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 15712 7840 16252 7868
rect 15712 7828 15718 7840
rect 14550 7760 14556 7812
rect 14608 7760 14614 7812
rect 16224 7800 16252 7840
rect 17218 7828 17224 7880
rect 17276 7828 17282 7880
rect 19058 7828 19064 7880
rect 19116 7828 19122 7880
rect 23290 7868 23296 7880
rect 22954 7840 23296 7868
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 23382 7828 23388 7880
rect 23440 7868 23446 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 23440 7840 24409 7868
rect 23440 7828 23446 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 29914 7828 29920 7880
rect 29972 7828 29978 7880
rect 31757 7871 31815 7877
rect 31757 7837 31769 7871
rect 31803 7868 31815 7871
rect 31846 7868 31852 7880
rect 31803 7840 31852 7868
rect 31803 7837 31815 7840
rect 31757 7831 31815 7837
rect 31846 7828 31852 7840
rect 31904 7868 31910 7880
rect 32861 7871 32919 7877
rect 32861 7868 32873 7871
rect 31904 7840 32873 7868
rect 31904 7828 31910 7840
rect 32861 7837 32873 7840
rect 32907 7868 32919 7871
rect 34054 7868 34060 7880
rect 32907 7840 34060 7868
rect 32907 7837 32919 7840
rect 32861 7831 32919 7837
rect 34054 7828 34060 7840
rect 34112 7868 34118 7880
rect 35360 7877 35388 7908
rect 35986 7896 35992 7908
rect 36044 7896 36050 7948
rect 34701 7871 34759 7877
rect 34701 7868 34713 7871
rect 34112 7840 34713 7868
rect 34112 7828 34118 7840
rect 34701 7837 34713 7840
rect 34747 7837 34759 7871
rect 35345 7871 35403 7877
rect 35345 7868 35357 7871
rect 34701 7831 34759 7837
rect 34900 7840 35357 7868
rect 17402 7800 17408 7812
rect 16224 7772 17408 7800
rect 17402 7760 17408 7772
rect 17460 7800 17466 7812
rect 17460 7772 17618 7800
rect 17460 7760 17466 7772
rect 20622 7760 20628 7812
rect 20680 7760 20686 7812
rect 21177 7803 21235 7809
rect 21177 7769 21189 7803
rect 21223 7800 21235 7803
rect 23750 7800 23756 7812
rect 21223 7772 22094 7800
rect 21223 7769 21235 7772
rect 21177 7763 21235 7769
rect 16022 7692 16028 7744
rect 16080 7692 16086 7744
rect 19705 7735 19763 7741
rect 19705 7701 19717 7735
rect 19751 7732 19763 7735
rect 20530 7732 20536 7744
rect 19751 7704 20536 7732
rect 19751 7701 19763 7704
rect 19705 7695 19763 7701
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 22066 7732 22094 7772
rect 23308 7772 23756 7800
rect 22186 7732 22192 7744
rect 22066 7704 22192 7732
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 23308 7741 23336 7772
rect 23750 7760 23756 7772
rect 23808 7760 23814 7812
rect 24673 7803 24731 7809
rect 24673 7769 24685 7803
rect 24719 7800 24731 7803
rect 24946 7800 24952 7812
rect 24719 7772 24952 7800
rect 24719 7769 24731 7772
rect 24673 7763 24731 7769
rect 24946 7760 24952 7772
rect 25004 7760 25010 7812
rect 25130 7760 25136 7812
rect 25188 7760 25194 7812
rect 27522 7760 27528 7812
rect 27580 7760 27586 7812
rect 27982 7760 27988 7812
rect 28040 7760 28046 7812
rect 30558 7760 30564 7812
rect 30616 7800 30622 7812
rect 32033 7803 32091 7809
rect 32033 7800 32045 7803
rect 30616 7772 32045 7800
rect 30616 7760 30622 7772
rect 32033 7769 32045 7772
rect 32079 7769 32091 7803
rect 32033 7763 32091 7769
rect 32950 7760 32956 7812
rect 33008 7760 33014 7812
rect 33318 7760 33324 7812
rect 33376 7800 33382 7812
rect 34900 7800 34928 7840
rect 35345 7837 35357 7840
rect 35391 7837 35403 7871
rect 35345 7831 35403 7837
rect 35434 7828 35440 7880
rect 35492 7868 35498 7880
rect 35805 7871 35863 7877
rect 35805 7868 35817 7871
rect 35492 7840 35817 7868
rect 35492 7828 35498 7840
rect 35805 7837 35817 7840
rect 35851 7837 35863 7871
rect 35805 7831 35863 7837
rect 33376 7772 34928 7800
rect 33376 7760 33382 7772
rect 36170 7760 36176 7812
rect 36228 7760 36234 7812
rect 23293 7735 23351 7741
rect 23293 7701 23305 7735
rect 23339 7701 23351 7735
rect 23293 7695 23351 7701
rect 26513 7735 26571 7741
rect 26513 7701 26525 7735
rect 26559 7732 26571 7735
rect 27890 7732 27896 7744
rect 26559 7704 27896 7732
rect 26559 7701 26571 7704
rect 26513 7695 26571 7701
rect 27890 7692 27896 7704
rect 27948 7692 27954 7744
rect 28442 7692 28448 7744
rect 28500 7732 28506 7744
rect 29549 7735 29607 7741
rect 29549 7732 29561 7735
rect 28500 7704 29561 7732
rect 28500 7692 28506 7704
rect 29549 7701 29561 7704
rect 29595 7701 29607 7735
rect 29549 7695 29607 7701
rect 30009 7735 30067 7741
rect 30009 7701 30021 7735
rect 30055 7732 30067 7735
rect 30190 7732 30196 7744
rect 30055 7704 30196 7732
rect 30055 7701 30067 7704
rect 30009 7695 30067 7701
rect 30190 7692 30196 7704
rect 30248 7692 30254 7744
rect 34241 7735 34299 7741
rect 34241 7701 34253 7735
rect 34287 7732 34299 7735
rect 34330 7732 34336 7744
rect 34287 7704 34336 7732
rect 34287 7701 34299 7704
rect 34241 7695 34299 7701
rect 34330 7692 34336 7704
rect 34388 7692 34394 7744
rect 1104 7642 37076 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 37076 7642
rect 1104 7568 37076 7590
rect 18966 7528 18972 7540
rect 15488 7500 18972 7528
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 15013 7463 15071 7469
rect 15013 7460 15025 7463
rect 14608 7432 15025 7460
rect 14608 7420 14614 7432
rect 15013 7429 15025 7432
rect 15059 7429 15071 7463
rect 15013 7423 15071 7429
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 15488 7401 15516 7500
rect 18966 7488 18972 7500
rect 19024 7488 19030 7540
rect 22465 7531 22523 7537
rect 22465 7497 22477 7531
rect 22511 7528 22523 7531
rect 23566 7528 23572 7540
rect 22511 7500 23572 7528
rect 22511 7497 22523 7500
rect 22465 7491 22523 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 25590 7488 25596 7540
rect 25648 7528 25654 7540
rect 26053 7531 26111 7537
rect 26053 7528 26065 7531
rect 25648 7500 26065 7528
rect 25648 7488 25654 7500
rect 26053 7497 26065 7500
rect 26099 7497 26111 7531
rect 26053 7491 26111 7497
rect 27433 7531 27491 7537
rect 27433 7497 27445 7531
rect 27479 7528 27491 7531
rect 27890 7528 27896 7540
rect 27479 7500 27896 7528
rect 27479 7497 27491 7500
rect 27433 7491 27491 7497
rect 27890 7488 27896 7500
rect 27948 7488 27954 7540
rect 29917 7531 29975 7537
rect 29917 7497 29929 7531
rect 29963 7528 29975 7531
rect 30098 7528 30104 7540
rect 29963 7500 30104 7528
rect 29963 7497 29975 7500
rect 29917 7491 29975 7497
rect 30098 7488 30104 7500
rect 30156 7488 30162 7540
rect 17402 7420 17408 7472
rect 17460 7420 17466 7472
rect 20622 7460 20628 7472
rect 20470 7432 20628 7460
rect 20622 7420 20628 7432
rect 20680 7420 20686 7472
rect 23290 7420 23296 7472
rect 23348 7420 23354 7472
rect 23937 7463 23995 7469
rect 23937 7429 23949 7463
rect 23983 7460 23995 7463
rect 24026 7460 24032 7472
rect 23983 7432 24032 7460
rect 23983 7429 23995 7432
rect 23937 7423 23995 7429
rect 24026 7420 24032 7432
rect 24084 7420 24090 7472
rect 24578 7420 24584 7472
rect 24636 7420 24642 7472
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 27341 7463 27399 7469
rect 27341 7429 27353 7463
rect 27387 7460 27399 7463
rect 27798 7460 27804 7472
rect 27387 7432 27804 7460
rect 27387 7429 27399 7432
rect 27341 7423 27399 7429
rect 27798 7420 27804 7432
rect 27856 7420 27862 7472
rect 28442 7420 28448 7472
rect 28500 7420 28506 7472
rect 29730 7460 29736 7472
rect 29670 7432 29736 7460
rect 29730 7420 29736 7432
rect 29788 7420 29794 7472
rect 31018 7420 31024 7472
rect 31076 7460 31082 7472
rect 31665 7463 31723 7469
rect 31665 7460 31677 7463
rect 31076 7432 31677 7460
rect 31076 7420 31082 7432
rect 31665 7429 31677 7432
rect 31711 7429 31723 7463
rect 31665 7423 31723 7429
rect 31846 7420 31852 7472
rect 31904 7420 31910 7472
rect 33686 7460 33692 7472
rect 33626 7432 33692 7460
rect 33686 7420 33692 7432
rect 33744 7420 33750 7472
rect 34054 7420 34060 7472
rect 34112 7460 34118 7472
rect 34149 7463 34207 7469
rect 34149 7460 34161 7463
rect 34112 7432 34161 7460
rect 34112 7420 34118 7432
rect 34149 7429 34161 7432
rect 34195 7429 34207 7463
rect 34149 7423 34207 7429
rect 34885 7463 34943 7469
rect 34885 7429 34897 7463
rect 34931 7460 34943 7463
rect 35253 7463 35311 7469
rect 35253 7460 35265 7463
rect 34931 7432 35265 7460
rect 34931 7429 34943 7432
rect 34885 7423 34943 7429
rect 35253 7429 35265 7432
rect 35299 7460 35311 7463
rect 35434 7460 35440 7472
rect 35299 7432 35440 7460
rect 35299 7429 35311 7432
rect 35253 7423 35311 7429
rect 35434 7420 35440 7432
rect 35492 7420 35498 7472
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15252 7364 15485 7392
rect 15252 7352 15258 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 15620 7364 15669 7392
rect 15620 7352 15626 7364
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16022 7392 16028 7404
rect 15795 7364 16028 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7392 21235 7395
rect 21450 7392 21456 7404
rect 21223 7364 21456 7392
rect 21223 7361 21235 7364
rect 21177 7355 21235 7361
rect 21450 7352 21456 7364
rect 21508 7392 21514 7404
rect 21508 7364 22094 7392
rect 21508 7352 21514 7364
rect 22066 7336 22094 7364
rect 27614 7352 27620 7404
rect 27672 7392 27678 7404
rect 28166 7392 28172 7404
rect 27672 7364 28172 7392
rect 27672 7352 27678 7364
rect 28166 7352 28172 7364
rect 28224 7352 28230 7404
rect 30282 7352 30288 7404
rect 30340 7352 30346 7404
rect 30558 7352 30564 7404
rect 30616 7392 30622 7404
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 30616 7364 31217 7392
rect 30616 7352 30622 7364
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 32122 7352 32128 7404
rect 32180 7352 32186 7404
rect 34330 7352 34336 7404
rect 34388 7352 34394 7404
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7324 17003 7327
rect 18506 7324 18512 7336
rect 16991 7296 18512 7324
rect 16991 7293 17003 7296
rect 16945 7287 17003 7293
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 20898 7284 20904 7336
rect 20956 7284 20962 7336
rect 22066 7296 22100 7336
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 24213 7327 24271 7333
rect 24213 7293 24225 7327
rect 24259 7324 24271 7327
rect 24305 7327 24363 7333
rect 24305 7324 24317 7327
rect 24259 7296 24317 7324
rect 24259 7293 24271 7296
rect 24213 7287 24271 7293
rect 24305 7293 24317 7296
rect 24351 7293 24363 7327
rect 24305 7287 24363 7293
rect 18417 7191 18475 7197
rect 18417 7157 18429 7191
rect 18463 7188 18475 7191
rect 18598 7188 18604 7200
rect 18463 7160 18604 7188
rect 18463 7157 18475 7160
rect 18417 7151 18475 7157
rect 18598 7148 18604 7160
rect 18656 7188 18662 7200
rect 19242 7188 19248 7200
rect 18656 7160 19248 7188
rect 18656 7148 18662 7160
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 19429 7191 19487 7197
rect 19429 7157 19441 7191
rect 19475 7188 19487 7191
rect 20438 7188 20444 7200
rect 19475 7160 20444 7188
rect 19475 7157 19487 7160
rect 19429 7151 19487 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 23382 7148 23388 7200
rect 23440 7188 23446 7200
rect 24228 7188 24256 7287
rect 27522 7284 27528 7336
rect 27580 7284 27586 7336
rect 30006 7284 30012 7336
rect 30064 7284 30070 7336
rect 31754 7284 31760 7336
rect 31812 7324 31818 7336
rect 32401 7327 32459 7333
rect 32401 7324 32413 7327
rect 31812 7296 32413 7324
rect 31812 7284 31818 7296
rect 32401 7293 32413 7296
rect 32447 7293 32459 7327
rect 32401 7287 32459 7293
rect 31389 7259 31447 7265
rect 31389 7225 31401 7259
rect 31435 7256 31447 7259
rect 31435 7228 32260 7256
rect 31435 7225 31447 7228
rect 31389 7219 31447 7225
rect 23440 7160 24256 7188
rect 23440 7148 23446 7160
rect 26970 7148 26976 7200
rect 27028 7148 27034 7200
rect 32232 7188 32260 7228
rect 34514 7216 34520 7268
rect 34572 7256 34578 7268
rect 35069 7259 35127 7265
rect 35069 7256 35081 7259
rect 34572 7228 35081 7256
rect 34572 7216 34578 7228
rect 35069 7225 35081 7228
rect 35115 7225 35127 7259
rect 35069 7219 35127 7225
rect 32490 7188 32496 7200
rect 32232 7160 32496 7188
rect 32490 7148 32496 7160
rect 32548 7148 32554 7200
rect 1104 7098 37076 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 37076 7098
rect 1104 7024 37076 7046
rect 22186 6944 22192 6996
rect 22244 6944 22250 6996
rect 26316 6987 26374 6993
rect 26316 6953 26328 6987
rect 26362 6984 26374 6987
rect 26970 6984 26976 6996
rect 26362 6956 26976 6984
rect 26362 6953 26374 6956
rect 26316 6947 26374 6953
rect 26970 6944 26976 6956
rect 27028 6944 27034 6996
rect 27798 6944 27804 6996
rect 27856 6944 27862 6996
rect 31113 6987 31171 6993
rect 31113 6984 31125 6987
rect 30300 6956 31125 6984
rect 30300 6928 30328 6956
rect 31113 6953 31125 6956
rect 31159 6953 31171 6987
rect 31113 6947 31171 6953
rect 34057 6987 34115 6993
rect 34057 6953 34069 6987
rect 34103 6984 34115 6987
rect 34333 6987 34391 6993
rect 34333 6984 34345 6987
rect 34103 6956 34345 6984
rect 34103 6953 34115 6956
rect 34057 6947 34115 6953
rect 34333 6953 34345 6956
rect 34379 6953 34391 6987
rect 34333 6947 34391 6953
rect 30282 6876 30288 6928
rect 30340 6876 30346 6928
rect 30377 6919 30435 6925
rect 30377 6885 30389 6919
rect 30423 6916 30435 6919
rect 30423 6888 30604 6916
rect 30423 6885 30435 6888
rect 30377 6879 30435 6885
rect 16022 6848 16028 6860
rect 15580 6820 16028 6848
rect 15580 6789 15608 6820
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 19058 6848 19064 6860
rect 16724 6820 19064 6848
rect 16724 6808 16730 6820
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 20438 6808 20444 6860
rect 20496 6848 20502 6860
rect 20496 6820 22094 6848
rect 20496 6808 20502 6820
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6780 15439 6783
rect 15565 6783 15623 6789
rect 15427 6752 15516 6780
rect 15427 6749 15439 6752
rect 15381 6743 15439 6749
rect 14826 6672 14832 6724
rect 14884 6712 14890 6724
rect 14921 6715 14979 6721
rect 14921 6712 14933 6715
rect 14884 6684 14933 6712
rect 14884 6672 14890 6684
rect 14921 6681 14933 6684
rect 14967 6681 14979 6715
rect 14921 6675 14979 6681
rect 15488 6644 15516 6752
rect 15565 6749 15577 6783
rect 15611 6749 15623 6783
rect 15565 6743 15623 6749
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6780 15715 6783
rect 15746 6780 15752 6792
rect 15703 6752 15752 6780
rect 15703 6749 15715 6752
rect 15657 6743 15715 6749
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 19024 6752 19257 6780
rect 19024 6740 19030 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6780 21051 6783
rect 21266 6780 21272 6792
rect 21039 6752 21272 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 21542 6740 21548 6792
rect 21600 6740 21606 6792
rect 21726 6740 21732 6792
rect 21784 6740 21790 6792
rect 21818 6740 21824 6792
rect 21876 6740 21882 6792
rect 22066 6780 22094 6820
rect 22462 6808 22468 6860
rect 22520 6848 22526 6860
rect 22833 6851 22891 6857
rect 22833 6848 22845 6851
rect 22520 6820 22845 6848
rect 22520 6808 22526 6820
rect 22833 6817 22845 6820
rect 22879 6848 22891 6851
rect 24118 6848 24124 6860
rect 22879 6820 24124 6848
rect 22879 6817 22891 6820
rect 22833 6811 22891 6817
rect 24118 6808 24124 6820
rect 24176 6808 24182 6860
rect 24946 6808 24952 6860
rect 25004 6808 25010 6860
rect 25685 6851 25743 6857
rect 25685 6817 25697 6851
rect 25731 6848 25743 6851
rect 25958 6848 25964 6860
rect 25731 6820 25964 6848
rect 25731 6817 25743 6820
rect 25685 6811 25743 6817
rect 25958 6808 25964 6820
rect 26016 6808 26022 6860
rect 28166 6848 28172 6860
rect 26068 6820 28172 6848
rect 26068 6792 26096 6820
rect 28166 6808 28172 6820
rect 28224 6808 28230 6860
rect 30006 6808 30012 6860
rect 30064 6848 30070 6860
rect 30469 6851 30527 6857
rect 30469 6848 30481 6851
rect 30064 6820 30481 6848
rect 30064 6808 30070 6820
rect 30469 6817 30481 6820
rect 30515 6817 30527 6851
rect 30469 6811 30527 6817
rect 22649 6783 22707 6789
rect 22649 6780 22661 6783
rect 22066 6752 22661 6780
rect 22649 6749 22661 6752
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 22922 6740 22928 6792
rect 22980 6780 22986 6792
rect 25314 6780 25320 6792
rect 22980 6752 25320 6780
rect 22980 6740 22986 6752
rect 25314 6740 25320 6752
rect 25372 6780 25378 6792
rect 25409 6783 25467 6789
rect 25409 6780 25421 6783
rect 25372 6752 25421 6780
rect 25372 6740 25378 6752
rect 25409 6749 25421 6752
rect 25455 6749 25467 6783
rect 25409 6743 25467 6749
rect 25590 6740 25596 6792
rect 25648 6740 25654 6792
rect 26050 6740 26056 6792
rect 26108 6740 26114 6792
rect 27338 6740 27344 6792
rect 27396 6780 27402 6792
rect 30576 6780 30604 6888
rect 30650 6808 30656 6860
rect 30708 6848 30714 6860
rect 31128 6848 31156 6947
rect 34146 6876 34152 6928
rect 34204 6876 34210 6928
rect 31481 6851 31539 6857
rect 30708 6820 31064 6848
rect 31128 6820 31432 6848
rect 30708 6808 30714 6820
rect 30929 6783 30987 6789
rect 30929 6780 30941 6783
rect 27396 6766 27462 6780
rect 27396 6752 27476 6766
rect 30576 6752 30941 6780
rect 27396 6740 27402 6752
rect 16942 6672 16948 6724
rect 17000 6672 17006 6724
rect 17402 6672 17408 6724
rect 17460 6672 17466 6724
rect 19518 6672 19524 6724
rect 19576 6712 19582 6724
rect 21085 6715 21143 6721
rect 21085 6712 21097 6715
rect 19576 6684 21097 6712
rect 19576 6672 19582 6684
rect 21085 6681 21097 6684
rect 21131 6681 21143 6715
rect 21085 6675 21143 6681
rect 17862 6644 17868 6656
rect 15488 6616 17868 6644
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 18414 6604 18420 6656
rect 18472 6604 18478 6656
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 22557 6647 22615 6653
rect 22557 6644 22569 6647
rect 20588 6616 22569 6644
rect 20588 6604 20594 6616
rect 22557 6613 22569 6616
rect 22603 6613 22615 6647
rect 27448 6644 27476 6752
rect 30009 6715 30067 6721
rect 30009 6681 30021 6715
rect 30055 6712 30067 6715
rect 30374 6712 30380 6724
rect 30055 6684 30380 6712
rect 30055 6681 30067 6684
rect 30009 6675 30067 6681
rect 30374 6672 30380 6684
rect 30432 6712 30438 6724
rect 30558 6712 30564 6724
rect 30432 6684 30564 6712
rect 30432 6672 30438 6684
rect 30558 6672 30564 6684
rect 30616 6672 30622 6724
rect 29730 6644 29736 6656
rect 27448 6616 29736 6644
rect 22557 6607 22615 6613
rect 29730 6604 29736 6616
rect 29788 6604 29794 6656
rect 30760 6644 30788 6752
rect 30929 6749 30941 6752
rect 30975 6749 30987 6783
rect 31036 6780 31064 6820
rect 31404 6789 31432 6820
rect 31481 6817 31493 6851
rect 31527 6848 31539 6851
rect 31754 6848 31760 6860
rect 31527 6820 31760 6848
rect 31527 6817 31539 6820
rect 31481 6811 31539 6817
rect 31754 6808 31760 6820
rect 31812 6808 31818 6860
rect 32122 6808 32128 6860
rect 32180 6848 32186 6860
rect 32309 6851 32367 6857
rect 32309 6848 32321 6851
rect 32180 6820 32321 6848
rect 32180 6808 32186 6820
rect 32309 6817 32321 6820
rect 32355 6848 32367 6851
rect 33042 6848 33048 6860
rect 32355 6820 33048 6848
rect 32355 6817 32367 6820
rect 32309 6811 32367 6817
rect 33042 6808 33048 6820
rect 33100 6808 33106 6860
rect 34348 6848 34376 6947
rect 34348 6820 34744 6848
rect 31113 6783 31171 6789
rect 31113 6780 31125 6783
rect 31036 6752 31125 6780
rect 30929 6743 30987 6749
rect 31113 6749 31125 6752
rect 31159 6749 31171 6783
rect 31113 6743 31171 6749
rect 31389 6783 31447 6789
rect 31389 6749 31401 6783
rect 31435 6749 31447 6783
rect 31389 6743 31447 6749
rect 31573 6783 31631 6789
rect 31573 6749 31585 6783
rect 31619 6780 31631 6783
rect 32214 6780 32220 6792
rect 31619 6752 32220 6780
rect 31619 6749 31631 6752
rect 31573 6743 31631 6749
rect 32214 6740 32220 6752
rect 32272 6740 32278 6792
rect 33686 6740 33692 6792
rect 33744 6780 33750 6792
rect 34330 6780 34336 6792
rect 33744 6752 34336 6780
rect 33744 6740 33750 6752
rect 34330 6740 34336 6752
rect 34388 6740 34394 6792
rect 34716 6789 34744 6820
rect 34900 6820 35388 6848
rect 34701 6783 34759 6789
rect 34701 6749 34713 6783
rect 34747 6749 34759 6783
rect 34701 6743 34759 6749
rect 32582 6672 32588 6724
rect 32640 6672 32646 6724
rect 34054 6672 34060 6724
rect 34112 6712 34118 6724
rect 34517 6715 34575 6721
rect 34517 6712 34529 6715
rect 34112 6684 34529 6712
rect 34112 6672 34118 6684
rect 34517 6681 34529 6684
rect 34563 6712 34575 6715
rect 34900 6712 34928 6820
rect 35360 6789 35388 6820
rect 34977 6783 35035 6789
rect 34977 6749 34989 6783
rect 35023 6780 35035 6783
rect 35345 6783 35403 6789
rect 35023 6752 35204 6780
rect 35023 6749 35035 6752
rect 34977 6743 35035 6749
rect 34563 6684 34928 6712
rect 34563 6681 34575 6684
rect 34517 6675 34575 6681
rect 33318 6644 33324 6656
rect 30760 6616 33324 6644
rect 33318 6604 33324 6616
rect 33376 6604 33382 6656
rect 34317 6647 34375 6653
rect 34317 6613 34329 6647
rect 34363 6644 34375 6647
rect 34606 6644 34612 6656
rect 34363 6616 34612 6644
rect 34363 6613 34375 6616
rect 34317 6607 34375 6613
rect 34606 6604 34612 6616
rect 34664 6604 34670 6656
rect 34790 6604 34796 6656
rect 34848 6604 34854 6656
rect 35176 6653 35204 6752
rect 35345 6749 35357 6783
rect 35391 6749 35403 6783
rect 35345 6743 35403 6749
rect 35161 6647 35219 6653
rect 35161 6613 35173 6647
rect 35207 6613 35219 6647
rect 35161 6607 35219 6613
rect 1104 6554 37076 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 37076 6554
rect 1104 6480 37076 6502
rect 14274 6400 14280 6452
rect 14332 6400 14338 6452
rect 18966 6440 18972 6452
rect 18340 6412 18972 6440
rect 14090 6372 14096 6384
rect 13832 6344 14096 6372
rect 13832 6313 13860 6344
rect 14090 6332 14096 6344
rect 14148 6372 14154 6384
rect 14292 6372 14320 6400
rect 15654 6372 15660 6384
rect 14148 6344 14320 6372
rect 15318 6344 15660 6372
rect 14148 6332 14154 6344
rect 15654 6332 15660 6344
rect 15712 6332 15718 6384
rect 16942 6332 16948 6384
rect 17000 6372 17006 6384
rect 17313 6375 17371 6381
rect 17313 6372 17325 6375
rect 17000 6344 17325 6372
rect 17000 6332 17006 6344
rect 17313 6341 17325 6344
rect 17359 6341 17371 6375
rect 18138 6372 18144 6384
rect 17313 6335 17371 6341
rect 17788 6344 18144 6372
rect 17788 6313 17816 6344
rect 18138 6332 18144 6344
rect 18196 6372 18202 6384
rect 18340 6372 18368 6412
rect 18966 6400 18972 6412
rect 19024 6440 19030 6452
rect 21542 6440 21548 6452
rect 19024 6412 21548 6440
rect 19024 6400 19030 6412
rect 21542 6400 21548 6412
rect 21600 6400 21606 6452
rect 25682 6440 25688 6452
rect 24780 6412 25688 6440
rect 18196 6344 18368 6372
rect 18432 6344 19196 6372
rect 18196 6332 18202 6344
rect 18432 6316 18460 6344
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 17773 6307 17831 6313
rect 17773 6273 17785 6307
rect 17819 6273 17831 6307
rect 17773 6267 17831 6273
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6304 18107 6307
rect 18414 6304 18420 6316
rect 18095 6276 18420 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14826 6236 14832 6248
rect 14139 6208 14832 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 17972 6236 18000 6267
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 18506 6264 18512 6316
rect 18564 6264 18570 6316
rect 19168 6313 19196 6344
rect 20898 6332 20904 6384
rect 20956 6372 20962 6384
rect 21177 6375 21235 6381
rect 21177 6372 21189 6375
rect 20956 6344 21189 6372
rect 20956 6332 20962 6344
rect 21177 6341 21189 6344
rect 21223 6341 21235 6375
rect 22922 6372 22928 6384
rect 21177 6335 21235 6341
rect 22112 6344 22928 6372
rect 18969 6307 19027 6313
rect 18969 6304 18981 6307
rect 18892 6276 18981 6304
rect 18322 6236 18328 6248
rect 17972 6208 18328 6236
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 17862 6128 17868 6180
rect 17920 6168 17926 6180
rect 18892 6168 18920 6276
rect 18969 6273 18981 6276
rect 19015 6273 19027 6307
rect 18969 6267 19027 6273
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 19242 6264 19248 6316
rect 19300 6264 19306 6316
rect 20438 6264 20444 6316
rect 20496 6264 20502 6316
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 20717 6307 20775 6313
rect 20717 6273 20729 6307
rect 20763 6304 20775 6307
rect 22112 6304 22140 6344
rect 22922 6332 22928 6344
rect 22980 6332 22986 6384
rect 20763 6276 22140 6304
rect 20763 6273 20775 6276
rect 20717 6267 20775 6273
rect 20548 6236 20576 6267
rect 22186 6264 22192 6316
rect 22244 6264 22250 6316
rect 24670 6264 24676 6316
rect 24728 6304 24734 6316
rect 24780 6304 24808 6412
rect 25682 6400 25688 6412
rect 25740 6400 25746 6452
rect 29730 6400 29736 6452
rect 29788 6440 29794 6452
rect 33873 6443 33931 6449
rect 29788 6412 30420 6440
rect 29788 6400 29794 6412
rect 27525 6375 27583 6381
rect 27525 6341 27537 6375
rect 27571 6372 27583 6375
rect 28534 6372 28540 6384
rect 27571 6344 28540 6372
rect 27571 6341 27583 6344
rect 27525 6335 27583 6341
rect 28534 6332 28540 6344
rect 28592 6332 28598 6384
rect 29748 6372 29776 6400
rect 30392 6384 30420 6412
rect 33873 6409 33885 6443
rect 33919 6440 33931 6443
rect 33919 6412 34284 6440
rect 33919 6409 33931 6412
rect 33873 6403 33931 6409
rect 29670 6344 29776 6372
rect 30374 6332 30380 6384
rect 30432 6372 30438 6384
rect 30432 6344 30958 6372
rect 30432 6332 30438 6344
rect 32582 6332 32588 6384
rect 32640 6372 32646 6384
rect 32769 6375 32827 6381
rect 32769 6372 32781 6375
rect 32640 6344 32781 6372
rect 32640 6332 32646 6344
rect 32769 6341 32781 6344
rect 32815 6341 32827 6375
rect 32769 6335 32827 6341
rect 33505 6375 33563 6381
rect 33505 6341 33517 6375
rect 33551 6372 33563 6375
rect 33594 6372 33600 6384
rect 33551 6344 33600 6372
rect 33551 6341 33563 6344
rect 33505 6335 33563 6341
rect 33594 6332 33600 6344
rect 33652 6332 33658 6384
rect 33778 6381 33784 6384
rect 33721 6375 33784 6381
rect 33721 6341 33733 6375
rect 33767 6341 33784 6375
rect 33721 6335 33784 6341
rect 33778 6332 33784 6335
rect 33836 6332 33842 6384
rect 34146 6372 34152 6384
rect 33980 6344 34152 6372
rect 24728 6290 24808 6304
rect 24728 6276 24794 6290
rect 24728 6264 24734 6276
rect 32214 6264 32220 6316
rect 32272 6304 32278 6316
rect 33137 6307 33195 6313
rect 33137 6304 33149 6307
rect 32272 6276 33149 6304
rect 32272 6264 32278 6276
rect 21818 6236 21824 6248
rect 20548 6208 21824 6236
rect 21818 6196 21824 6208
rect 21876 6196 21882 6248
rect 22278 6196 22284 6248
rect 22336 6196 22342 6248
rect 22462 6196 22468 6248
rect 22520 6196 22526 6248
rect 23106 6196 23112 6248
rect 23164 6236 23170 6248
rect 23382 6236 23388 6248
rect 23164 6208 23388 6236
rect 23164 6196 23170 6208
rect 23382 6196 23388 6208
rect 23440 6196 23446 6248
rect 23661 6239 23719 6245
rect 23661 6205 23673 6239
rect 23707 6236 23719 6239
rect 24394 6236 24400 6248
rect 23707 6208 24400 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 24394 6196 24400 6208
rect 24452 6196 24458 6248
rect 27430 6196 27436 6248
rect 27488 6236 27494 6248
rect 27617 6239 27675 6245
rect 27617 6236 27629 6239
rect 27488 6208 27629 6236
rect 27488 6196 27494 6208
rect 27617 6205 27629 6208
rect 27663 6205 27675 6239
rect 27617 6199 27675 6205
rect 27706 6196 27712 6248
rect 27764 6236 27770 6248
rect 27801 6239 27859 6245
rect 27801 6236 27813 6239
rect 27764 6208 27813 6236
rect 27764 6196 27770 6208
rect 27801 6205 27813 6208
rect 27847 6236 27859 6239
rect 28074 6236 28080 6248
rect 27847 6208 28080 6236
rect 27847 6205 27859 6208
rect 27801 6199 27859 6205
rect 28074 6196 28080 6208
rect 28132 6196 28138 6248
rect 28166 6196 28172 6248
rect 28224 6196 28230 6248
rect 28445 6239 28503 6245
rect 28445 6205 28457 6239
rect 28491 6236 28503 6239
rect 30098 6236 30104 6248
rect 28491 6208 30104 6236
rect 28491 6205 28503 6208
rect 28445 6199 28503 6205
rect 30098 6196 30104 6208
rect 30156 6196 30162 6248
rect 30193 6239 30251 6245
rect 30193 6205 30205 6239
rect 30239 6205 30251 6239
rect 30193 6199 30251 6205
rect 17920 6140 18920 6168
rect 17920 6128 17926 6140
rect 22094 6128 22100 6180
rect 22152 6168 22158 6180
rect 23124 6168 23152 6196
rect 22152 6140 23152 6168
rect 22152 6128 22158 6140
rect 29454 6128 29460 6180
rect 29512 6168 29518 6180
rect 30208 6168 30236 6199
rect 30466 6196 30472 6248
rect 30524 6196 30530 6248
rect 31941 6239 31999 6245
rect 31941 6205 31953 6239
rect 31987 6236 31999 6239
rect 32674 6236 32680 6248
rect 31987 6208 32680 6236
rect 31987 6205 31999 6208
rect 31941 6199 31999 6205
rect 32674 6196 32680 6208
rect 32732 6196 32738 6248
rect 29512 6140 30236 6168
rect 32968 6168 32996 6276
rect 33137 6273 33149 6276
rect 33183 6273 33195 6307
rect 33137 6267 33195 6273
rect 33321 6307 33379 6313
rect 33321 6273 33333 6307
rect 33367 6304 33379 6307
rect 33980 6304 34008 6344
rect 34146 6332 34152 6344
rect 34204 6332 34210 6384
rect 34256 6381 34284 6412
rect 34241 6375 34299 6381
rect 34241 6341 34253 6375
rect 34287 6341 34299 6375
rect 34241 6335 34299 6341
rect 34330 6332 34336 6384
rect 34388 6372 34394 6384
rect 34388 6344 34730 6372
rect 34388 6332 34394 6344
rect 33367 6276 34008 6304
rect 33367 6273 33379 6276
rect 33321 6267 33379 6273
rect 33042 6196 33048 6248
rect 33100 6236 33106 6248
rect 33965 6239 34023 6245
rect 33965 6236 33977 6239
rect 33100 6208 33977 6236
rect 33100 6196 33106 6208
rect 33965 6205 33977 6208
rect 34011 6205 34023 6239
rect 34790 6236 34796 6248
rect 33965 6199 34023 6205
rect 34072 6208 34796 6236
rect 34072 6168 34100 6208
rect 34790 6196 34796 6208
rect 34848 6196 34854 6248
rect 32968 6140 34100 6168
rect 29512 6128 29518 6140
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 15436 6072 15577 6100
rect 15436 6060 15442 6072
rect 15565 6069 15577 6072
rect 15611 6100 15623 6103
rect 15746 6100 15752 6112
rect 15611 6072 15752 6100
rect 15611 6069 15623 6072
rect 15565 6063 15623 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 21821 6103 21879 6109
rect 21821 6069 21833 6103
rect 21867 6100 21879 6103
rect 23290 6100 23296 6112
rect 21867 6072 23296 6100
rect 21867 6069 21879 6072
rect 21821 6063 21879 6069
rect 23290 6060 23296 6072
rect 23348 6060 23354 6112
rect 25130 6060 25136 6112
rect 25188 6060 25194 6112
rect 27154 6060 27160 6112
rect 27212 6060 27218 6112
rect 29914 6060 29920 6112
rect 29972 6060 29978 6112
rect 30208 6100 30236 6140
rect 36722 6128 36728 6180
rect 36780 6128 36786 6180
rect 32122 6100 32128 6112
rect 30208 6072 32128 6100
rect 32122 6060 32128 6072
rect 32180 6060 32186 6112
rect 32217 6103 32275 6109
rect 32217 6069 32229 6103
rect 32263 6100 32275 6103
rect 32306 6100 32312 6112
rect 32263 6072 32312 6100
rect 32263 6069 32275 6072
rect 32217 6063 32275 6069
rect 32306 6060 32312 6072
rect 32364 6060 32370 6112
rect 33686 6060 33692 6112
rect 33744 6060 33750 6112
rect 33778 6060 33784 6112
rect 33836 6100 33842 6112
rect 35713 6103 35771 6109
rect 35713 6100 35725 6103
rect 33836 6072 35725 6100
rect 33836 6060 33842 6072
rect 35713 6069 35725 6072
rect 35759 6069 35771 6103
rect 35713 6063 35771 6069
rect 1104 6010 37076 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 37076 6010
rect 1104 5936 37076 5958
rect 20993 5899 21051 5905
rect 20993 5865 21005 5899
rect 21039 5896 21051 5899
rect 21818 5896 21824 5908
rect 21039 5868 21824 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 21818 5856 21824 5868
rect 21876 5856 21882 5908
rect 25948 5899 26006 5905
rect 25948 5865 25960 5899
rect 25994 5896 26006 5899
rect 27525 5899 27583 5905
rect 27525 5896 27537 5899
rect 25994 5868 27537 5896
rect 25994 5865 26006 5868
rect 25948 5859 26006 5865
rect 27525 5865 27537 5868
rect 27571 5865 27583 5899
rect 27525 5859 27583 5865
rect 30193 5899 30251 5905
rect 30193 5865 30205 5899
rect 30239 5896 30251 5899
rect 30466 5896 30472 5908
rect 30239 5868 30472 5896
rect 30239 5865 30251 5868
rect 30193 5859 30251 5865
rect 30466 5856 30472 5868
rect 30524 5856 30530 5908
rect 33594 5856 33600 5908
rect 33652 5856 33658 5908
rect 33686 5856 33692 5908
rect 33744 5896 33750 5908
rect 34606 5896 34612 5908
rect 33744 5868 34612 5896
rect 33744 5856 33750 5868
rect 34606 5856 34612 5868
rect 34664 5896 34670 5908
rect 35342 5896 35348 5908
rect 34664 5868 35348 5896
rect 34664 5856 34670 5868
rect 35342 5856 35348 5868
rect 35400 5856 35406 5908
rect 27430 5788 27436 5840
rect 27488 5788 27494 5840
rect 33778 5828 33784 5840
rect 33152 5800 33784 5828
rect 15105 5763 15163 5769
rect 15105 5729 15117 5763
rect 15151 5760 15163 5763
rect 15838 5760 15844 5772
rect 15151 5732 15844 5760
rect 15151 5729 15163 5732
rect 15105 5723 15163 5729
rect 15838 5720 15844 5732
rect 15896 5760 15902 5772
rect 15896 5732 16160 5760
rect 15896 5720 15902 5732
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 14829 5655 14887 5661
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5692 15071 5695
rect 15378 5692 15384 5704
rect 15059 5664 15384 5692
rect 15059 5661 15071 5664
rect 15013 5655 15071 5661
rect 14366 5584 14372 5636
rect 14424 5584 14430 5636
rect 14844 5624 14872 5655
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 16132 5701 16160 5732
rect 16574 5720 16580 5772
rect 16632 5720 16638 5772
rect 19058 5720 19064 5772
rect 19116 5760 19122 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 19116 5732 19257 5760
rect 19116 5720 19122 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19518 5720 19524 5772
rect 19576 5720 19582 5772
rect 21361 5763 21419 5769
rect 21361 5729 21373 5763
rect 21407 5760 21419 5763
rect 22278 5760 22284 5772
rect 21407 5732 22284 5760
rect 21407 5729 21419 5732
rect 21361 5723 21419 5729
rect 22278 5720 22284 5732
rect 22336 5760 22342 5772
rect 23937 5763 23995 5769
rect 23937 5760 23949 5763
rect 22336 5732 23949 5760
rect 22336 5720 22342 5732
rect 23937 5729 23949 5732
rect 23983 5729 23995 5763
rect 23937 5723 23995 5729
rect 24394 5720 24400 5772
rect 24452 5720 24458 5772
rect 25130 5720 25136 5772
rect 25188 5720 25194 5772
rect 26050 5760 26056 5772
rect 25700 5732 26056 5760
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16209 5695 16267 5701
rect 16209 5661 16221 5695
rect 16255 5661 16267 5695
rect 16209 5655 16267 5661
rect 15194 5624 15200 5636
rect 14844 5596 15200 5624
rect 15194 5584 15200 5596
rect 15252 5584 15258 5636
rect 15473 5627 15531 5633
rect 15473 5593 15485 5627
rect 15519 5624 15531 5627
rect 15562 5624 15568 5636
rect 15519 5596 15568 5624
rect 15519 5593 15531 5596
rect 15473 5587 15531 5593
rect 15562 5584 15568 5596
rect 15620 5584 15626 5636
rect 16224 5624 16252 5655
rect 23106 5652 23112 5704
rect 23164 5652 23170 5704
rect 23661 5695 23719 5701
rect 23661 5661 23673 5695
rect 23707 5661 23719 5695
rect 23661 5655 23719 5661
rect 16758 5624 16764 5636
rect 16224 5596 16764 5624
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 16850 5584 16856 5636
rect 16908 5584 16914 5636
rect 17402 5584 17408 5636
rect 17460 5584 17466 5636
rect 20530 5584 20536 5636
rect 20588 5584 20594 5636
rect 22278 5584 22284 5636
rect 22336 5584 22342 5636
rect 22833 5627 22891 5633
rect 22833 5593 22845 5627
rect 22879 5624 22891 5627
rect 23201 5627 23259 5633
rect 23201 5624 23213 5627
rect 22879 5596 23213 5624
rect 22879 5593 22891 5596
rect 22833 5587 22891 5593
rect 23201 5593 23213 5596
rect 23247 5593 23259 5627
rect 23201 5587 23259 5593
rect 18322 5516 18328 5568
rect 18380 5516 18386 5568
rect 21542 5516 21548 5568
rect 21600 5556 21606 5568
rect 23676 5556 23704 5655
rect 23842 5652 23848 5704
rect 23900 5652 23906 5704
rect 24854 5652 24860 5704
rect 24912 5652 24918 5704
rect 24946 5652 24952 5704
rect 25004 5692 25010 5704
rect 25041 5695 25099 5701
rect 25041 5692 25053 5695
rect 25004 5664 25053 5692
rect 25004 5652 25010 5664
rect 25041 5661 25053 5664
rect 25087 5661 25099 5695
rect 25041 5655 25099 5661
rect 25406 5652 25412 5704
rect 25464 5692 25470 5704
rect 25700 5701 25728 5732
rect 26050 5720 26056 5732
rect 26108 5720 26114 5772
rect 25685 5695 25743 5701
rect 25685 5692 25697 5695
rect 25464 5664 25697 5692
rect 25464 5652 25470 5664
rect 25685 5661 25697 5664
rect 25731 5661 25743 5695
rect 27338 5692 27344 5704
rect 27094 5664 27344 5692
rect 25685 5655 25743 5661
rect 27338 5652 27344 5664
rect 27396 5652 27402 5704
rect 27448 5692 27476 5788
rect 33152 5772 33180 5800
rect 33778 5788 33784 5800
rect 33836 5788 33842 5840
rect 27798 5720 27804 5772
rect 27856 5760 27862 5772
rect 27985 5763 28043 5769
rect 27985 5760 27997 5763
rect 27856 5732 27997 5760
rect 27856 5720 27862 5732
rect 27985 5729 27997 5732
rect 28031 5729 28043 5763
rect 27985 5723 28043 5729
rect 28074 5720 28080 5772
rect 28132 5760 28138 5772
rect 28169 5763 28227 5769
rect 28169 5760 28181 5763
rect 28132 5732 28181 5760
rect 28132 5720 28138 5732
rect 28169 5729 28181 5732
rect 28215 5729 28227 5763
rect 28169 5723 28227 5729
rect 27893 5695 27951 5701
rect 27893 5692 27905 5695
rect 27448 5664 27905 5692
rect 27893 5661 27905 5664
rect 27939 5661 27951 5695
rect 28184 5692 28212 5723
rect 30282 5720 30288 5772
rect 30340 5760 30346 5772
rect 30653 5763 30711 5769
rect 30653 5760 30665 5763
rect 30340 5732 30665 5760
rect 30340 5720 30346 5732
rect 30653 5729 30665 5732
rect 30699 5729 30711 5763
rect 30653 5723 30711 5729
rect 30837 5763 30895 5769
rect 30837 5729 30849 5763
rect 30883 5760 30895 5763
rect 31021 5763 31079 5769
rect 31021 5760 31033 5763
rect 30883 5732 31033 5760
rect 30883 5729 30895 5732
rect 30837 5723 30895 5729
rect 31021 5729 31033 5732
rect 31067 5760 31079 5763
rect 32306 5760 32312 5772
rect 31067 5732 32312 5760
rect 31067 5729 31079 5732
rect 31021 5723 31079 5729
rect 32306 5720 32312 5732
rect 32364 5720 32370 5772
rect 33134 5720 33140 5772
rect 33192 5720 33198 5772
rect 33321 5763 33379 5769
rect 33321 5729 33333 5763
rect 33367 5760 33379 5763
rect 34701 5763 34759 5769
rect 34701 5760 34713 5763
rect 33367 5732 34713 5760
rect 33367 5729 33379 5732
rect 33321 5723 33379 5729
rect 34701 5729 34713 5732
rect 34747 5729 34759 5763
rect 34701 5723 34759 5729
rect 28445 5695 28503 5701
rect 28445 5692 28457 5695
rect 28184 5664 28457 5692
rect 27893 5655 27951 5661
rect 28445 5661 28457 5664
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 28460 5624 28488 5655
rect 28534 5652 28540 5704
rect 28592 5652 28598 5704
rect 31110 5652 31116 5704
rect 31168 5692 31174 5704
rect 31297 5695 31355 5701
rect 31297 5692 31309 5695
rect 31168 5664 31309 5692
rect 31168 5652 31174 5664
rect 31297 5661 31309 5664
rect 31343 5661 31355 5695
rect 31297 5655 31355 5661
rect 33226 5652 33232 5704
rect 33284 5652 33290 5704
rect 33410 5652 33416 5704
rect 33468 5652 33474 5704
rect 33689 5695 33747 5701
rect 33689 5692 33701 5695
rect 33612 5664 33701 5692
rect 29822 5624 29828 5636
rect 28460 5596 29828 5624
rect 29822 5584 29828 5596
rect 29880 5624 29886 5636
rect 29880 5596 30604 5624
rect 29880 5584 29886 5596
rect 21600 5528 23704 5556
rect 28721 5559 28779 5565
rect 21600 5516 21606 5528
rect 28721 5525 28733 5559
rect 28767 5556 28779 5559
rect 29546 5556 29552 5568
rect 28767 5528 29552 5556
rect 28767 5525 28779 5528
rect 28721 5519 28779 5525
rect 29546 5516 29552 5528
rect 29604 5516 29610 5568
rect 30576 5565 30604 5596
rect 33318 5584 33324 5636
rect 33376 5624 33382 5636
rect 33612 5624 33640 5664
rect 33689 5661 33701 5664
rect 33735 5661 33747 5695
rect 33689 5655 33747 5661
rect 33778 5652 33784 5704
rect 33836 5692 33842 5704
rect 33965 5695 34023 5701
rect 33965 5692 33977 5695
rect 33836 5664 33977 5692
rect 33836 5652 33842 5664
rect 33965 5661 33977 5664
rect 34011 5661 34023 5695
rect 33965 5655 34023 5661
rect 34514 5624 34520 5636
rect 33376 5596 34520 5624
rect 33376 5584 33382 5596
rect 34514 5584 34520 5596
rect 34572 5584 34578 5636
rect 34885 5627 34943 5633
rect 34885 5593 34897 5627
rect 34931 5624 34943 5627
rect 35066 5624 35072 5636
rect 34931 5596 35072 5624
rect 34931 5593 34943 5596
rect 34885 5587 34943 5593
rect 35066 5584 35072 5596
rect 35124 5584 35130 5636
rect 30561 5559 30619 5565
rect 30561 5525 30573 5559
rect 30607 5556 30619 5559
rect 36170 5556 36176 5568
rect 30607 5528 36176 5556
rect 30607 5525 30619 5528
rect 30561 5519 30619 5525
rect 36170 5516 36176 5528
rect 36228 5516 36234 5568
rect 1104 5466 37076 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 37076 5466
rect 1104 5392 37076 5414
rect 15838 5312 15844 5364
rect 15896 5312 15902 5364
rect 23106 5352 23112 5364
rect 18984 5324 23112 5352
rect 14366 5244 14372 5296
rect 14424 5244 14430 5296
rect 15654 5284 15660 5296
rect 15594 5256 15660 5284
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 16850 5244 16856 5296
rect 16908 5284 16914 5296
rect 16945 5287 17003 5293
rect 16945 5284 16957 5287
rect 16908 5256 16957 5284
rect 16908 5244 16914 5256
rect 16945 5253 16957 5256
rect 16991 5253 17003 5287
rect 18138 5284 18144 5296
rect 16945 5247 17003 5253
rect 17420 5256 18144 5284
rect 14090 5176 14096 5228
rect 14148 5176 14154 5228
rect 17420 5225 17448 5256
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17589 5219 17647 5225
rect 17589 5185 17601 5219
rect 17635 5185 17647 5219
rect 17589 5179 17647 5185
rect 17681 5219 17739 5225
rect 17681 5185 17693 5219
rect 17727 5216 17739 5219
rect 18322 5216 18328 5228
rect 17727 5188 18328 5216
rect 17727 5185 17739 5188
rect 17681 5179 17739 5185
rect 16758 5108 16764 5160
rect 16816 5148 16822 5160
rect 17604 5148 17632 5179
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 18984 5225 19012 5324
rect 23106 5312 23112 5324
rect 23164 5352 23170 5364
rect 28166 5352 28172 5364
rect 23164 5324 23612 5352
rect 23164 5312 23170 5324
rect 23290 5244 23296 5296
rect 23348 5244 23354 5296
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5185 19027 5219
rect 20530 5216 20536 5228
rect 20378 5188 20536 5216
rect 18969 5179 19027 5185
rect 20530 5176 20536 5188
rect 20588 5216 20594 5228
rect 22278 5216 22284 5228
rect 20588 5188 22284 5216
rect 20588 5176 20594 5188
rect 16816 5120 17632 5148
rect 19245 5151 19303 5157
rect 16816 5108 16822 5120
rect 19245 5117 19257 5151
rect 19291 5148 19303 5151
rect 20806 5148 20812 5160
rect 19291 5120 20812 5148
rect 19291 5117 19303 5120
rect 19245 5111 19303 5117
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 21821 5151 21879 5157
rect 21821 5117 21833 5151
rect 21867 5148 21879 5151
rect 22094 5148 22100 5160
rect 21867 5120 22100 5148
rect 21867 5117 21879 5120
rect 21821 5111 21879 5117
rect 22094 5108 22100 5120
rect 22152 5108 22158 5160
rect 22204 5148 22232 5188
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 23584 5225 23612 5324
rect 23676 5324 24808 5352
rect 23569 5219 23627 5225
rect 23569 5185 23581 5219
rect 23615 5185 23627 5219
rect 23569 5179 23627 5185
rect 23676 5148 23704 5324
rect 24670 5244 24676 5296
rect 24728 5284 24734 5296
rect 24780 5284 24808 5324
rect 27080 5324 28172 5352
rect 27080 5284 27108 5324
rect 28166 5312 28172 5324
rect 28224 5312 28230 5364
rect 28534 5312 28540 5364
rect 28592 5352 28598 5364
rect 28721 5355 28779 5361
rect 28721 5352 28733 5355
rect 28592 5324 28733 5352
rect 28592 5312 28598 5324
rect 28721 5321 28733 5324
rect 28767 5321 28779 5355
rect 30006 5352 30012 5364
rect 28721 5315 28779 5321
rect 29840 5324 30012 5352
rect 24728 5256 24808 5284
rect 26988 5256 27108 5284
rect 24728 5244 24734 5256
rect 25406 5176 25412 5228
rect 25464 5176 25470 5228
rect 26988 5225 27016 5256
rect 27154 5244 27160 5296
rect 27212 5284 27218 5296
rect 27249 5287 27307 5293
rect 27249 5284 27261 5287
rect 27212 5256 27261 5284
rect 27212 5244 27218 5256
rect 27249 5253 27261 5256
rect 27295 5253 27307 5287
rect 29730 5284 29736 5296
rect 28474 5256 29736 5284
rect 27249 5247 27307 5253
rect 29730 5244 29736 5256
rect 29788 5244 29794 5296
rect 29840 5293 29868 5324
rect 30006 5312 30012 5324
rect 30064 5312 30070 5364
rect 30098 5312 30104 5364
rect 30156 5352 30162 5364
rect 32306 5361 32312 5364
rect 30193 5355 30251 5361
rect 30193 5352 30205 5355
rect 30156 5324 30205 5352
rect 30156 5312 30162 5324
rect 30193 5321 30205 5324
rect 30239 5321 30251 5355
rect 30193 5315 30251 5321
rect 32293 5355 32312 5361
rect 32293 5321 32305 5355
rect 32293 5315 32312 5321
rect 32306 5312 32312 5315
rect 32364 5312 32370 5364
rect 29825 5287 29883 5293
rect 29825 5253 29837 5287
rect 29871 5253 29883 5287
rect 29825 5247 29883 5253
rect 29914 5244 29920 5296
rect 29972 5244 29978 5296
rect 30024 5284 30052 5312
rect 30024 5256 30328 5284
rect 26973 5219 27031 5225
rect 26973 5185 26985 5219
rect 27019 5185 27031 5219
rect 26973 5179 27031 5185
rect 29546 5176 29552 5228
rect 29604 5176 29610 5228
rect 29642 5219 29700 5225
rect 29642 5185 29654 5219
rect 29688 5185 29700 5219
rect 29642 5179 29700 5185
rect 30055 5219 30113 5225
rect 30055 5185 30067 5219
rect 30101 5216 30113 5219
rect 30190 5216 30196 5228
rect 30101 5188 30196 5216
rect 30101 5185 30113 5188
rect 30055 5179 30113 5185
rect 22204 5120 23704 5148
rect 24394 5108 24400 5160
rect 24452 5148 24458 5160
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 24452 5120 25145 5148
rect 24452 5108 24458 5120
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 29656 5148 29684 5179
rect 30190 5176 30196 5188
rect 30248 5176 30254 5228
rect 30300 5225 30328 5256
rect 30374 5244 30380 5296
rect 30432 5284 30438 5296
rect 30432 5256 31524 5284
rect 30432 5244 30438 5256
rect 30285 5219 30343 5225
rect 30285 5185 30297 5219
rect 30331 5185 30343 5219
rect 30285 5179 30343 5185
rect 30469 5219 30527 5225
rect 30469 5185 30481 5219
rect 30515 5185 30527 5219
rect 30469 5179 30527 5185
rect 25133 5111 25191 5117
rect 26206 5120 29684 5148
rect 20717 5083 20775 5089
rect 20717 5049 20729 5083
rect 20763 5080 20775 5083
rect 21726 5080 21732 5092
rect 20763 5052 21732 5080
rect 20763 5049 20775 5052
rect 20717 5043 20775 5049
rect 21726 5040 21732 5052
rect 21784 5040 21790 5092
rect 23661 5015 23719 5021
rect 23661 4981 23673 5015
rect 23707 5012 23719 5015
rect 23842 5012 23848 5024
rect 23707 4984 23848 5012
rect 23707 4981 23719 4984
rect 23661 4975 23719 4981
rect 23842 4972 23848 4984
rect 23900 5012 23906 5024
rect 24486 5012 24492 5024
rect 23900 4984 24492 5012
rect 23900 4972 23906 4984
rect 24486 4972 24492 4984
rect 24544 4972 24550 5024
rect 24946 4972 24952 5024
rect 25004 5012 25010 5024
rect 26206 5012 26234 5120
rect 30484 5092 30512 5179
rect 30834 5176 30840 5228
rect 30892 5176 30898 5228
rect 31018 5176 31024 5228
rect 31076 5176 31082 5228
rect 31110 5176 31116 5228
rect 31168 5176 31174 5228
rect 31496 5225 31524 5256
rect 32490 5244 32496 5296
rect 32548 5244 32554 5296
rect 33318 5284 33324 5296
rect 32968 5256 33324 5284
rect 32968 5225 32996 5256
rect 33318 5244 33324 5256
rect 33376 5244 33382 5296
rect 34241 5287 34299 5293
rect 34241 5284 34253 5287
rect 34164 5256 34253 5284
rect 31389 5219 31447 5225
rect 31389 5185 31401 5219
rect 31435 5185 31447 5219
rect 31389 5179 31447 5185
rect 31481 5219 31539 5225
rect 31481 5185 31493 5219
rect 31527 5185 31539 5219
rect 31481 5179 31539 5185
rect 32953 5219 33011 5225
rect 32953 5185 32965 5219
rect 32999 5185 33011 5219
rect 32953 5179 33011 5185
rect 30653 5151 30711 5157
rect 30653 5117 30665 5151
rect 30699 5148 30711 5151
rect 31404 5148 31432 5179
rect 33134 5176 33140 5228
rect 33192 5176 33198 5228
rect 33410 5176 33416 5228
rect 33468 5176 33474 5228
rect 34164 5225 34192 5256
rect 34241 5253 34253 5256
rect 34287 5284 34299 5287
rect 35066 5284 35072 5296
rect 34287 5256 35072 5284
rect 34287 5253 34299 5256
rect 34241 5247 34299 5253
rect 35066 5244 35072 5256
rect 35124 5244 35130 5296
rect 34149 5219 34207 5225
rect 34149 5185 34161 5219
rect 34195 5185 34207 5219
rect 34149 5179 34207 5185
rect 34698 5176 34704 5228
rect 34756 5176 34762 5228
rect 34882 5176 34888 5228
rect 34940 5176 34946 5228
rect 35161 5219 35219 5225
rect 35161 5216 35173 5219
rect 34992 5188 35173 5216
rect 30699 5120 31432 5148
rect 30699 5117 30711 5120
rect 30653 5111 30711 5117
rect 34054 5108 34060 5160
rect 34112 5108 34118 5160
rect 34422 5108 34428 5160
rect 34480 5148 34486 5160
rect 34793 5151 34851 5157
rect 34793 5148 34805 5151
rect 34480 5120 34805 5148
rect 34480 5108 34486 5120
rect 34793 5117 34805 5120
rect 34839 5117 34851 5151
rect 34793 5111 34851 5117
rect 30466 5040 30472 5092
rect 30524 5080 30530 5092
rect 32125 5083 32183 5089
rect 32125 5080 32137 5083
rect 30524 5052 32137 5080
rect 30524 5040 30530 5052
rect 32125 5049 32137 5052
rect 32171 5049 32183 5083
rect 32125 5043 32183 5049
rect 34330 5040 34336 5092
rect 34388 5080 34394 5092
rect 34992 5080 35020 5188
rect 35161 5185 35173 5188
rect 35207 5185 35219 5219
rect 35161 5179 35219 5185
rect 34388 5052 35020 5080
rect 34388 5040 34394 5052
rect 25004 4984 26234 5012
rect 25004 4972 25010 4984
rect 30650 4972 30656 5024
rect 30708 5012 30714 5024
rect 31205 5015 31263 5021
rect 31205 5012 31217 5015
rect 30708 4984 31217 5012
rect 30708 4972 30714 4984
rect 31205 4981 31217 4984
rect 31251 4981 31263 5015
rect 31205 4975 31263 4981
rect 32306 4972 32312 5024
rect 32364 4972 32370 5024
rect 33226 4972 33232 5024
rect 33284 5012 33290 5024
rect 34790 5012 34796 5024
rect 33284 4984 34796 5012
rect 33284 4972 33290 4984
rect 34790 4972 34796 4984
rect 34848 4972 34854 5024
rect 35161 5015 35219 5021
rect 35161 4981 35173 5015
rect 35207 5012 35219 5015
rect 35526 5012 35532 5024
rect 35207 4984 35532 5012
rect 35207 4981 35219 4984
rect 35161 4975 35219 4981
rect 35526 4972 35532 4984
rect 35584 4972 35590 5024
rect 1104 4922 37076 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 37076 4922
rect 1104 4848 37076 4870
rect 16758 4768 16764 4820
rect 16816 4808 16822 4820
rect 17037 4811 17095 4817
rect 17037 4808 17049 4811
rect 16816 4780 17049 4808
rect 16816 4768 16822 4780
rect 17037 4777 17049 4780
rect 17083 4777 17095 4811
rect 17037 4771 17095 4777
rect 35253 4811 35311 4817
rect 35253 4777 35265 4811
rect 35299 4808 35311 4811
rect 35529 4811 35587 4817
rect 35529 4808 35541 4811
rect 35299 4780 35541 4808
rect 35299 4777 35311 4780
rect 35253 4771 35311 4777
rect 35529 4777 35541 4780
rect 35575 4777 35587 4811
rect 35529 4771 35587 4777
rect 21542 4740 21548 4752
rect 21284 4712 21548 4740
rect 14090 4632 14096 4684
rect 14148 4672 14154 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 14148 4644 15301 4672
rect 14148 4632 14154 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 15562 4632 15568 4684
rect 15620 4632 15626 4684
rect 20806 4632 20812 4684
rect 20864 4632 20870 4684
rect 21284 4613 21312 4712
rect 21542 4700 21548 4712
rect 21600 4700 21606 4752
rect 30374 4700 30380 4752
rect 30432 4700 30438 4752
rect 32306 4740 32312 4752
rect 31864 4712 32312 4740
rect 22094 4672 22100 4684
rect 21468 4644 22100 4672
rect 21468 4613 21496 4644
rect 22094 4632 22100 4644
rect 22152 4632 22158 4684
rect 24394 4632 24400 4684
rect 24452 4632 24458 4684
rect 24486 4632 24492 4684
rect 24544 4672 24550 4684
rect 25133 4675 25191 4681
rect 25133 4672 25145 4675
rect 24544 4644 25145 4672
rect 24544 4632 24550 4644
rect 25133 4641 25145 4644
rect 25179 4641 25191 4675
rect 30392 4672 30420 4700
rect 25133 4635 25191 4641
rect 30300 4644 30420 4672
rect 21269 4607 21327 4613
rect 21269 4573 21281 4607
rect 21315 4573 21327 4607
rect 21269 4567 21327 4573
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4573 21511 4607
rect 21453 4567 21511 4573
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4604 21603 4607
rect 21726 4604 21732 4616
rect 21591 4576 21732 4604
rect 21591 4573 21603 4576
rect 21545 4567 21603 4573
rect 21726 4564 21732 4576
rect 21784 4564 21790 4616
rect 24857 4607 24915 4613
rect 24857 4573 24869 4607
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 15654 4496 15660 4548
rect 15712 4536 15718 4548
rect 24872 4536 24900 4567
rect 25038 4564 25044 4616
rect 25096 4564 25102 4616
rect 30300 4613 30328 4644
rect 30834 4632 30840 4684
rect 30892 4672 30898 4684
rect 31864 4681 31892 4712
rect 32306 4700 32312 4712
rect 32364 4740 32370 4752
rect 34057 4743 34115 4749
rect 34057 4740 34069 4743
rect 32364 4712 34069 4740
rect 32364 4700 32370 4712
rect 34057 4709 34069 4712
rect 34103 4709 34115 4743
rect 34057 4703 34115 4709
rect 34698 4700 34704 4752
rect 34756 4740 34762 4752
rect 34756 4712 35112 4740
rect 34756 4700 34762 4712
rect 31573 4675 31631 4681
rect 31573 4672 31585 4675
rect 30892 4644 31585 4672
rect 30892 4632 30898 4644
rect 31573 4641 31585 4644
rect 31619 4641 31631 4675
rect 31573 4635 31631 4641
rect 31849 4675 31907 4681
rect 31849 4641 31861 4675
rect 31895 4641 31907 4675
rect 31849 4635 31907 4641
rect 31938 4632 31944 4684
rect 31996 4672 32002 4684
rect 32585 4675 32643 4681
rect 32585 4672 32597 4675
rect 31996 4644 32597 4672
rect 31996 4632 32002 4644
rect 32585 4641 32597 4644
rect 32631 4641 32643 4675
rect 34422 4672 34428 4684
rect 32585 4635 32643 4641
rect 33520 4644 34428 4672
rect 30101 4607 30159 4613
rect 30101 4573 30113 4607
rect 30147 4573 30159 4607
rect 30101 4567 30159 4573
rect 30285 4607 30343 4613
rect 30285 4573 30297 4607
rect 30331 4573 30343 4607
rect 30285 4567 30343 4573
rect 30377 4607 30435 4613
rect 30377 4573 30389 4607
rect 30423 4604 30435 4607
rect 30466 4604 30472 4616
rect 30423 4576 30472 4604
rect 30423 4573 30435 4576
rect 30377 4567 30435 4573
rect 25314 4536 25320 4548
rect 15712 4508 16054 4536
rect 24872 4508 25320 4536
rect 15712 4496 15718 4508
rect 25314 4496 25320 4508
rect 25372 4496 25378 4548
rect 29454 4496 29460 4548
rect 29512 4536 29518 4548
rect 29641 4539 29699 4545
rect 29641 4536 29653 4539
rect 29512 4508 29653 4536
rect 29512 4496 29518 4508
rect 29641 4505 29653 4508
rect 29687 4505 29699 4539
rect 30116 4536 30144 4567
rect 30466 4564 30472 4576
rect 30524 4564 30530 4616
rect 32030 4564 32036 4616
rect 32088 4604 32094 4616
rect 32125 4607 32183 4613
rect 32125 4604 32137 4607
rect 32088 4576 32137 4604
rect 32088 4564 32094 4576
rect 32125 4573 32137 4576
rect 32171 4573 32183 4607
rect 32125 4567 32183 4573
rect 32217 4607 32275 4613
rect 32217 4573 32229 4607
rect 32263 4604 32275 4607
rect 33134 4604 33140 4616
rect 32263 4576 33140 4604
rect 32263 4573 32275 4576
rect 32217 4567 32275 4573
rect 30116 4508 30420 4536
rect 29641 4499 29699 4505
rect 30392 4480 30420 4508
rect 31018 4496 31024 4548
rect 31076 4536 31082 4548
rect 32232 4536 32260 4567
rect 33134 4564 33140 4576
rect 33192 4564 33198 4616
rect 33226 4564 33232 4616
rect 33284 4564 33290 4616
rect 33318 4564 33324 4616
rect 33376 4604 33382 4616
rect 33520 4613 33548 4644
rect 34422 4632 34428 4644
rect 34480 4672 34486 4684
rect 35084 4681 35112 4712
rect 34977 4675 35035 4681
rect 34977 4672 34989 4675
rect 34480 4644 34989 4672
rect 34480 4632 34486 4644
rect 34977 4641 34989 4644
rect 35023 4641 35035 4675
rect 34977 4635 35035 4641
rect 35069 4675 35127 4681
rect 35069 4641 35081 4675
rect 35115 4641 35127 4675
rect 35069 4635 35127 4641
rect 33505 4607 33563 4613
rect 33505 4604 33517 4607
rect 33376 4576 33517 4604
rect 33376 4564 33382 4576
rect 33505 4573 33517 4576
rect 33551 4573 33563 4607
rect 33505 4567 33563 4573
rect 33597 4607 33655 4613
rect 33597 4573 33609 4607
rect 33643 4604 33655 4607
rect 33686 4604 33692 4616
rect 33643 4576 33692 4604
rect 33643 4573 33655 4576
rect 33597 4567 33655 4573
rect 33686 4564 33692 4576
rect 33744 4564 33750 4616
rect 34793 4607 34851 4613
rect 34793 4573 34805 4607
rect 34839 4573 34851 4607
rect 34793 4567 34851 4573
rect 31076 4508 32260 4536
rect 31076 4496 31082 4508
rect 33410 4496 33416 4548
rect 33468 4536 33474 4548
rect 34330 4536 34336 4548
rect 33468 4508 34336 4536
rect 33468 4496 33474 4508
rect 34330 4496 34336 4508
rect 34388 4536 34394 4548
rect 34808 4536 34836 4567
rect 34882 4564 34888 4616
rect 34940 4564 34946 4616
rect 35342 4564 35348 4616
rect 35400 4604 35406 4616
rect 35400 4576 35756 4604
rect 35400 4564 35406 4576
rect 35526 4545 35532 4548
rect 34388 4508 34836 4536
rect 35513 4539 35532 4545
rect 34388 4496 34394 4508
rect 35513 4505 35525 4539
rect 35513 4499 35532 4505
rect 35526 4496 35532 4499
rect 35584 4496 35590 4548
rect 35728 4545 35756 4576
rect 35713 4539 35771 4545
rect 35713 4505 35725 4539
rect 35759 4505 35771 4539
rect 35713 4499 35771 4505
rect 30374 4428 30380 4480
rect 30432 4428 30438 4480
rect 31294 4428 31300 4480
rect 31352 4468 31358 4480
rect 31941 4471 31999 4477
rect 31941 4468 31953 4471
rect 31352 4440 31953 4468
rect 31352 4428 31358 4440
rect 31941 4437 31953 4440
rect 31987 4437 31999 4471
rect 31941 4431 31999 4437
rect 32306 4428 32312 4480
rect 32364 4428 32370 4480
rect 32490 4428 32496 4480
rect 32548 4428 32554 4480
rect 35342 4428 35348 4480
rect 35400 4428 35406 4480
rect 1104 4378 37076 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 37076 4378
rect 1104 4304 37076 4326
rect 30374 4224 30380 4276
rect 30432 4224 30438 4276
rect 31097 4267 31155 4273
rect 31097 4233 31109 4267
rect 31143 4264 31155 4267
rect 31754 4264 31760 4276
rect 31143 4236 31760 4264
rect 31143 4233 31155 4236
rect 31097 4227 31155 4233
rect 31754 4224 31760 4236
rect 31812 4224 31818 4276
rect 31849 4267 31907 4273
rect 31849 4233 31861 4267
rect 31895 4264 31907 4267
rect 31938 4264 31944 4276
rect 31895 4236 31944 4264
rect 31895 4233 31907 4236
rect 31849 4227 31907 4233
rect 31938 4224 31944 4236
rect 31996 4224 32002 4276
rect 32217 4267 32275 4273
rect 32217 4233 32229 4267
rect 32263 4264 32275 4267
rect 32306 4264 32312 4276
rect 32263 4236 32312 4264
rect 32263 4233 32275 4236
rect 32217 4227 32275 4233
rect 32306 4224 32312 4236
rect 32364 4224 32370 4276
rect 32398 4224 32404 4276
rect 32456 4264 32462 4276
rect 32456 4236 33180 4264
rect 32456 4224 32462 4236
rect 30282 4196 30288 4208
rect 29946 4168 30288 4196
rect 30282 4156 30288 4168
rect 30340 4196 30346 4208
rect 30340 4168 30420 4196
rect 30340 4156 30346 4168
rect 28166 4088 28172 4140
rect 28224 4128 28230 4140
rect 28445 4131 28503 4137
rect 28445 4128 28457 4131
rect 28224 4100 28457 4128
rect 28224 4088 28230 4100
rect 28445 4097 28457 4100
rect 28491 4097 28503 4131
rect 30392 4128 30420 4168
rect 31294 4156 31300 4208
rect 31352 4156 31358 4208
rect 32030 4156 32036 4208
rect 32088 4196 32094 4208
rect 33152 4205 33180 4236
rect 33318 4224 33324 4276
rect 33376 4224 33382 4276
rect 33410 4224 33416 4276
rect 33468 4264 33474 4276
rect 33597 4267 33655 4273
rect 33597 4264 33609 4267
rect 33468 4236 33609 4264
rect 33468 4224 33474 4236
rect 33597 4233 33609 4236
rect 33643 4233 33655 4267
rect 33597 4227 33655 4233
rect 33045 4199 33103 4205
rect 33045 4196 33057 4199
rect 32088 4168 33057 4196
rect 32088 4156 32094 4168
rect 33045 4165 33057 4168
rect 33091 4165 33103 4199
rect 33045 4159 33103 4165
rect 33137 4199 33195 4205
rect 33137 4165 33149 4199
rect 33183 4196 33195 4199
rect 33686 4196 33692 4208
rect 33183 4168 33692 4196
rect 33183 4165 33195 4168
rect 33137 4159 33195 4165
rect 33686 4156 33692 4168
rect 33744 4156 33750 4208
rect 35069 4199 35127 4205
rect 35069 4165 35081 4199
rect 35115 4196 35127 4199
rect 35342 4196 35348 4208
rect 35115 4168 35348 4196
rect 35115 4165 35127 4168
rect 35069 4159 35127 4165
rect 35342 4156 35348 4168
rect 35400 4156 35406 4208
rect 30742 4128 30748 4140
rect 30392 4100 30748 4128
rect 28445 4091 28503 4097
rect 30742 4088 30748 4100
rect 30800 4088 30806 4140
rect 32490 4128 32496 4140
rect 30852 4100 32496 4128
rect 28721 4063 28779 4069
rect 28721 4029 28733 4063
rect 28767 4060 28779 4063
rect 29454 4060 29460 4072
rect 28767 4032 29460 4060
rect 28767 4029 28779 4032
rect 28721 4023 28779 4029
rect 29454 4020 29460 4032
rect 29512 4020 29518 4072
rect 30852 4069 30880 4100
rect 32490 4088 32496 4100
rect 32548 4128 32554 4140
rect 32769 4131 32827 4137
rect 32769 4128 32781 4131
rect 32548 4100 32781 4128
rect 32548 4088 32554 4100
rect 32769 4097 32781 4100
rect 32815 4097 32827 4131
rect 32769 4091 32827 4097
rect 32953 4131 33011 4137
rect 32953 4097 32965 4131
rect 32999 4097 33011 4131
rect 32953 4091 33011 4097
rect 30193 4063 30251 4069
rect 30193 4029 30205 4063
rect 30239 4060 30251 4063
rect 30837 4063 30895 4069
rect 30837 4060 30849 4063
rect 30239 4032 30849 4060
rect 30239 4029 30251 4032
rect 30193 4023 30251 4029
rect 30837 4029 30849 4032
rect 30883 4029 30895 4063
rect 30837 4023 30895 4029
rect 31389 4063 31447 4069
rect 31389 4029 31401 4063
rect 31435 4060 31447 4063
rect 31846 4060 31852 4072
rect 31435 4032 31852 4060
rect 31435 4029 31447 4032
rect 31389 4023 31447 4029
rect 31846 4020 31852 4032
rect 31904 4060 31910 4072
rect 32398 4060 32404 4072
rect 31904 4032 32404 4060
rect 31904 4020 31910 4032
rect 32398 4020 32404 4032
rect 32456 4020 32462 4072
rect 32674 4020 32680 4072
rect 32732 4060 32738 4072
rect 32968 4060 32996 4091
rect 33962 4088 33968 4140
rect 34020 4088 34026 4140
rect 32732 4032 32996 4060
rect 32732 4020 32738 4032
rect 33042 4020 33048 4072
rect 33100 4060 33106 4072
rect 35345 4063 35403 4069
rect 35345 4060 35357 4063
rect 33100 4032 35357 4060
rect 33100 4020 33106 4032
rect 35345 4029 35357 4032
rect 35391 4029 35403 4063
rect 35345 4023 35403 4029
rect 30466 3884 30472 3936
rect 30524 3924 30530 3936
rect 30929 3927 30987 3933
rect 30929 3924 30941 3927
rect 30524 3896 30941 3924
rect 30524 3884 30530 3896
rect 30929 3893 30941 3896
rect 30975 3893 30987 3927
rect 30929 3887 30987 3893
rect 31113 3927 31171 3933
rect 31113 3893 31125 3927
rect 31159 3924 31171 3927
rect 33594 3924 33600 3936
rect 31159 3896 33600 3924
rect 31159 3893 31171 3896
rect 31113 3887 31171 3893
rect 33594 3884 33600 3896
rect 33652 3884 33658 3936
rect 1104 3834 37076 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 37076 3834
rect 1104 3760 37076 3782
rect 31754 3680 31760 3732
rect 31812 3720 31818 3732
rect 32493 3723 32551 3729
rect 32493 3720 32505 3723
rect 31812 3692 32505 3720
rect 31812 3680 31818 3692
rect 32493 3689 32505 3692
rect 32539 3720 32551 3723
rect 32950 3720 32956 3732
rect 32539 3692 32956 3720
rect 32539 3689 32551 3692
rect 32493 3683 32551 3689
rect 32950 3680 32956 3692
rect 33008 3680 33014 3732
rect 33594 3612 33600 3664
rect 33652 3652 33658 3664
rect 33652 3624 34008 3652
rect 33652 3612 33658 3624
rect 30285 3587 30343 3593
rect 30285 3553 30297 3587
rect 30331 3584 30343 3587
rect 30650 3584 30656 3596
rect 30331 3556 30656 3584
rect 30331 3553 30343 3556
rect 30285 3547 30343 3553
rect 30650 3544 30656 3556
rect 30708 3544 30714 3596
rect 31757 3587 31815 3593
rect 31757 3553 31769 3587
rect 31803 3584 31815 3587
rect 31846 3584 31852 3596
rect 31803 3556 31852 3584
rect 31803 3553 31815 3556
rect 31757 3547 31815 3553
rect 31846 3544 31852 3556
rect 31904 3544 31910 3596
rect 32677 3587 32735 3593
rect 32677 3584 32689 3587
rect 32140 3556 32689 3584
rect 30006 3476 30012 3528
rect 30064 3476 30070 3528
rect 32140 3525 32168 3556
rect 32677 3553 32689 3556
rect 32723 3553 32735 3587
rect 33226 3584 33232 3596
rect 32677 3547 32735 3553
rect 32876 3556 33232 3584
rect 32125 3519 32183 3525
rect 32125 3485 32137 3519
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 32401 3519 32459 3525
rect 32401 3485 32413 3519
rect 32447 3485 32459 3519
rect 32401 3479 32459 3485
rect 32585 3519 32643 3525
rect 32585 3485 32597 3519
rect 32631 3516 32643 3519
rect 32876 3516 32904 3556
rect 33226 3544 33232 3556
rect 33284 3544 33290 3596
rect 33873 3587 33931 3593
rect 33873 3584 33885 3587
rect 33336 3556 33885 3584
rect 32631 3488 32904 3516
rect 32631 3485 32643 3488
rect 32585 3479 32643 3485
rect 30926 3408 30932 3460
rect 30984 3408 30990 3460
rect 32416 3448 32444 3479
rect 32950 3476 32956 3528
rect 33008 3516 33014 3528
rect 33336 3525 33364 3556
rect 33873 3553 33885 3556
rect 33919 3553 33931 3587
rect 33873 3547 33931 3553
rect 33980 3525 34008 3624
rect 33137 3519 33195 3525
rect 33137 3516 33149 3519
rect 33008 3488 33149 3516
rect 33008 3476 33014 3488
rect 33137 3485 33149 3488
rect 33183 3485 33195 3519
rect 33137 3479 33195 3485
rect 33321 3519 33379 3525
rect 33321 3485 33333 3519
rect 33367 3485 33379 3519
rect 33321 3479 33379 3485
rect 33413 3519 33471 3525
rect 33413 3485 33425 3519
rect 33459 3516 33471 3519
rect 33781 3519 33839 3525
rect 33781 3516 33793 3519
rect 33459 3488 33793 3516
rect 33459 3485 33471 3488
rect 33413 3479 33471 3485
rect 33781 3485 33793 3488
rect 33827 3485 33839 3519
rect 33781 3479 33839 3485
rect 33965 3519 34023 3525
rect 33965 3485 33977 3519
rect 34011 3485 34023 3519
rect 33965 3479 34023 3485
rect 33686 3448 33692 3460
rect 32416 3420 33692 3448
rect 33686 3408 33692 3420
rect 33744 3408 33750 3460
rect 33796 3448 33824 3479
rect 34698 3448 34704 3460
rect 33796 3420 34704 3448
rect 34698 3408 34704 3420
rect 34756 3408 34762 3460
rect 32033 3383 32091 3389
rect 32033 3349 32045 3383
rect 32079 3380 32091 3383
rect 32398 3380 32404 3392
rect 32079 3352 32404 3380
rect 32079 3349 32091 3352
rect 32033 3343 32091 3349
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 1104 3290 37076 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 37076 3290
rect 1104 3216 37076 3238
rect 33873 3179 33931 3185
rect 33873 3145 33885 3179
rect 33919 3176 33931 3179
rect 34698 3176 34704 3188
rect 33919 3148 34704 3176
rect 33919 3145 33931 3148
rect 33873 3139 33931 3145
rect 34698 3136 34704 3148
rect 34756 3136 34762 3188
rect 30466 3068 30472 3120
rect 30524 3068 30530 3120
rect 30926 3068 30932 3120
rect 30984 3068 30990 3120
rect 32398 3068 32404 3120
rect 32456 3068 32462 3120
rect 33962 3108 33968 3120
rect 33626 3080 33968 3108
rect 33962 3068 33968 3080
rect 34020 3068 34026 3120
rect 30006 2932 30012 2984
rect 30064 2972 30070 2984
rect 30193 2975 30251 2981
rect 30193 2972 30205 2975
rect 30064 2944 30205 2972
rect 30064 2932 30070 2944
rect 30193 2941 30205 2944
rect 30239 2972 30251 2975
rect 31941 2975 31999 2981
rect 30239 2944 31892 2972
rect 30239 2941 30251 2944
rect 30193 2935 30251 2941
rect 31864 2904 31892 2944
rect 31941 2941 31953 2975
rect 31987 2972 31999 2975
rect 32030 2972 32036 2984
rect 31987 2944 32036 2972
rect 31987 2941 31999 2944
rect 31941 2935 31999 2941
rect 32030 2932 32036 2944
rect 32088 2932 32094 2984
rect 32125 2975 32183 2981
rect 32125 2941 32137 2975
rect 32171 2972 32183 2975
rect 33042 2972 33048 2984
rect 32171 2944 33048 2972
rect 32171 2941 32183 2944
rect 32125 2935 32183 2941
rect 32140 2904 32168 2935
rect 33042 2932 33048 2944
rect 33100 2932 33106 2984
rect 31864 2876 32168 2904
rect 1104 2746 37076 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 37076 2746
rect 1104 2672 37076 2694
rect 23477 2635 23535 2641
rect 23477 2601 23489 2635
rect 23523 2632 23535 2635
rect 24946 2632 24952 2644
rect 23523 2604 24952 2632
rect 23523 2601 23535 2604
rect 23477 2595 23535 2601
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 23256 2400 23305 2428
rect 23256 2388 23262 2400
rect 23293 2397 23305 2400
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 1104 2202 37076 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 37076 2202
rect 1104 2128 37076 2150
<< via1 >>
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 31944 37884 31996 37936
rect 32956 37884 33008 37936
rect 12532 37816 12584 37868
rect 16028 37859 16080 37868
rect 16028 37825 16037 37859
rect 16037 37825 16071 37859
rect 16071 37825 16080 37859
rect 16028 37816 16080 37825
rect 16396 37816 16448 37868
rect 18604 37859 18656 37868
rect 18604 37825 18613 37859
rect 18613 37825 18647 37859
rect 18647 37825 18656 37859
rect 18604 37816 18656 37825
rect 23848 37816 23900 37868
rect 25228 37859 25280 37868
rect 25228 37825 25237 37859
rect 25237 37825 25271 37859
rect 25271 37825 25280 37859
rect 25228 37816 25280 37825
rect 28080 37816 28132 37868
rect 29736 37859 29788 37868
rect 29736 37825 29745 37859
rect 29745 37825 29779 37859
rect 29779 37825 29788 37859
rect 29736 37816 29788 37825
rect 31668 37816 31720 37868
rect 32864 37816 32916 37868
rect 13084 37748 13136 37800
rect 13728 37791 13780 37800
rect 13728 37757 13737 37791
rect 13737 37757 13771 37791
rect 13771 37757 13780 37791
rect 13728 37748 13780 37757
rect 18696 37791 18748 37800
rect 18696 37757 18705 37791
rect 18705 37757 18739 37791
rect 18739 37757 18748 37791
rect 18696 37748 18748 37757
rect 18880 37791 18932 37800
rect 18880 37757 18889 37791
rect 18889 37757 18923 37791
rect 18923 37757 18932 37791
rect 18880 37748 18932 37757
rect 23664 37791 23716 37800
rect 23664 37757 23673 37791
rect 23673 37757 23707 37791
rect 23707 37757 23716 37791
rect 23664 37748 23716 37757
rect 24860 37748 24912 37800
rect 27252 37748 27304 37800
rect 29184 37791 29236 37800
rect 29184 37757 29193 37791
rect 29193 37757 29227 37791
rect 29227 37757 29236 37791
rect 29184 37748 29236 37757
rect 30380 37748 30432 37800
rect 31852 37748 31904 37800
rect 32220 37680 32272 37732
rect 13452 37612 13504 37664
rect 16212 37612 16264 37664
rect 17500 37612 17552 37664
rect 22376 37612 22428 37664
rect 25412 37655 25464 37664
rect 25412 37621 25421 37655
rect 25421 37621 25455 37655
rect 25455 37621 25464 37655
rect 25412 37612 25464 37621
rect 27712 37612 27764 37664
rect 27988 37612 28040 37664
rect 31576 37655 31628 37664
rect 31576 37621 31585 37655
rect 31585 37621 31619 37655
rect 31619 37621 31628 37655
rect 31576 37612 31628 37621
rect 32312 37655 32364 37664
rect 32312 37621 32321 37655
rect 32321 37621 32355 37655
rect 32355 37621 32364 37655
rect 32312 37612 32364 37621
rect 32496 37655 32548 37664
rect 32496 37621 32505 37655
rect 32505 37621 32539 37655
rect 32539 37621 32548 37655
rect 32496 37612 32548 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 15476 37408 15528 37460
rect 16028 37408 16080 37460
rect 18604 37408 18656 37460
rect 23664 37408 23716 37460
rect 24400 37451 24452 37460
rect 24400 37417 24409 37451
rect 24409 37417 24443 37451
rect 24443 37417 24452 37451
rect 24400 37408 24452 37417
rect 28080 37451 28132 37460
rect 28080 37417 28089 37451
rect 28089 37417 28123 37451
rect 28123 37417 28132 37451
rect 28080 37408 28132 37417
rect 31944 37408 31996 37460
rect 23848 37383 23900 37392
rect 23848 37349 23857 37383
rect 23857 37349 23891 37383
rect 23891 37349 23900 37383
rect 23848 37340 23900 37349
rect 13452 37315 13504 37324
rect 13452 37281 13461 37315
rect 13461 37281 13495 37315
rect 13495 37281 13504 37315
rect 13452 37272 13504 37281
rect 16212 37315 16264 37324
rect 16212 37281 16221 37315
rect 16221 37281 16255 37315
rect 16255 37281 16264 37315
rect 16212 37272 16264 37281
rect 17500 37315 17552 37324
rect 17500 37281 17509 37315
rect 17509 37281 17543 37315
rect 17543 37281 17552 37315
rect 17500 37272 17552 37281
rect 21548 37272 21600 37324
rect 22376 37315 22428 37324
rect 22376 37281 22385 37315
rect 22385 37281 22419 37315
rect 22419 37281 22428 37315
rect 22376 37272 22428 37281
rect 848 37204 900 37256
rect 14648 37204 14700 37256
rect 3332 37136 3384 37188
rect 12992 37136 13044 37188
rect 15568 37136 15620 37188
rect 19432 37136 19484 37188
rect 21272 37136 21324 37188
rect 21456 37136 21508 37188
rect 12532 37068 12584 37120
rect 15200 37068 15252 37120
rect 16488 37068 16540 37120
rect 18788 37068 18840 37120
rect 19892 37068 19944 37120
rect 20076 37111 20128 37120
rect 20076 37077 20085 37111
rect 20085 37077 20119 37111
rect 20119 37077 20128 37111
rect 20076 37068 20128 37077
rect 20536 37068 20588 37120
rect 26148 37247 26200 37256
rect 26148 37213 26157 37247
rect 26157 37213 26191 37247
rect 26191 37213 26200 37247
rect 26148 37204 26200 37213
rect 27528 37204 27580 37256
rect 30472 37272 30524 37324
rect 30564 37272 30616 37324
rect 28540 37247 28592 37256
rect 28540 37213 28549 37247
rect 28549 37213 28583 37247
rect 28583 37213 28592 37247
rect 28540 37204 28592 37213
rect 28724 37247 28776 37256
rect 28724 37213 28733 37247
rect 28733 37213 28767 37247
rect 28767 37213 28776 37247
rect 28724 37204 28776 37213
rect 29828 37247 29880 37256
rect 29828 37213 29837 37247
rect 29837 37213 29871 37247
rect 29871 37213 29880 37247
rect 29828 37204 29880 37213
rect 22284 37136 22336 37188
rect 22008 37068 22060 37120
rect 25872 37179 25924 37188
rect 25872 37145 25881 37179
rect 25881 37145 25915 37179
rect 25915 37145 25924 37179
rect 25872 37136 25924 37145
rect 26516 37179 26568 37188
rect 26516 37145 26525 37179
rect 26525 37145 26559 37179
rect 26559 37145 26568 37179
rect 26516 37136 26568 37145
rect 28908 37136 28960 37188
rect 29736 37136 29788 37188
rect 30564 37136 30616 37188
rect 33968 37204 34020 37256
rect 31576 37136 31628 37188
rect 26608 37068 26660 37120
rect 28264 37068 28316 37120
rect 29828 37068 29880 37120
rect 31484 37068 31536 37120
rect 33232 37068 33284 37120
rect 33416 37111 33468 37120
rect 33416 37077 33425 37111
rect 33425 37077 33459 37111
rect 33459 37077 33468 37111
rect 33416 37068 33468 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 12532 36907 12584 36916
rect 12532 36873 12541 36907
rect 12541 36873 12575 36907
rect 12575 36873 12584 36907
rect 12532 36864 12584 36873
rect 16396 36864 16448 36916
rect 18604 36864 18656 36916
rect 18696 36864 18748 36916
rect 12348 36796 12400 36848
rect 12992 36796 13044 36848
rect 15568 36796 15620 36848
rect 12440 36771 12492 36780
rect 12440 36737 12449 36771
rect 12449 36737 12483 36771
rect 12483 36737 12492 36771
rect 12440 36728 12492 36737
rect 14648 36771 14700 36780
rect 14648 36737 14657 36771
rect 14657 36737 14691 36771
rect 14691 36737 14700 36771
rect 14648 36728 14700 36737
rect 13728 36660 13780 36712
rect 14372 36703 14424 36712
rect 14372 36669 14381 36703
rect 14381 36669 14415 36703
rect 14415 36669 14424 36703
rect 14372 36660 14424 36669
rect 11704 36524 11756 36576
rect 13084 36524 13136 36576
rect 16396 36728 16448 36780
rect 17132 36703 17184 36712
rect 17132 36669 17141 36703
rect 17141 36669 17175 36703
rect 17175 36669 17184 36703
rect 17132 36660 17184 36669
rect 17684 36660 17736 36712
rect 18788 36728 18840 36780
rect 19524 36796 19576 36848
rect 22008 36864 22060 36916
rect 21824 36796 21876 36848
rect 19892 36660 19944 36712
rect 20536 36703 20588 36712
rect 20536 36669 20545 36703
rect 20545 36669 20579 36703
rect 20579 36669 20588 36703
rect 20536 36660 20588 36669
rect 20812 36703 20864 36712
rect 20812 36669 20821 36703
rect 20821 36669 20855 36703
rect 20855 36669 20864 36703
rect 20812 36660 20864 36669
rect 20996 36703 21048 36712
rect 20996 36669 21005 36703
rect 21005 36669 21039 36703
rect 21039 36669 21048 36703
rect 20996 36660 21048 36669
rect 15200 36524 15252 36576
rect 17500 36524 17552 36576
rect 20076 36524 20128 36576
rect 21272 36728 21324 36780
rect 22284 36728 22336 36780
rect 23848 36864 23900 36916
rect 25412 36864 25464 36916
rect 24400 36796 24452 36848
rect 25872 36864 25924 36916
rect 26516 36864 26568 36916
rect 21456 36635 21508 36644
rect 21456 36601 21465 36635
rect 21465 36601 21499 36635
rect 21499 36601 21508 36635
rect 21456 36592 21508 36601
rect 21364 36524 21416 36576
rect 25964 36728 26016 36780
rect 32956 36907 33008 36916
rect 32956 36873 32965 36907
rect 32965 36873 32999 36907
rect 32999 36873 33008 36907
rect 32956 36864 33008 36873
rect 34796 36864 34848 36916
rect 27712 36839 27764 36848
rect 27712 36805 27721 36839
rect 27721 36805 27755 36839
rect 27755 36805 27764 36839
rect 27712 36796 27764 36805
rect 29000 36796 29052 36848
rect 30564 36796 30616 36848
rect 26516 36771 26568 36780
rect 26516 36737 26525 36771
rect 26525 36737 26559 36771
rect 26559 36737 26568 36771
rect 26516 36728 26568 36737
rect 26608 36771 26660 36780
rect 26608 36737 26622 36771
rect 26622 36737 26656 36771
rect 26656 36737 26660 36771
rect 26608 36728 26660 36737
rect 27068 36771 27120 36780
rect 27068 36737 27077 36771
rect 27077 36737 27111 36771
rect 27111 36737 27120 36771
rect 27068 36728 27120 36737
rect 27344 36728 27396 36780
rect 24124 36703 24176 36712
rect 24124 36669 24133 36703
rect 24133 36669 24167 36703
rect 24167 36669 24176 36703
rect 24124 36660 24176 36669
rect 25504 36703 25556 36712
rect 25504 36669 25513 36703
rect 25513 36669 25547 36703
rect 25547 36669 25556 36703
rect 25504 36660 25556 36669
rect 24676 36592 24728 36644
rect 24860 36592 24912 36644
rect 26148 36592 26200 36644
rect 27252 36635 27304 36644
rect 27252 36601 27261 36635
rect 27261 36601 27295 36635
rect 27295 36601 27304 36635
rect 27252 36592 27304 36601
rect 27344 36592 27396 36644
rect 29552 36703 29604 36712
rect 29552 36669 29561 36703
rect 29561 36669 29595 36703
rect 29595 36669 29604 36703
rect 29552 36660 29604 36669
rect 29736 36771 29788 36780
rect 29736 36737 29745 36771
rect 29745 36737 29779 36771
rect 29779 36737 29788 36771
rect 29736 36728 29788 36737
rect 30380 36771 30432 36780
rect 30380 36737 30389 36771
rect 30389 36737 30423 36771
rect 30423 36737 30432 36771
rect 31024 36771 31076 36780
rect 30380 36728 30432 36737
rect 31024 36737 31033 36771
rect 31033 36737 31067 36771
rect 31067 36737 31076 36771
rect 31024 36728 31076 36737
rect 31116 36728 31168 36780
rect 32312 36839 32364 36848
rect 32312 36805 32353 36839
rect 32353 36805 32364 36839
rect 32312 36796 32364 36805
rect 33416 36796 33468 36848
rect 33968 36796 34020 36848
rect 31668 36660 31720 36712
rect 32036 36728 32088 36780
rect 32128 36660 32180 36712
rect 33140 36728 33192 36780
rect 33232 36771 33284 36780
rect 33232 36737 33241 36771
rect 33241 36737 33275 36771
rect 33275 36737 33284 36771
rect 33232 36728 33284 36737
rect 33508 36703 33560 36712
rect 33508 36669 33517 36703
rect 33517 36669 33551 36703
rect 33551 36669 33560 36703
rect 33508 36660 33560 36669
rect 25228 36567 25280 36576
rect 25228 36533 25237 36567
rect 25237 36533 25271 36567
rect 25271 36533 25280 36567
rect 25228 36524 25280 36533
rect 27436 36524 27488 36576
rect 30104 36524 30156 36576
rect 31300 36524 31352 36576
rect 32404 36524 32456 36576
rect 32864 36524 32916 36576
rect 33324 36524 33376 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 12440 36320 12492 36372
rect 12992 36320 13044 36372
rect 14372 36320 14424 36372
rect 18512 36320 18564 36372
rect 18788 36320 18840 36372
rect 20996 36320 21048 36372
rect 21824 36320 21876 36372
rect 25504 36320 25556 36372
rect 25964 36320 26016 36372
rect 26516 36320 26568 36372
rect 24952 36252 25004 36304
rect 11704 36227 11756 36236
rect 11704 36193 11713 36227
rect 11713 36193 11747 36227
rect 11747 36193 11756 36227
rect 11704 36184 11756 36193
rect 13728 36184 13780 36236
rect 16396 36184 16448 36236
rect 16488 36184 16540 36236
rect 17500 36227 17552 36236
rect 17500 36193 17509 36227
rect 17509 36193 17543 36227
rect 17543 36193 17552 36227
rect 17500 36184 17552 36193
rect 20904 36184 20956 36236
rect 25412 36184 25464 36236
rect 26148 36184 26200 36236
rect 27620 36184 27672 36236
rect 13084 36116 13136 36168
rect 15476 36116 15528 36168
rect 19984 36159 20036 36168
rect 19984 36125 19993 36159
rect 19993 36125 20027 36159
rect 20027 36125 20036 36159
rect 19984 36116 20036 36125
rect 25780 36116 25832 36168
rect 12348 36048 12400 36100
rect 11520 35980 11572 36032
rect 18144 35980 18196 36032
rect 19524 36048 19576 36100
rect 20536 36048 20588 36100
rect 21272 36048 21324 36100
rect 24768 36048 24820 36100
rect 24676 35980 24728 36032
rect 25964 36159 26016 36168
rect 25964 36125 25973 36159
rect 25973 36125 26007 36159
rect 26007 36125 26016 36159
rect 25964 36116 26016 36125
rect 29184 36320 29236 36372
rect 29552 36320 29604 36372
rect 29920 36320 29972 36372
rect 30932 36320 30984 36372
rect 31024 36320 31076 36372
rect 28724 36252 28776 36304
rect 28724 36116 28776 36168
rect 29552 36184 29604 36236
rect 30104 36227 30156 36236
rect 30104 36193 30113 36227
rect 30113 36193 30147 36227
rect 30147 36193 30156 36227
rect 30104 36184 30156 36193
rect 30472 36184 30524 36236
rect 29368 36116 29420 36168
rect 25504 36023 25556 36032
rect 25504 35989 25513 36023
rect 25513 35989 25547 36023
rect 25547 35989 25556 36023
rect 25504 35980 25556 35989
rect 28816 36048 28868 36100
rect 31116 36184 31168 36236
rect 28908 35980 28960 36032
rect 29000 35980 29052 36032
rect 30932 36159 30984 36168
rect 30932 36125 30941 36159
rect 30941 36125 30975 36159
rect 30975 36125 30984 36159
rect 30932 36116 30984 36125
rect 31392 36091 31444 36100
rect 31392 36057 31401 36091
rect 31401 36057 31435 36091
rect 31435 36057 31444 36091
rect 31392 36048 31444 36057
rect 32036 36320 32088 36372
rect 33508 36363 33560 36372
rect 33508 36329 33517 36363
rect 33517 36329 33551 36363
rect 33551 36329 33560 36363
rect 33508 36320 33560 36329
rect 31852 36252 31904 36304
rect 32128 36184 32180 36236
rect 32312 36184 32364 36236
rect 34796 36252 34848 36304
rect 31852 36048 31904 36100
rect 33140 36116 33192 36168
rect 33324 36159 33376 36168
rect 33324 36125 33333 36159
rect 33333 36125 33367 36159
rect 33367 36125 33376 36159
rect 33324 36116 33376 36125
rect 33600 36159 33652 36168
rect 33600 36125 33609 36159
rect 33609 36125 33643 36159
rect 33643 36125 33652 36159
rect 33600 36116 33652 36125
rect 34796 36116 34848 36168
rect 32404 36048 32456 36100
rect 32220 36023 32272 36032
rect 32220 35989 32229 36023
rect 32229 35989 32263 36023
rect 32263 35989 32272 36023
rect 32220 35980 32272 35989
rect 32772 36023 32824 36032
rect 32772 35989 32781 36023
rect 32781 35989 32815 36023
rect 32815 35989 32824 36023
rect 32772 35980 32824 35989
rect 32864 35980 32916 36032
rect 34612 35980 34664 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 12992 35819 13044 35828
rect 12992 35785 13001 35819
rect 13001 35785 13035 35819
rect 13035 35785 13044 35819
rect 12992 35776 13044 35785
rect 18512 35776 18564 35828
rect 20904 35819 20956 35828
rect 20904 35785 20913 35819
rect 20913 35785 20947 35819
rect 20947 35785 20956 35819
rect 20904 35776 20956 35785
rect 20996 35776 21048 35828
rect 21364 35819 21416 35828
rect 21364 35785 21373 35819
rect 21373 35785 21407 35819
rect 21407 35785 21416 35819
rect 21364 35776 21416 35785
rect 24124 35776 24176 35828
rect 16948 35708 17000 35760
rect 20812 35708 20864 35760
rect 22284 35708 22336 35760
rect 11888 35640 11940 35692
rect 19064 35640 19116 35692
rect 13728 35572 13780 35624
rect 16212 35615 16264 35624
rect 16212 35581 16221 35615
rect 16221 35581 16255 35615
rect 16255 35581 16264 35615
rect 16212 35572 16264 35581
rect 16396 35615 16448 35624
rect 16396 35581 16405 35615
rect 16405 35581 16439 35615
rect 16439 35581 16448 35615
rect 16396 35572 16448 35581
rect 18880 35615 18932 35624
rect 18880 35581 18889 35615
rect 18889 35581 18923 35615
rect 18923 35581 18932 35615
rect 18880 35572 18932 35581
rect 20260 35572 20312 35624
rect 23572 35683 23624 35692
rect 23572 35649 23581 35683
rect 23581 35649 23615 35683
rect 23615 35649 23624 35683
rect 23572 35640 23624 35649
rect 21456 35615 21508 35624
rect 21456 35581 21465 35615
rect 21465 35581 21499 35615
rect 21499 35581 21508 35615
rect 21456 35572 21508 35581
rect 25228 35708 25280 35760
rect 27620 35708 27672 35760
rect 27712 35640 27764 35692
rect 27988 35683 28040 35692
rect 27988 35649 27997 35683
rect 27997 35649 28031 35683
rect 28031 35649 28040 35683
rect 27988 35640 28040 35649
rect 25136 35572 25188 35624
rect 25412 35615 25464 35624
rect 25412 35581 25421 35615
rect 25421 35581 25455 35615
rect 25455 35581 25464 35615
rect 25412 35572 25464 35581
rect 26240 35572 26292 35624
rect 27252 35572 27304 35624
rect 31760 35776 31812 35828
rect 33140 35776 33192 35828
rect 34244 35776 34296 35828
rect 30564 35708 30616 35760
rect 31392 35708 31444 35760
rect 28540 35640 28592 35692
rect 27068 35547 27120 35556
rect 27068 35513 27077 35547
rect 27077 35513 27111 35547
rect 27111 35513 27120 35547
rect 27068 35504 27120 35513
rect 13360 35436 13412 35488
rect 15476 35436 15528 35488
rect 17592 35436 17644 35488
rect 27436 35436 27488 35488
rect 27712 35436 27764 35488
rect 29368 35436 29420 35488
rect 29736 35683 29788 35692
rect 29736 35649 29745 35683
rect 29745 35649 29779 35683
rect 29779 35649 29788 35683
rect 29736 35640 29788 35649
rect 29828 35683 29880 35692
rect 29828 35649 29837 35683
rect 29837 35649 29871 35683
rect 29871 35649 29880 35683
rect 29828 35640 29880 35649
rect 31576 35640 31628 35692
rect 31760 35640 31812 35692
rect 31852 35504 31904 35556
rect 32220 35640 32272 35692
rect 32312 35572 32364 35624
rect 33232 35708 33284 35760
rect 33324 35683 33376 35692
rect 33324 35649 33333 35683
rect 33333 35649 33367 35683
rect 33367 35649 33376 35683
rect 33324 35640 33376 35649
rect 32036 35504 32088 35556
rect 32772 35547 32824 35556
rect 32772 35513 32781 35547
rect 32781 35513 32815 35547
rect 32815 35513 32824 35547
rect 32772 35504 32824 35513
rect 31576 35479 31628 35488
rect 31576 35445 31585 35479
rect 31585 35445 31619 35479
rect 31619 35445 31628 35479
rect 31576 35436 31628 35445
rect 33048 35436 33100 35488
rect 33600 35683 33652 35692
rect 33600 35649 33609 35683
rect 33609 35649 33643 35683
rect 33643 35649 33652 35683
rect 33600 35640 33652 35649
rect 33968 35708 34020 35760
rect 34060 35708 34112 35760
rect 34428 35708 34480 35760
rect 34152 35436 34204 35488
rect 35624 35436 35676 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 11888 35275 11940 35284
rect 11888 35241 11897 35275
rect 11897 35241 11931 35275
rect 11931 35241 11940 35275
rect 11888 35232 11940 35241
rect 16948 35275 17000 35284
rect 16948 35241 16957 35275
rect 16957 35241 16991 35275
rect 16991 35241 17000 35275
rect 16948 35232 17000 35241
rect 19064 35275 19116 35284
rect 19064 35241 19073 35275
rect 19073 35241 19107 35275
rect 19107 35241 19116 35275
rect 19064 35232 19116 35241
rect 11520 35096 11572 35148
rect 14188 35096 14240 35148
rect 15200 35139 15252 35148
rect 15200 35105 15209 35139
rect 15209 35105 15243 35139
rect 15243 35105 15252 35139
rect 15200 35096 15252 35105
rect 17592 35139 17644 35148
rect 17592 35105 17601 35139
rect 17601 35105 17635 35139
rect 17635 35105 17644 35139
rect 17592 35096 17644 35105
rect 18144 35096 18196 35148
rect 12348 34960 12400 35012
rect 13360 35003 13412 35012
rect 13360 34969 13369 35003
rect 13369 34969 13403 35003
rect 13403 34969 13412 35003
rect 13360 34960 13412 34969
rect 15476 35003 15528 35012
rect 15476 34969 15485 35003
rect 15485 34969 15519 35003
rect 15519 34969 15528 35003
rect 15476 34960 15528 34969
rect 15568 34960 15620 35012
rect 19800 35139 19852 35148
rect 19800 35105 19809 35139
rect 19809 35105 19843 35139
rect 19843 35105 19852 35139
rect 19800 35096 19852 35105
rect 18880 35028 18932 35080
rect 16396 34892 16448 34944
rect 19524 34960 19576 35012
rect 19156 34892 19208 34944
rect 20536 34892 20588 34944
rect 25964 35232 26016 35284
rect 26240 35275 26292 35284
rect 26240 35241 26249 35275
rect 26249 35241 26283 35275
rect 26283 35241 26292 35275
rect 26240 35232 26292 35241
rect 25412 35096 25464 35148
rect 29736 35232 29788 35284
rect 33600 35232 33652 35284
rect 28632 35164 28684 35216
rect 24400 35071 24452 35080
rect 24400 35037 24409 35071
rect 24409 35037 24443 35071
rect 24443 35037 24452 35071
rect 24400 35028 24452 35037
rect 24952 34960 25004 35012
rect 25136 34960 25188 35012
rect 25964 34960 26016 35012
rect 28448 35028 28500 35080
rect 28724 35071 28776 35080
rect 28724 35037 28733 35071
rect 28733 35037 28767 35071
rect 28767 35037 28776 35071
rect 28724 35028 28776 35037
rect 28816 35071 28868 35080
rect 28816 35037 28825 35071
rect 28825 35037 28859 35071
rect 28859 35037 28868 35071
rect 28816 35028 28868 35037
rect 29184 35028 29236 35080
rect 30472 35028 30524 35080
rect 31392 35164 31444 35216
rect 31760 35139 31812 35148
rect 31760 35105 31769 35139
rect 31769 35105 31803 35139
rect 31803 35105 31812 35139
rect 31760 35096 31812 35105
rect 31944 35139 31996 35148
rect 31944 35105 31953 35139
rect 31953 35105 31987 35139
rect 31987 35105 31996 35139
rect 31944 35096 31996 35105
rect 32036 35096 32088 35148
rect 29092 34960 29144 35012
rect 28172 34892 28224 34944
rect 30012 34892 30064 34944
rect 30104 34935 30156 34944
rect 30104 34901 30113 34935
rect 30113 34901 30147 34935
rect 30147 34901 30156 34935
rect 30104 34892 30156 34901
rect 30656 34935 30708 34944
rect 30656 34901 30665 34935
rect 30665 34901 30699 34935
rect 30699 34901 30708 34935
rect 30656 34892 30708 34901
rect 31852 35071 31904 35080
rect 31852 35037 31861 35071
rect 31861 35037 31895 35071
rect 31895 35037 31904 35071
rect 31852 35028 31904 35037
rect 32128 35028 32180 35080
rect 32036 34960 32088 35012
rect 32680 35096 32732 35148
rect 33324 35164 33376 35216
rect 33508 35139 33560 35148
rect 33508 35105 33517 35139
rect 33517 35105 33551 35139
rect 33551 35105 33560 35139
rect 33508 35096 33560 35105
rect 33876 35139 33928 35148
rect 33876 35105 33885 35139
rect 33885 35105 33919 35139
rect 33919 35105 33928 35139
rect 33876 35096 33928 35105
rect 33232 35028 33284 35080
rect 33324 35071 33376 35080
rect 33324 35037 33333 35071
rect 33333 35037 33367 35071
rect 33367 35037 33376 35071
rect 33324 35028 33376 35037
rect 33600 35071 33652 35080
rect 33600 35037 33609 35071
rect 33609 35037 33643 35071
rect 33643 35037 33652 35071
rect 33600 35028 33652 35037
rect 33048 34960 33100 35012
rect 34796 35071 34848 35080
rect 34796 35037 34805 35071
rect 34805 35037 34839 35071
rect 34839 35037 34848 35071
rect 34796 35028 34848 35037
rect 35532 35071 35584 35080
rect 35532 35037 35541 35071
rect 35541 35037 35575 35071
rect 35575 35037 35584 35071
rect 35532 35028 35584 35037
rect 35624 35071 35676 35080
rect 35624 35037 35633 35071
rect 35633 35037 35667 35071
rect 35667 35037 35676 35071
rect 35624 35028 35676 35037
rect 31852 34892 31904 34944
rect 33600 34892 33652 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 11888 34688 11940 34740
rect 16212 34688 16264 34740
rect 13544 34620 13596 34672
rect 13084 34595 13136 34604
rect 13084 34561 13093 34595
rect 13093 34561 13127 34595
rect 13127 34561 13136 34595
rect 13084 34552 13136 34561
rect 14188 34595 14240 34604
rect 14188 34561 14197 34595
rect 14197 34561 14231 34595
rect 14231 34561 14240 34595
rect 14188 34552 14240 34561
rect 15568 34552 15620 34604
rect 13360 34527 13412 34536
rect 13360 34493 13369 34527
rect 13369 34493 13403 34527
rect 13403 34493 13412 34527
rect 13360 34484 13412 34493
rect 13820 34416 13872 34468
rect 18880 34688 18932 34740
rect 19800 34688 19852 34740
rect 19340 34620 19392 34672
rect 19524 34620 19576 34672
rect 20536 34731 20588 34740
rect 20536 34697 20545 34731
rect 20545 34697 20579 34731
rect 20579 34697 20588 34731
rect 20536 34688 20588 34697
rect 25504 34688 25556 34740
rect 24676 34620 24728 34672
rect 25228 34620 25280 34672
rect 25964 34620 26016 34672
rect 27620 34620 27672 34672
rect 27804 34620 27856 34672
rect 28448 34731 28500 34740
rect 28448 34697 28457 34731
rect 28457 34697 28491 34731
rect 28491 34697 28500 34731
rect 28448 34688 28500 34697
rect 30656 34688 30708 34740
rect 31852 34688 31904 34740
rect 32220 34688 32272 34740
rect 33232 34688 33284 34740
rect 33416 34688 33468 34740
rect 34612 34688 34664 34740
rect 29460 34620 29512 34672
rect 31668 34620 31720 34672
rect 33048 34663 33100 34672
rect 20628 34595 20680 34604
rect 20628 34561 20637 34595
rect 20637 34561 20671 34595
rect 20671 34561 20680 34595
rect 20628 34552 20680 34561
rect 23480 34552 23532 34604
rect 26148 34552 26200 34604
rect 28908 34552 28960 34604
rect 29368 34595 29420 34604
rect 29368 34561 29377 34595
rect 29377 34561 29411 34595
rect 29411 34561 29420 34595
rect 29368 34552 29420 34561
rect 17776 34484 17828 34536
rect 19156 34484 19208 34536
rect 22560 34527 22612 34536
rect 22560 34493 22569 34527
rect 22569 34493 22603 34527
rect 22603 34493 22612 34527
rect 22560 34484 22612 34493
rect 12072 34348 12124 34400
rect 12716 34391 12768 34400
rect 12716 34357 12725 34391
rect 12725 34357 12759 34391
rect 12759 34357 12768 34391
rect 12716 34348 12768 34357
rect 24860 34416 24912 34468
rect 28172 34527 28224 34536
rect 28172 34493 28181 34527
rect 28181 34493 28215 34527
rect 28215 34493 28224 34527
rect 28172 34484 28224 34493
rect 28264 34527 28316 34536
rect 28264 34493 28273 34527
rect 28273 34493 28307 34527
rect 28307 34493 28316 34527
rect 28264 34484 28316 34493
rect 25780 34416 25832 34468
rect 29000 34484 29052 34536
rect 29092 34527 29144 34536
rect 29092 34493 29101 34527
rect 29101 34493 29135 34527
rect 29135 34493 29144 34527
rect 29092 34484 29144 34493
rect 29276 34484 29328 34536
rect 30104 34552 30156 34604
rect 30472 34595 30524 34604
rect 30472 34561 30481 34595
rect 30481 34561 30515 34595
rect 30515 34561 30524 34595
rect 30472 34552 30524 34561
rect 30932 34595 30984 34604
rect 30932 34561 30941 34595
rect 30941 34561 30975 34595
rect 30975 34561 30984 34595
rect 30932 34552 30984 34561
rect 31576 34595 31628 34604
rect 31576 34561 31585 34595
rect 31585 34561 31619 34595
rect 31619 34561 31628 34595
rect 31576 34552 31628 34561
rect 31944 34595 31996 34604
rect 31944 34561 31953 34595
rect 31953 34561 31987 34595
rect 31987 34561 31996 34595
rect 31944 34552 31996 34561
rect 32220 34552 32272 34604
rect 32496 34552 32548 34604
rect 33048 34629 33057 34663
rect 33057 34629 33091 34663
rect 33091 34629 33100 34663
rect 33048 34620 33100 34629
rect 34520 34620 34572 34672
rect 33232 34595 33284 34604
rect 33232 34561 33241 34595
rect 33241 34561 33275 34595
rect 33275 34561 33284 34595
rect 33232 34552 33284 34561
rect 33416 34595 33468 34604
rect 33416 34561 33425 34595
rect 33425 34561 33459 34595
rect 33459 34561 33468 34595
rect 33416 34552 33468 34561
rect 33692 34595 33744 34604
rect 33692 34561 33701 34595
rect 33701 34561 33735 34595
rect 33735 34561 33744 34595
rect 33692 34552 33744 34561
rect 33968 34595 34020 34604
rect 33968 34561 33977 34595
rect 33977 34561 34011 34595
rect 34011 34561 34020 34595
rect 33968 34552 34020 34561
rect 29736 34484 29788 34536
rect 30012 34484 30064 34536
rect 30564 34484 30616 34536
rect 32036 34484 32088 34536
rect 34336 34484 34388 34536
rect 33232 34416 33284 34468
rect 19616 34348 19668 34400
rect 21456 34348 21508 34400
rect 22100 34391 22152 34400
rect 22100 34357 22109 34391
rect 22109 34357 22143 34391
rect 22143 34357 22152 34391
rect 22100 34348 22152 34357
rect 25044 34391 25096 34400
rect 25044 34357 25053 34391
rect 25053 34357 25087 34391
rect 25087 34357 25096 34391
rect 25044 34348 25096 34357
rect 30288 34348 30340 34400
rect 30472 34348 30524 34400
rect 33048 34348 33100 34400
rect 34060 34348 34112 34400
rect 34336 34348 34388 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 13544 34187 13596 34196
rect 13544 34153 13553 34187
rect 13553 34153 13587 34187
rect 13587 34153 13596 34187
rect 13544 34144 13596 34153
rect 14280 34144 14332 34196
rect 23480 34144 23532 34196
rect 28172 34144 28224 34196
rect 30012 34144 30064 34196
rect 29368 34076 29420 34128
rect 11520 34008 11572 34060
rect 12072 34051 12124 34060
rect 12072 34017 12081 34051
rect 12081 34017 12115 34051
rect 12115 34017 12124 34051
rect 12072 34008 12124 34017
rect 14188 34008 14240 34060
rect 15568 34008 15620 34060
rect 18880 33940 18932 33992
rect 12348 33804 12400 33856
rect 15384 33872 15436 33924
rect 15568 33915 15620 33924
rect 15568 33881 15577 33915
rect 15577 33881 15611 33915
rect 15611 33881 15620 33915
rect 15568 33872 15620 33881
rect 15936 33915 15988 33924
rect 15936 33881 15945 33915
rect 15945 33881 15979 33915
rect 15979 33881 15988 33915
rect 15936 33872 15988 33881
rect 16396 33872 16448 33924
rect 17776 33872 17828 33924
rect 19340 34051 19392 34060
rect 19340 34017 19349 34051
rect 19349 34017 19383 34051
rect 19383 34017 19392 34051
rect 19340 34008 19392 34017
rect 19984 34008 20036 34060
rect 20628 34008 20680 34060
rect 25044 34008 25096 34060
rect 25136 34008 25188 34060
rect 28540 34008 28592 34060
rect 29184 34008 29236 34060
rect 21548 33983 21600 33992
rect 21548 33949 21557 33983
rect 21557 33949 21591 33983
rect 21591 33949 21600 33983
rect 21548 33940 21600 33949
rect 24400 33983 24452 33992
rect 24400 33949 24409 33983
rect 24409 33949 24443 33983
rect 24443 33949 24452 33983
rect 24400 33940 24452 33949
rect 29276 33983 29328 33992
rect 29276 33949 29285 33983
rect 29285 33949 29319 33983
rect 29319 33949 29328 33983
rect 29276 33940 29328 33949
rect 29368 33983 29420 33992
rect 29368 33949 29377 33983
rect 29377 33949 29411 33983
rect 29411 33949 29420 33983
rect 29368 33940 29420 33949
rect 31944 34144 31996 34196
rect 33416 34144 33468 34196
rect 31484 34051 31536 34060
rect 31484 34017 31493 34051
rect 31493 34017 31527 34051
rect 31527 34017 31536 34051
rect 31484 34008 31536 34017
rect 32772 34008 32824 34060
rect 31300 33940 31352 33992
rect 34612 34008 34664 34060
rect 34336 33983 34388 33992
rect 34336 33949 34345 33983
rect 34345 33949 34379 33983
rect 34379 33949 34388 33983
rect 34336 33940 34388 33949
rect 35716 33983 35768 33992
rect 35716 33949 35725 33983
rect 35725 33949 35759 33983
rect 35759 33949 35768 33983
rect 35716 33940 35768 33949
rect 19524 33872 19576 33924
rect 19708 33872 19760 33924
rect 21272 33872 21324 33924
rect 22100 33872 22152 33924
rect 17408 33847 17460 33856
rect 17408 33813 17417 33847
rect 17417 33813 17451 33847
rect 17451 33813 17460 33847
rect 17408 33804 17460 33813
rect 20628 33804 20680 33856
rect 25228 33872 25280 33924
rect 25964 33872 26016 33924
rect 22192 33804 22244 33856
rect 25504 33804 25556 33856
rect 29644 33872 29696 33924
rect 30380 33804 30432 33856
rect 30656 33804 30708 33856
rect 34520 33872 34572 33924
rect 35256 33872 35308 33924
rect 34428 33804 34480 33856
rect 34612 33804 34664 33856
rect 35440 33847 35492 33856
rect 35440 33813 35449 33847
rect 35449 33813 35483 33847
rect 35483 33813 35492 33847
rect 35440 33804 35492 33813
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 12716 33600 12768 33652
rect 13084 33600 13136 33652
rect 12348 33532 12400 33584
rect 14280 33575 14332 33584
rect 14280 33541 14289 33575
rect 14289 33541 14323 33575
rect 14323 33541 14332 33575
rect 14280 33532 14332 33541
rect 15936 33600 15988 33652
rect 17408 33600 17460 33652
rect 17684 33600 17736 33652
rect 19616 33600 19668 33652
rect 19708 33643 19760 33652
rect 19708 33609 19717 33643
rect 19717 33609 19751 33643
rect 19751 33609 19760 33643
rect 19708 33600 19760 33609
rect 20444 33600 20496 33652
rect 22560 33600 22612 33652
rect 17776 33532 17828 33584
rect 19524 33532 19576 33584
rect 20352 33532 20404 33584
rect 21548 33532 21600 33584
rect 25228 33600 25280 33652
rect 26148 33600 26200 33652
rect 11520 33507 11572 33516
rect 11520 33473 11529 33507
rect 11529 33473 11563 33507
rect 11563 33473 11572 33507
rect 11520 33464 11572 33473
rect 15384 33464 15436 33516
rect 16396 33464 16448 33516
rect 17040 33464 17092 33516
rect 19708 33464 19760 33516
rect 20628 33464 20680 33516
rect 21456 33464 21508 33516
rect 13912 33396 13964 33448
rect 17684 33439 17736 33448
rect 17684 33405 17693 33439
rect 17693 33405 17727 33439
rect 17727 33405 17736 33439
rect 17684 33396 17736 33405
rect 18052 33396 18104 33448
rect 20260 33439 20312 33448
rect 20260 33405 20269 33439
rect 20269 33405 20303 33439
rect 20303 33405 20312 33439
rect 20260 33396 20312 33405
rect 22284 33439 22336 33448
rect 22284 33405 22293 33439
rect 22293 33405 22327 33439
rect 22327 33405 22336 33439
rect 22284 33396 22336 33405
rect 24400 33464 24452 33516
rect 25136 33532 25188 33584
rect 27712 33464 27764 33516
rect 30380 33532 30432 33584
rect 30656 33532 30708 33584
rect 33048 33600 33100 33652
rect 32772 33532 32824 33584
rect 33692 33600 33744 33652
rect 34428 33643 34480 33652
rect 34428 33609 34437 33643
rect 34437 33609 34471 33643
rect 34471 33609 34480 33643
rect 34428 33600 34480 33609
rect 34704 33600 34756 33652
rect 22928 33439 22980 33448
rect 22928 33405 22937 33439
rect 22937 33405 22971 33439
rect 22971 33405 22980 33439
rect 22928 33396 22980 33405
rect 24860 33439 24912 33448
rect 24860 33405 24869 33439
rect 24869 33405 24903 33439
rect 24903 33405 24912 33439
rect 24860 33396 24912 33405
rect 26056 33396 26108 33448
rect 19800 33328 19852 33380
rect 18512 33260 18564 33312
rect 21088 33260 21140 33312
rect 24400 33303 24452 33312
rect 24400 33269 24409 33303
rect 24409 33269 24443 33303
rect 24443 33269 24452 33303
rect 24400 33260 24452 33269
rect 28080 33303 28132 33312
rect 28080 33269 28089 33303
rect 28089 33269 28123 33303
rect 28123 33269 28132 33303
rect 28080 33260 28132 33269
rect 29368 33507 29420 33516
rect 29368 33473 29377 33507
rect 29377 33473 29411 33507
rect 29411 33473 29420 33507
rect 29368 33464 29420 33473
rect 29460 33464 29512 33516
rect 29644 33507 29696 33516
rect 29644 33473 29653 33507
rect 29653 33473 29687 33507
rect 29687 33473 29696 33507
rect 29644 33464 29696 33473
rect 29828 33507 29880 33516
rect 29828 33473 29837 33507
rect 29837 33473 29871 33507
rect 29871 33473 29880 33507
rect 29828 33464 29880 33473
rect 31392 33464 31444 33516
rect 33508 33464 33560 33516
rect 34704 33464 34756 33516
rect 29092 33396 29144 33448
rect 31576 33439 31628 33448
rect 31576 33405 31585 33439
rect 31585 33405 31619 33439
rect 31619 33405 31628 33439
rect 31576 33396 31628 33405
rect 33600 33396 33652 33448
rect 34060 33439 34112 33448
rect 34060 33405 34069 33439
rect 34069 33405 34103 33439
rect 34103 33405 34112 33439
rect 34060 33396 34112 33405
rect 34152 33439 34204 33448
rect 34152 33405 34161 33439
rect 34161 33405 34195 33439
rect 34195 33405 34204 33439
rect 34152 33396 34204 33405
rect 34796 33396 34848 33448
rect 35256 33439 35308 33448
rect 35256 33405 35265 33439
rect 35265 33405 35299 33439
rect 35299 33405 35308 33439
rect 35256 33396 35308 33405
rect 34520 33328 34572 33380
rect 29000 33260 29052 33312
rect 32404 33260 32456 33312
rect 34612 33303 34664 33312
rect 34612 33269 34621 33303
rect 34621 33269 34655 33303
rect 34655 33269 34664 33303
rect 34612 33260 34664 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 17040 33099 17092 33108
rect 17040 33065 17049 33099
rect 17049 33065 17083 33099
rect 17083 33065 17092 33099
rect 17040 33056 17092 33065
rect 22560 33099 22612 33108
rect 22560 33065 22569 33099
rect 22569 33065 22603 33099
rect 22603 33065 22612 33099
rect 22560 33056 22612 33065
rect 22928 33056 22980 33108
rect 24860 33056 24912 33108
rect 28540 33099 28592 33108
rect 28540 33065 28549 33099
rect 28549 33065 28583 33099
rect 28583 33065 28592 33099
rect 28540 33056 28592 33065
rect 19616 32988 19668 33040
rect 13084 32920 13136 32972
rect 13360 32963 13412 32972
rect 13360 32929 13369 32963
rect 13369 32929 13403 32963
rect 13403 32929 13412 32963
rect 13360 32920 13412 32929
rect 18512 32963 18564 32972
rect 18512 32929 18521 32963
rect 18521 32929 18555 32963
rect 18555 32929 18564 32963
rect 18512 32920 18564 32929
rect 19708 32963 19760 32972
rect 19708 32929 19717 32963
rect 19717 32929 19751 32963
rect 19751 32929 19760 32963
rect 19708 32920 19760 32929
rect 21088 32963 21140 32972
rect 21088 32929 21097 32963
rect 21097 32929 21131 32963
rect 21131 32929 21140 32963
rect 21088 32920 21140 32929
rect 24676 32988 24728 33040
rect 25780 32963 25832 32972
rect 25780 32929 25789 32963
rect 25789 32929 25823 32963
rect 25823 32929 25832 32963
rect 25780 32920 25832 32929
rect 27804 32988 27856 33040
rect 28816 33056 28868 33108
rect 30104 33099 30156 33108
rect 30104 33065 30113 33099
rect 30113 33065 30147 33099
rect 30147 33065 30156 33099
rect 30104 33056 30156 33065
rect 30288 33099 30340 33108
rect 30288 33065 30297 33099
rect 30297 33065 30331 33099
rect 30331 33065 30340 33099
rect 30288 33056 30340 33065
rect 34704 33056 34756 33108
rect 29644 32988 29696 33040
rect 29000 32963 29052 32972
rect 29000 32929 29009 32963
rect 29009 32929 29043 32963
rect 29043 32929 29052 32963
rect 29000 32920 29052 32929
rect 30012 32920 30064 32972
rect 31852 32988 31904 33040
rect 33600 32988 33652 33040
rect 31576 32920 31628 32972
rect 33324 32920 33376 32972
rect 34336 32920 34388 32972
rect 35256 32920 35308 32972
rect 13912 32852 13964 32904
rect 19064 32852 19116 32904
rect 22192 32852 22244 32904
rect 23572 32852 23624 32904
rect 24400 32852 24452 32904
rect 25136 32852 25188 32904
rect 26056 32895 26108 32904
rect 26056 32861 26065 32895
rect 26065 32861 26099 32895
rect 26099 32861 26108 32895
rect 26056 32852 26108 32861
rect 16396 32784 16448 32836
rect 18236 32784 18288 32836
rect 26148 32784 26200 32836
rect 29184 32895 29236 32904
rect 29184 32861 29193 32895
rect 29193 32861 29227 32895
rect 29227 32861 29236 32895
rect 29184 32852 29236 32861
rect 29736 32852 29788 32904
rect 30196 32895 30248 32904
rect 30196 32861 30205 32895
rect 30205 32861 30239 32895
rect 30239 32861 30248 32895
rect 30196 32852 30248 32861
rect 30932 32852 30984 32904
rect 31116 32895 31168 32904
rect 31116 32861 31125 32895
rect 31125 32861 31159 32895
rect 31159 32861 31168 32895
rect 31116 32852 31168 32861
rect 32404 32895 32456 32904
rect 32404 32861 32413 32895
rect 32413 32861 32447 32895
rect 32447 32861 32456 32895
rect 32404 32852 32456 32861
rect 28908 32827 28960 32836
rect 28908 32793 28917 32827
rect 28917 32793 28951 32827
rect 28951 32793 28960 32827
rect 28908 32784 28960 32793
rect 30380 32784 30432 32836
rect 31668 32784 31720 32836
rect 33232 32784 33284 32836
rect 35440 32852 35492 32904
rect 35164 32784 35216 32836
rect 12072 32716 12124 32768
rect 13084 32759 13136 32768
rect 13084 32725 13093 32759
rect 13093 32725 13127 32759
rect 13127 32725 13136 32759
rect 13084 32716 13136 32725
rect 19524 32716 19576 32768
rect 23480 32716 23532 32768
rect 25688 32759 25740 32768
rect 25688 32725 25697 32759
rect 25697 32725 25731 32759
rect 25731 32725 25740 32759
rect 25688 32716 25740 32725
rect 28816 32716 28868 32768
rect 30564 32716 30616 32768
rect 30748 32716 30800 32768
rect 35348 32716 35400 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 18052 32555 18104 32564
rect 18052 32521 18061 32555
rect 18061 32521 18095 32555
rect 18095 32521 18104 32555
rect 18052 32512 18104 32521
rect 22284 32512 22336 32564
rect 25780 32512 25832 32564
rect 15568 32444 15620 32496
rect 16396 32444 16448 32496
rect 19524 32487 19576 32496
rect 19524 32453 19533 32487
rect 19533 32453 19567 32487
rect 19567 32453 19576 32487
rect 19524 32444 19576 32453
rect 20352 32487 20404 32496
rect 20352 32453 20361 32487
rect 20361 32453 20395 32487
rect 20395 32453 20404 32487
rect 20352 32444 20404 32453
rect 24860 32444 24912 32496
rect 27712 32444 27764 32496
rect 27896 32444 27948 32496
rect 29000 32512 29052 32564
rect 29184 32444 29236 32496
rect 14280 32376 14332 32428
rect 17040 32419 17092 32428
rect 17040 32385 17049 32419
rect 17049 32385 17083 32419
rect 17083 32385 17092 32419
rect 17040 32376 17092 32385
rect 26056 32376 26108 32428
rect 11612 32308 11664 32360
rect 13176 32351 13228 32360
rect 13176 32317 13185 32351
rect 13185 32317 13219 32351
rect 13219 32317 13228 32351
rect 13176 32308 13228 32317
rect 15292 32308 15344 32360
rect 15936 32308 15988 32360
rect 17408 32308 17460 32360
rect 13912 32172 13964 32224
rect 14188 32172 14240 32224
rect 14832 32172 14884 32224
rect 15568 32172 15620 32224
rect 19064 32172 19116 32224
rect 22100 32308 22152 32360
rect 22468 32351 22520 32360
rect 22468 32317 22477 32351
rect 22477 32317 22511 32351
rect 22511 32317 22520 32351
rect 22468 32308 22520 32317
rect 28080 32308 28132 32360
rect 29920 32419 29972 32428
rect 29920 32385 29929 32419
rect 29929 32385 29963 32419
rect 29963 32385 29972 32419
rect 29920 32376 29972 32385
rect 31300 32512 31352 32564
rect 31392 32444 31444 32496
rect 32864 32512 32916 32564
rect 29828 32308 29880 32360
rect 30564 32308 30616 32360
rect 30748 32419 30800 32428
rect 30748 32385 30757 32419
rect 30757 32385 30791 32419
rect 30791 32385 30800 32419
rect 30748 32376 30800 32385
rect 31668 32376 31720 32428
rect 32588 32419 32640 32428
rect 32588 32385 32597 32419
rect 32597 32385 32631 32419
rect 32631 32385 32640 32419
rect 32588 32376 32640 32385
rect 33968 32444 34020 32496
rect 34428 32376 34480 32428
rect 32312 32240 32364 32292
rect 20996 32172 21048 32224
rect 29920 32215 29972 32224
rect 29920 32181 29929 32215
rect 29929 32181 29963 32215
rect 29963 32181 29972 32215
rect 29920 32172 29972 32181
rect 30104 32172 30156 32224
rect 30288 32172 30340 32224
rect 30380 32172 30432 32224
rect 34612 32308 34664 32360
rect 35164 32419 35216 32428
rect 35164 32385 35173 32419
rect 35173 32385 35207 32419
rect 35207 32385 35216 32419
rect 35164 32376 35216 32385
rect 35256 32376 35308 32428
rect 34520 32240 34572 32292
rect 34152 32172 34204 32224
rect 35348 32172 35400 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 13084 31968 13136 32020
rect 13544 32011 13596 32020
rect 13544 31977 13553 32011
rect 13553 31977 13587 32011
rect 13587 31977 13596 32011
rect 13544 31968 13596 31977
rect 17040 32011 17092 32020
rect 17040 31977 17049 32011
rect 17049 31977 17083 32011
rect 17083 31977 17092 32011
rect 17040 31968 17092 31977
rect 22284 31968 22336 32020
rect 26056 31968 26108 32020
rect 13820 31900 13872 31952
rect 12072 31875 12124 31884
rect 12072 31841 12081 31875
rect 12081 31841 12115 31875
rect 12115 31841 12124 31875
rect 12072 31832 12124 31841
rect 11612 31764 11664 31816
rect 14280 31832 14332 31884
rect 14832 31832 14884 31884
rect 15568 31875 15620 31884
rect 15568 31841 15577 31875
rect 15577 31841 15611 31875
rect 15611 31841 15620 31875
rect 15568 31832 15620 31841
rect 19064 31832 19116 31884
rect 20996 31875 21048 31884
rect 20996 31841 21005 31875
rect 21005 31841 21039 31875
rect 21039 31841 21048 31875
rect 20996 31832 21048 31841
rect 22192 31832 22244 31884
rect 23572 31875 23624 31884
rect 23572 31841 23581 31875
rect 23581 31841 23615 31875
rect 23615 31841 23624 31875
rect 23572 31832 23624 31841
rect 24768 31832 24820 31884
rect 25688 31832 25740 31884
rect 26976 31832 27028 31884
rect 27620 31968 27672 32020
rect 27988 31875 28040 31884
rect 27988 31841 27997 31875
rect 27997 31841 28031 31875
rect 28031 31841 28040 31875
rect 27988 31832 28040 31841
rect 14188 31764 14240 31816
rect 15292 31807 15344 31816
rect 15292 31773 15301 31807
rect 15301 31773 15335 31807
rect 15335 31773 15344 31807
rect 15292 31764 15344 31773
rect 25228 31764 25280 31816
rect 30288 31968 30340 32020
rect 32588 31968 32640 32020
rect 29920 31900 29972 31952
rect 34612 31900 34664 31952
rect 31392 31832 31444 31884
rect 29184 31807 29236 31816
rect 29184 31773 29193 31807
rect 29193 31773 29227 31807
rect 29227 31773 29236 31807
rect 29184 31764 29236 31773
rect 29828 31764 29880 31816
rect 30104 31807 30156 31816
rect 30104 31773 30113 31807
rect 30113 31773 30147 31807
rect 30147 31773 30156 31807
rect 30104 31764 30156 31773
rect 30472 31807 30524 31816
rect 30472 31773 30481 31807
rect 30481 31773 30515 31807
rect 30515 31773 30524 31807
rect 30472 31764 30524 31773
rect 34152 31832 34204 31884
rect 14464 31671 14516 31680
rect 14464 31637 14473 31671
rect 14473 31637 14507 31671
rect 14507 31637 14516 31671
rect 14464 31628 14516 31637
rect 15936 31628 15988 31680
rect 16304 31628 16356 31680
rect 18880 31696 18932 31748
rect 25780 31696 25832 31748
rect 26976 31696 27028 31748
rect 30656 31696 30708 31748
rect 22560 31628 22612 31680
rect 24400 31671 24452 31680
rect 24400 31637 24409 31671
rect 24409 31637 24443 31671
rect 24443 31637 24452 31671
rect 24400 31628 24452 31637
rect 24492 31628 24544 31680
rect 27896 31671 27948 31680
rect 27896 31637 27905 31671
rect 27905 31637 27939 31671
rect 27939 31637 27948 31671
rect 27896 31628 27948 31637
rect 30288 31628 30340 31680
rect 33968 31764 34020 31816
rect 35440 31875 35492 31884
rect 35440 31841 35449 31875
rect 35449 31841 35483 31875
rect 35483 31841 35492 31875
rect 35440 31832 35492 31841
rect 32864 31739 32916 31748
rect 32864 31705 32873 31739
rect 32873 31705 32907 31739
rect 32907 31705 32916 31739
rect 32864 31696 32916 31705
rect 33600 31628 33652 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 13176 31424 13228 31476
rect 13544 31424 13596 31476
rect 9404 31356 9456 31408
rect 14832 31424 14884 31476
rect 15936 31467 15988 31476
rect 15936 31433 15945 31467
rect 15945 31433 15979 31467
rect 15979 31433 15988 31467
rect 15936 31424 15988 31433
rect 17040 31424 17092 31476
rect 14464 31399 14516 31408
rect 14464 31365 14473 31399
rect 14473 31365 14507 31399
rect 14507 31365 14516 31399
rect 14464 31356 14516 31365
rect 16304 31356 16356 31408
rect 19064 31424 19116 31476
rect 22100 31424 22152 31476
rect 8116 31263 8168 31272
rect 8116 31229 8125 31263
rect 8125 31229 8159 31263
rect 8159 31229 8168 31263
rect 8116 31220 8168 31229
rect 8944 31220 8996 31272
rect 9680 31084 9732 31136
rect 14188 31331 14240 31340
rect 14188 31297 14197 31331
rect 14197 31297 14231 31331
rect 14231 31297 14240 31331
rect 14188 31288 14240 31297
rect 17960 31288 18012 31340
rect 18880 31356 18932 31408
rect 22192 31356 22244 31408
rect 22560 31356 22612 31408
rect 24492 31424 24544 31476
rect 25780 31467 25832 31476
rect 25780 31433 25789 31467
rect 25789 31433 25823 31467
rect 25823 31433 25832 31467
rect 25780 31424 25832 31433
rect 29000 31424 29052 31476
rect 32864 31424 32916 31476
rect 24400 31356 24452 31408
rect 25320 31356 25372 31408
rect 27528 31356 27580 31408
rect 27712 31356 27764 31408
rect 30288 31399 30340 31408
rect 30288 31365 30297 31399
rect 30297 31365 30331 31399
rect 30331 31365 30340 31399
rect 30288 31356 30340 31365
rect 26332 31288 26384 31340
rect 13820 31220 13872 31272
rect 17408 31263 17460 31272
rect 17408 31229 17417 31263
rect 17417 31229 17451 31263
rect 17451 31229 17460 31263
rect 17408 31220 17460 31229
rect 18328 31263 18380 31272
rect 18328 31229 18337 31263
rect 18337 31229 18371 31263
rect 18371 31229 18380 31263
rect 18328 31220 18380 31229
rect 19064 31220 19116 31272
rect 16396 31152 16448 31204
rect 9956 31084 10008 31136
rect 16028 31084 16080 31136
rect 19340 31084 19392 31136
rect 19616 31084 19668 31136
rect 20168 31263 20220 31272
rect 20168 31229 20177 31263
rect 20177 31229 20211 31263
rect 20211 31229 20220 31263
rect 20168 31220 20220 31229
rect 24400 31220 24452 31272
rect 25780 31220 25832 31272
rect 26056 31220 26108 31272
rect 26516 31263 26568 31272
rect 26516 31229 26525 31263
rect 26525 31229 26559 31263
rect 26559 31229 26568 31263
rect 26516 31220 26568 31229
rect 27252 31263 27304 31272
rect 27252 31229 27261 31263
rect 27261 31229 27295 31263
rect 27295 31229 27304 31263
rect 27252 31220 27304 31229
rect 28908 31220 28960 31272
rect 30564 31331 30616 31340
rect 30564 31297 30573 31331
rect 30573 31297 30607 31331
rect 30607 31297 30616 31331
rect 30564 31288 30616 31297
rect 31668 31288 31720 31340
rect 32312 31288 32364 31340
rect 34796 31356 34848 31408
rect 34520 31331 34572 31340
rect 34520 31297 34529 31331
rect 34529 31297 34563 31331
rect 34563 31297 34572 31331
rect 34520 31288 34572 31297
rect 34612 31331 34664 31340
rect 34612 31297 34621 31331
rect 34621 31297 34655 31331
rect 34655 31297 34664 31331
rect 34612 31288 34664 31297
rect 29644 31220 29696 31272
rect 32588 31220 32640 31272
rect 33140 31263 33192 31272
rect 33140 31229 33149 31263
rect 33149 31229 33183 31263
rect 33183 31229 33192 31263
rect 33140 31220 33192 31229
rect 25872 31127 25924 31136
rect 25872 31093 25881 31127
rect 25881 31093 25915 31127
rect 25915 31093 25924 31127
rect 25872 31084 25924 31093
rect 27896 31084 27948 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 8944 30923 8996 30932
rect 8944 30889 8953 30923
rect 8953 30889 8987 30923
rect 8987 30889 8996 30923
rect 8944 30880 8996 30889
rect 13360 30880 13412 30932
rect 3516 30676 3568 30728
rect 5632 30744 5684 30796
rect 8208 30744 8260 30796
rect 8576 30744 8628 30796
rect 16396 30880 16448 30932
rect 18328 30880 18380 30932
rect 20168 30880 20220 30932
rect 22468 30880 22520 30932
rect 19340 30812 19392 30864
rect 15292 30744 15344 30796
rect 16488 30744 16540 30796
rect 18236 30744 18288 30796
rect 20260 30812 20312 30864
rect 26332 30880 26384 30932
rect 27252 30880 27304 30932
rect 30380 30880 30432 30932
rect 31116 30880 31168 30932
rect 26516 30812 26568 30864
rect 20904 30787 20956 30796
rect 20904 30753 20913 30787
rect 20913 30753 20947 30787
rect 20947 30753 20956 30787
rect 20904 30744 20956 30753
rect 25872 30744 25924 30796
rect 27988 30744 28040 30796
rect 30564 30744 30616 30796
rect 33048 30812 33100 30864
rect 32404 30744 32456 30796
rect 4620 30676 4672 30728
rect 9772 30719 9824 30728
rect 9772 30685 9781 30719
rect 9781 30685 9815 30719
rect 9815 30685 9824 30719
rect 9772 30676 9824 30685
rect 9956 30719 10008 30728
rect 9956 30685 9965 30719
rect 9965 30685 9999 30719
rect 9999 30685 10008 30719
rect 9956 30676 10008 30685
rect 19616 30719 19668 30728
rect 19616 30685 19625 30719
rect 19625 30685 19659 30719
rect 19659 30685 19668 30719
rect 19616 30676 19668 30685
rect 24400 30719 24452 30728
rect 24400 30685 24409 30719
rect 24409 30685 24443 30719
rect 24443 30685 24452 30719
rect 24400 30676 24452 30685
rect 27896 30676 27948 30728
rect 32588 30719 32640 30728
rect 32588 30685 32597 30719
rect 32597 30685 32631 30719
rect 32631 30685 32640 30719
rect 32588 30676 32640 30685
rect 33600 30719 33652 30728
rect 33600 30685 33609 30719
rect 33609 30685 33643 30719
rect 33643 30685 33652 30719
rect 33600 30676 33652 30685
rect 34612 30676 34664 30728
rect 35348 30676 35400 30728
rect 4712 30608 4764 30660
rect 6368 30651 6420 30660
rect 6368 30617 6377 30651
rect 6377 30617 6411 30651
rect 6411 30617 6420 30651
rect 6368 30608 6420 30617
rect 4160 30540 4212 30592
rect 6736 30540 6788 30592
rect 7472 30608 7524 30660
rect 8300 30540 8352 30592
rect 8484 30583 8536 30592
rect 8484 30549 8493 30583
rect 8493 30549 8527 30583
rect 8527 30549 8536 30583
rect 8484 30540 8536 30549
rect 16028 30608 16080 30660
rect 16304 30608 16356 30660
rect 17592 30651 17644 30660
rect 17592 30617 17601 30651
rect 17601 30617 17635 30651
rect 17635 30617 17644 30651
rect 17592 30608 17644 30617
rect 18880 30608 18932 30660
rect 22100 30608 22152 30660
rect 25228 30608 25280 30660
rect 28908 30608 28960 30660
rect 12624 30540 12676 30592
rect 13176 30583 13228 30592
rect 13176 30549 13185 30583
rect 13185 30549 13219 30583
rect 13219 30549 13228 30583
rect 13176 30540 13228 30549
rect 13728 30540 13780 30592
rect 17960 30540 18012 30592
rect 18328 30540 18380 30592
rect 20812 30540 20864 30592
rect 27620 30540 27672 30592
rect 31116 30608 31168 30660
rect 31576 30608 31628 30660
rect 31944 30608 31996 30660
rect 34520 30608 34572 30660
rect 31484 30540 31536 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 4712 30336 4764 30388
rect 6368 30379 6420 30388
rect 6368 30345 6377 30379
rect 6377 30345 6411 30379
rect 6411 30345 6420 30379
rect 6368 30336 6420 30345
rect 8576 30379 8628 30388
rect 2596 30200 2648 30252
rect 5908 30268 5960 30320
rect 7472 30268 7524 30320
rect 8576 30345 8585 30379
rect 8585 30345 8619 30379
rect 8619 30345 8628 30379
rect 8576 30336 8628 30345
rect 9588 30336 9640 30388
rect 8760 30311 8812 30320
rect 8760 30277 8787 30311
rect 8787 30277 8812 30311
rect 8760 30268 8812 30277
rect 2964 30200 3016 30252
rect 3332 30243 3384 30252
rect 3332 30209 3341 30243
rect 3341 30209 3375 30243
rect 3375 30209 3384 30243
rect 3332 30200 3384 30209
rect 5632 30243 5684 30252
rect 5632 30209 5641 30243
rect 5641 30209 5675 30243
rect 5675 30209 5684 30243
rect 5632 30200 5684 30209
rect 5816 30243 5868 30252
rect 5816 30209 5825 30243
rect 5825 30209 5859 30243
rect 5859 30209 5868 30243
rect 5816 30200 5868 30209
rect 7840 30200 7892 30252
rect 8116 30243 8168 30252
rect 8116 30209 8125 30243
rect 8125 30209 8159 30243
rect 8159 30209 8168 30243
rect 8116 30200 8168 30209
rect 3792 30132 3844 30184
rect 5724 30175 5776 30184
rect 5724 30141 5733 30175
rect 5733 30141 5767 30175
rect 5767 30141 5776 30175
rect 5724 30132 5776 30141
rect 6736 30064 6788 30116
rect 8300 30107 8352 30116
rect 8300 30073 8309 30107
rect 8309 30073 8343 30107
rect 8343 30073 8352 30107
rect 8300 30064 8352 30073
rect 9680 30268 9732 30320
rect 13268 30268 13320 30320
rect 16212 30336 16264 30388
rect 17592 30336 17644 30388
rect 18236 30379 18288 30388
rect 18236 30345 18245 30379
rect 18245 30345 18279 30379
rect 18279 30345 18288 30379
rect 18236 30336 18288 30345
rect 18328 30379 18380 30388
rect 18328 30345 18337 30379
rect 18337 30345 18371 30379
rect 18371 30345 18380 30379
rect 18328 30336 18380 30345
rect 26332 30379 26384 30388
rect 26332 30345 26341 30379
rect 26341 30345 26375 30379
rect 26375 30345 26384 30379
rect 26332 30336 26384 30345
rect 32404 30379 32456 30388
rect 32404 30345 32413 30379
rect 32413 30345 32447 30379
rect 32447 30345 32456 30379
rect 32404 30336 32456 30345
rect 15292 30268 15344 30320
rect 9404 30243 9456 30252
rect 9404 30209 9413 30243
rect 9413 30209 9447 30243
rect 9447 30209 9456 30243
rect 9404 30200 9456 30209
rect 10784 30200 10836 30252
rect 11612 30243 11664 30252
rect 11612 30209 11621 30243
rect 11621 30209 11655 30243
rect 11655 30209 11664 30243
rect 11612 30200 11664 30209
rect 22192 30268 22244 30320
rect 24400 30200 24452 30252
rect 9128 30132 9180 30184
rect 9772 30132 9824 30184
rect 10508 30175 10560 30184
rect 10508 30141 10517 30175
rect 10517 30141 10551 30175
rect 10551 30141 10560 30175
rect 10508 30132 10560 30141
rect 9220 30064 9272 30116
rect 12624 30132 12676 30184
rect 15200 30175 15252 30184
rect 15200 30141 15209 30175
rect 15209 30141 15243 30175
rect 15243 30141 15252 30175
rect 15200 30132 15252 30141
rect 18420 30175 18472 30184
rect 18420 30141 18429 30175
rect 18429 30141 18463 30175
rect 18463 30141 18472 30175
rect 18420 30132 18472 30141
rect 20904 30132 20956 30184
rect 23664 30175 23716 30184
rect 23664 30141 23673 30175
rect 23673 30141 23707 30175
rect 23707 30141 23716 30175
rect 23664 30132 23716 30141
rect 25044 30132 25096 30184
rect 26516 30175 26568 30184
rect 26516 30141 26525 30175
rect 26525 30141 26559 30175
rect 26559 30141 26568 30175
rect 26516 30132 26568 30141
rect 24860 30064 24912 30116
rect 4712 29996 4764 30048
rect 5172 30039 5224 30048
rect 5172 30005 5181 30039
rect 5181 30005 5215 30039
rect 5215 30005 5224 30039
rect 5172 29996 5224 30005
rect 8484 29996 8536 30048
rect 9496 29996 9548 30048
rect 9956 29996 10008 30048
rect 12992 29996 13044 30048
rect 13176 29996 13228 30048
rect 13728 30039 13780 30048
rect 13728 30005 13737 30039
rect 13737 30005 13771 30039
rect 13771 30005 13780 30039
rect 13728 29996 13780 30005
rect 22560 29996 22612 30048
rect 25872 30039 25924 30048
rect 25872 30005 25881 30039
rect 25881 30005 25915 30039
rect 25915 30005 25924 30039
rect 25872 29996 25924 30005
rect 30564 30268 30616 30320
rect 31576 30200 31628 30252
rect 33508 30336 33560 30388
rect 33968 30336 34020 30388
rect 34520 30268 34572 30320
rect 34152 30243 34204 30252
rect 34152 30209 34161 30243
rect 34161 30209 34195 30243
rect 34195 30209 34204 30243
rect 34152 30200 34204 30209
rect 31484 30132 31536 30184
rect 30840 29996 30892 30048
rect 31944 30039 31996 30048
rect 31944 30005 31953 30039
rect 31953 30005 31987 30039
rect 31987 30005 31996 30039
rect 31944 29996 31996 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3792 29835 3844 29844
rect 3792 29801 3801 29835
rect 3801 29801 3835 29835
rect 3835 29801 3844 29835
rect 3792 29792 3844 29801
rect 4528 29792 4580 29844
rect 5172 29792 5224 29844
rect 7840 29835 7892 29844
rect 7840 29801 7849 29835
rect 7849 29801 7883 29835
rect 7883 29801 7892 29835
rect 7840 29792 7892 29801
rect 8116 29835 8168 29844
rect 8116 29801 8125 29835
rect 8125 29801 8159 29835
rect 8159 29801 8168 29835
rect 8116 29792 8168 29801
rect 8208 29792 8260 29844
rect 4528 29656 4580 29708
rect 4712 29656 4764 29708
rect 1400 29588 1452 29640
rect 4252 29588 4304 29640
rect 4620 29588 4672 29640
rect 2596 29520 2648 29572
rect 4896 29631 4948 29640
rect 4896 29597 4905 29631
rect 4905 29597 4939 29631
rect 4939 29597 4948 29631
rect 4896 29588 4948 29597
rect 8484 29724 8536 29776
rect 15200 29792 15252 29844
rect 27620 29835 27672 29844
rect 27620 29801 27629 29835
rect 27629 29801 27663 29835
rect 27663 29801 27672 29835
rect 27620 29792 27672 29801
rect 24768 29724 24820 29776
rect 3608 29495 3660 29504
rect 3608 29461 3617 29495
rect 3617 29461 3651 29495
rect 3651 29461 3660 29495
rect 3608 29452 3660 29461
rect 4160 29452 4212 29504
rect 5540 29520 5592 29572
rect 5908 29520 5960 29572
rect 6092 29452 6144 29504
rect 8300 29631 8352 29640
rect 8300 29597 8309 29631
rect 8309 29597 8343 29631
rect 8343 29597 8352 29631
rect 8300 29588 8352 29597
rect 8484 29631 8536 29640
rect 8484 29597 8493 29631
rect 8493 29597 8527 29631
rect 8527 29597 8536 29631
rect 8484 29588 8536 29597
rect 9956 29699 10008 29708
rect 9956 29665 9965 29699
rect 9965 29665 9999 29699
rect 9999 29665 10008 29699
rect 9956 29656 10008 29665
rect 10416 29656 10468 29708
rect 9220 29588 9272 29640
rect 8760 29520 8812 29572
rect 9404 29520 9456 29572
rect 8484 29452 8536 29504
rect 9128 29452 9180 29504
rect 9312 29495 9364 29504
rect 9312 29461 9321 29495
rect 9321 29461 9355 29495
rect 9355 29461 9364 29495
rect 9312 29452 9364 29461
rect 10416 29520 10468 29572
rect 13820 29656 13872 29708
rect 14648 29699 14700 29708
rect 14648 29665 14657 29699
rect 14657 29665 14691 29699
rect 14691 29665 14700 29699
rect 14648 29656 14700 29665
rect 16488 29656 16540 29708
rect 20904 29656 20956 29708
rect 25044 29699 25096 29708
rect 25044 29665 25053 29699
rect 25053 29665 25087 29699
rect 25087 29665 25096 29699
rect 25044 29656 25096 29665
rect 25228 29724 25280 29776
rect 11520 29631 11572 29640
rect 11520 29597 11529 29631
rect 11529 29597 11563 29631
rect 11563 29597 11572 29631
rect 11520 29588 11572 29597
rect 10600 29452 10652 29504
rect 11796 29563 11848 29572
rect 11796 29529 11805 29563
rect 11805 29529 11839 29563
rect 11839 29529 11848 29563
rect 11796 29520 11848 29529
rect 13268 29588 13320 29640
rect 13728 29588 13780 29640
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 20812 29588 20864 29640
rect 22192 29588 22244 29640
rect 25412 29588 25464 29640
rect 16212 29520 16264 29572
rect 17224 29563 17276 29572
rect 17224 29529 17233 29563
rect 17233 29529 17267 29563
rect 17267 29529 17276 29563
rect 17224 29520 17276 29529
rect 19524 29563 19576 29572
rect 19524 29529 19533 29563
rect 19533 29529 19567 29563
rect 19567 29529 19576 29563
rect 19524 29520 19576 29529
rect 23296 29563 23348 29572
rect 23296 29529 23305 29563
rect 23305 29529 23339 29563
rect 23339 29529 23348 29563
rect 23296 29520 23348 29529
rect 13268 29495 13320 29504
rect 13268 29461 13277 29495
rect 13277 29461 13311 29495
rect 13311 29461 13320 29495
rect 13268 29452 13320 29461
rect 15660 29452 15712 29504
rect 15752 29495 15804 29504
rect 15752 29461 15761 29495
rect 15761 29461 15795 29495
rect 15795 29461 15804 29495
rect 15752 29452 15804 29461
rect 20168 29452 20220 29504
rect 22652 29452 22704 29504
rect 25136 29520 25188 29572
rect 24768 29452 24820 29504
rect 25780 29656 25832 29708
rect 29092 29656 29144 29708
rect 31760 29588 31812 29640
rect 33048 29656 33100 29708
rect 33876 29656 33928 29708
rect 34612 29588 34664 29640
rect 26608 29520 26660 29572
rect 27988 29520 28040 29572
rect 27620 29452 27672 29504
rect 29552 29495 29604 29504
rect 29552 29461 29561 29495
rect 29561 29461 29595 29495
rect 29595 29461 29604 29495
rect 29552 29452 29604 29461
rect 29920 29495 29972 29504
rect 29920 29461 29929 29495
rect 29929 29461 29963 29495
rect 29963 29461 29972 29495
rect 29920 29452 29972 29461
rect 30104 29452 30156 29504
rect 32496 29452 32548 29504
rect 33416 29452 33468 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 2964 29180 3016 29232
rect 4252 29291 4304 29300
rect 4252 29257 4261 29291
rect 4261 29257 4295 29291
rect 4295 29257 4304 29291
rect 4252 29248 4304 29257
rect 3976 29180 4028 29232
rect 1400 29087 1452 29096
rect 1400 29053 1409 29087
rect 1409 29053 1443 29087
rect 1443 29053 1452 29087
rect 1400 29044 1452 29053
rect 1676 29087 1728 29096
rect 1676 29053 1685 29087
rect 1685 29053 1719 29087
rect 1719 29053 1728 29087
rect 1676 29044 1728 29053
rect 2872 28976 2924 29028
rect 5356 29180 5408 29232
rect 5540 29291 5592 29300
rect 5540 29257 5549 29291
rect 5549 29257 5583 29291
rect 5583 29257 5592 29291
rect 5540 29248 5592 29257
rect 5908 29248 5960 29300
rect 6460 29248 6512 29300
rect 5816 29180 5868 29232
rect 9312 29248 9364 29300
rect 10508 29291 10560 29300
rect 10508 29257 10517 29291
rect 10517 29257 10551 29291
rect 10551 29257 10560 29291
rect 10508 29248 10560 29257
rect 10784 29223 10836 29232
rect 10784 29189 10793 29223
rect 10793 29189 10827 29223
rect 10827 29189 10836 29223
rect 10784 29180 10836 29189
rect 5724 29155 5776 29164
rect 5724 29121 5733 29155
rect 5733 29121 5767 29155
rect 5767 29121 5776 29155
rect 5724 29112 5776 29121
rect 6092 29112 6144 29164
rect 3608 28908 3660 28960
rect 5908 28951 5960 28960
rect 5908 28917 5917 28951
rect 5917 28917 5951 28951
rect 5951 28917 5960 28951
rect 5908 28908 5960 28917
rect 7748 29087 7800 29096
rect 7748 29053 7757 29087
rect 7757 29053 7791 29087
rect 7791 29053 7800 29087
rect 7748 29044 7800 29053
rect 9220 29019 9272 29028
rect 9220 28985 9229 29019
rect 9229 28985 9263 29019
rect 9263 28985 9272 29019
rect 10600 29155 10652 29164
rect 10600 29121 10609 29155
rect 10609 29121 10643 29155
rect 10643 29121 10652 29155
rect 10600 29112 10652 29121
rect 11796 29248 11848 29300
rect 13268 29248 13320 29300
rect 15660 29291 15712 29300
rect 15660 29257 15669 29291
rect 15669 29257 15703 29291
rect 15703 29257 15712 29291
rect 15660 29248 15712 29257
rect 17224 29248 17276 29300
rect 19524 29248 19576 29300
rect 20168 29248 20220 29300
rect 22192 29248 22244 29300
rect 12992 29223 13044 29232
rect 12992 29189 13001 29223
rect 13001 29189 13035 29223
rect 13035 29189 13044 29223
rect 12992 29180 13044 29189
rect 16212 29180 16264 29232
rect 23480 29248 23532 29300
rect 24768 29248 24820 29300
rect 26608 29248 26660 29300
rect 27528 29248 27580 29300
rect 28908 29248 28960 29300
rect 23848 29180 23900 29232
rect 25136 29223 25188 29232
rect 25136 29189 25145 29223
rect 25145 29189 25179 29223
rect 25179 29189 25188 29223
rect 25136 29180 25188 29189
rect 30104 29248 30156 29300
rect 34612 29248 34664 29300
rect 9680 29087 9732 29096
rect 9680 29053 9689 29087
rect 9689 29053 9723 29087
rect 9723 29053 9732 29087
rect 9680 29044 9732 29053
rect 9772 29044 9824 29096
rect 15752 29112 15804 29164
rect 17316 29112 17368 29164
rect 19892 29112 19944 29164
rect 21272 29155 21324 29164
rect 21272 29121 21281 29155
rect 21281 29121 21315 29155
rect 21315 29121 21324 29155
rect 21272 29112 21324 29121
rect 22652 29112 22704 29164
rect 25412 29155 25464 29164
rect 25412 29121 25421 29155
rect 25421 29121 25455 29155
rect 25455 29121 25464 29155
rect 25412 29112 25464 29121
rect 26148 29112 26200 29164
rect 13176 29087 13228 29096
rect 13176 29053 13185 29087
rect 13185 29053 13219 29087
rect 13219 29053 13228 29087
rect 13176 29044 13228 29053
rect 9220 28976 9272 28985
rect 10232 28976 10284 29028
rect 8208 28908 8260 28960
rect 9588 28951 9640 28960
rect 9588 28917 9597 28951
rect 9597 28917 9631 28951
rect 9631 28917 9640 28951
rect 9588 28908 9640 28917
rect 14188 29087 14240 29096
rect 14188 29053 14197 29087
rect 14197 29053 14231 29087
rect 14231 29053 14240 29087
rect 14188 29044 14240 29053
rect 14648 29044 14700 29096
rect 16856 29044 16908 29096
rect 20260 29087 20312 29096
rect 20260 29053 20269 29087
rect 20269 29053 20303 29087
rect 20303 29053 20312 29087
rect 20260 29044 20312 29053
rect 20904 29044 20956 29096
rect 21456 29087 21508 29096
rect 21456 29053 21465 29087
rect 21465 29053 21499 29087
rect 21499 29053 21508 29087
rect 21456 29044 21508 29053
rect 27252 29087 27304 29096
rect 27252 29053 27261 29087
rect 27261 29053 27295 29087
rect 27295 29053 27304 29087
rect 27252 29044 27304 29053
rect 30472 29087 30524 29096
rect 30472 29053 30481 29087
rect 30481 29053 30515 29087
rect 30515 29053 30524 29087
rect 30472 29044 30524 29053
rect 17960 28976 18012 29028
rect 18420 28976 18472 29028
rect 30840 29087 30892 29096
rect 30840 29053 30849 29087
rect 30849 29053 30883 29087
rect 30883 29053 30892 29087
rect 30840 29044 30892 29053
rect 32496 29223 32548 29232
rect 32496 29189 32505 29223
rect 32505 29189 32539 29223
rect 32539 29189 32548 29223
rect 32496 29180 32548 29189
rect 33508 29180 33560 29232
rect 31392 29112 31444 29164
rect 31944 29112 31996 29164
rect 31852 28976 31904 29028
rect 33140 29044 33192 29096
rect 14740 28908 14792 28960
rect 18788 28908 18840 28960
rect 20720 28908 20772 28960
rect 27620 28908 27672 28960
rect 29000 28951 29052 28960
rect 29000 28917 29009 28951
rect 29009 28917 29043 28951
rect 29043 28917 29052 28951
rect 29000 28908 29052 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1676 28704 1728 28756
rect 2872 28543 2924 28552
rect 2872 28509 2881 28543
rect 2881 28509 2915 28543
rect 2915 28509 2924 28543
rect 2872 28500 2924 28509
rect 3608 28568 3660 28620
rect 4068 28704 4120 28756
rect 6000 28747 6052 28756
rect 6000 28713 6009 28747
rect 6009 28713 6043 28747
rect 6043 28713 6052 28747
rect 6000 28704 6052 28713
rect 6736 28704 6788 28756
rect 7748 28704 7800 28756
rect 8300 28747 8352 28756
rect 8300 28713 8309 28747
rect 8309 28713 8343 28747
rect 8343 28713 8352 28747
rect 8300 28704 8352 28713
rect 14188 28704 14240 28756
rect 17316 28747 17368 28756
rect 17316 28713 17325 28747
rect 17325 28713 17359 28747
rect 17359 28713 17368 28747
rect 17316 28704 17368 28713
rect 21272 28704 21324 28756
rect 23296 28704 23348 28756
rect 23664 28704 23716 28756
rect 4804 28636 4856 28688
rect 3976 28611 4028 28620
rect 3976 28577 3985 28611
rect 3985 28577 4019 28611
rect 4019 28577 4028 28611
rect 3976 28568 4028 28577
rect 3516 28432 3568 28484
rect 3700 28432 3752 28484
rect 4620 28500 4672 28552
rect 13176 28611 13228 28620
rect 13176 28577 13185 28611
rect 13185 28577 13219 28611
rect 13219 28577 13228 28611
rect 13176 28568 13228 28577
rect 16396 28568 16448 28620
rect 18788 28611 18840 28620
rect 18788 28577 18797 28611
rect 18797 28577 18831 28611
rect 18831 28577 18840 28611
rect 18788 28568 18840 28577
rect 19248 28568 19300 28620
rect 19340 28568 19392 28620
rect 20720 28611 20772 28620
rect 20720 28577 20729 28611
rect 20729 28577 20763 28611
rect 20763 28577 20772 28611
rect 20720 28568 20772 28577
rect 21456 28568 21508 28620
rect 22560 28611 22612 28620
rect 22560 28577 22569 28611
rect 22569 28577 22603 28611
rect 22603 28577 22612 28611
rect 22560 28568 22612 28577
rect 27252 28747 27304 28756
rect 27252 28713 27261 28747
rect 27261 28713 27295 28747
rect 27295 28713 27304 28747
rect 27252 28704 27304 28713
rect 30472 28704 30524 28756
rect 26516 28636 26568 28688
rect 25872 28611 25924 28620
rect 25872 28577 25881 28611
rect 25881 28577 25915 28611
rect 25915 28577 25924 28611
rect 25872 28568 25924 28577
rect 26148 28611 26200 28620
rect 26148 28577 26157 28611
rect 26157 28577 26191 28611
rect 26191 28577 26200 28611
rect 26148 28568 26200 28577
rect 27988 28568 28040 28620
rect 29092 28636 29144 28688
rect 30104 28679 30156 28688
rect 30104 28645 30113 28679
rect 30113 28645 30147 28679
rect 30147 28645 30156 28679
rect 30104 28636 30156 28645
rect 29276 28568 29328 28620
rect 29920 28568 29972 28620
rect 30840 28568 30892 28620
rect 33416 28611 33468 28620
rect 33416 28577 33425 28611
rect 33425 28577 33459 28611
rect 33459 28577 33468 28611
rect 33416 28568 33468 28577
rect 8116 28543 8168 28552
rect 8116 28509 8125 28543
rect 8125 28509 8159 28543
rect 8159 28509 8168 28543
rect 8116 28500 8168 28509
rect 8760 28500 8812 28552
rect 13268 28500 13320 28552
rect 15660 28500 15712 28552
rect 22652 28543 22704 28552
rect 22652 28509 22661 28543
rect 22661 28509 22695 28543
rect 22695 28509 22704 28543
rect 22652 28500 22704 28509
rect 23480 28500 23532 28552
rect 27620 28543 27672 28552
rect 27620 28509 27629 28543
rect 27629 28509 27663 28543
rect 27663 28509 27672 28543
rect 27620 28500 27672 28509
rect 29000 28543 29052 28552
rect 29000 28509 29009 28543
rect 29009 28509 29043 28543
rect 29043 28509 29052 28543
rect 29000 28500 29052 28509
rect 31852 28543 31904 28552
rect 31852 28509 31861 28543
rect 31861 28509 31895 28543
rect 31895 28509 31904 28543
rect 31852 28500 31904 28509
rect 5724 28432 5776 28484
rect 6092 28432 6144 28484
rect 15752 28432 15804 28484
rect 18328 28432 18380 28484
rect 19892 28475 19944 28484
rect 19892 28441 19901 28475
rect 19901 28441 19935 28475
rect 19935 28441 19944 28475
rect 19892 28432 19944 28441
rect 20168 28432 20220 28484
rect 20812 28432 20864 28484
rect 23848 28432 23900 28484
rect 30932 28432 30984 28484
rect 32680 28475 32732 28484
rect 32680 28441 32689 28475
rect 32689 28441 32723 28475
rect 32723 28441 32732 28475
rect 32680 28432 32732 28441
rect 33968 28500 34020 28552
rect 33784 28432 33836 28484
rect 35348 28432 35400 28484
rect 2228 28364 2280 28416
rect 4528 28364 4580 28416
rect 5356 28364 5408 28416
rect 5816 28407 5868 28416
rect 5816 28373 5825 28407
rect 5825 28373 5859 28407
rect 5859 28373 5868 28407
rect 5816 28364 5868 28373
rect 11980 28364 12032 28416
rect 13452 28364 13504 28416
rect 19524 28407 19576 28416
rect 19524 28373 19533 28407
rect 19533 28373 19567 28407
rect 19567 28373 19576 28407
rect 19524 28364 19576 28373
rect 22560 28364 22612 28416
rect 25044 28364 25096 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 2872 28160 2924 28212
rect 5908 28160 5960 28212
rect 6092 28160 6144 28212
rect 2228 28067 2280 28076
rect 2228 28033 2237 28067
rect 2237 28033 2271 28067
rect 2271 28033 2280 28067
rect 2228 28024 2280 28033
rect 3424 28135 3476 28144
rect 3424 28101 3433 28135
rect 3433 28101 3467 28135
rect 3467 28101 3476 28135
rect 3424 28092 3476 28101
rect 3700 28092 3752 28144
rect 5264 28135 5316 28144
rect 5264 28101 5273 28135
rect 5273 28101 5307 28135
rect 5307 28101 5316 28135
rect 5264 28092 5316 28101
rect 5356 28092 5408 28144
rect 5724 28135 5776 28144
rect 5724 28101 5733 28135
rect 5733 28101 5767 28135
rect 5767 28101 5776 28135
rect 5724 28092 5776 28101
rect 3056 27956 3108 28008
rect 3608 28024 3660 28076
rect 3976 28067 4028 28076
rect 3976 28033 3985 28067
rect 3985 28033 4019 28067
rect 4019 28033 4028 28067
rect 3976 28024 4028 28033
rect 4068 28024 4120 28076
rect 4528 28024 4580 28076
rect 16856 28160 16908 28212
rect 29276 28160 29328 28212
rect 33416 28160 33468 28212
rect 5908 27999 5960 28008
rect 5908 27965 5917 27999
rect 5917 27965 5951 27999
rect 5951 27965 5960 27999
rect 5908 27956 5960 27965
rect 6828 27999 6880 28008
rect 6828 27965 6837 27999
rect 6837 27965 6871 27999
rect 6871 27965 6880 27999
rect 6828 27956 6880 27965
rect 8208 27956 8260 28008
rect 9036 27999 9088 28008
rect 9036 27965 9045 27999
rect 9045 27965 9079 27999
rect 9079 27965 9088 27999
rect 9036 27956 9088 27965
rect 9128 27956 9180 28008
rect 5632 27888 5684 27940
rect 6000 27888 6052 27940
rect 10048 27888 10100 27940
rect 11980 28135 12032 28144
rect 11980 28101 11989 28135
rect 11989 28101 12023 28135
rect 12023 28101 12032 28135
rect 11980 28092 12032 28101
rect 11520 28024 11572 28076
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 12440 27956 12492 28008
rect 13728 28092 13780 28144
rect 18236 28092 18288 28144
rect 28908 28092 28960 28144
rect 29552 28092 29604 28144
rect 32680 28092 32732 28144
rect 33140 28092 33192 28144
rect 16120 28024 16172 28076
rect 22652 28024 22704 28076
rect 25136 28024 25188 28076
rect 30012 28024 30064 28076
rect 30932 28067 30984 28076
rect 30932 28033 30941 28067
rect 30941 28033 30975 28067
rect 30975 28033 30984 28067
rect 30932 28024 30984 28033
rect 14740 27999 14792 28008
rect 14740 27965 14749 27999
rect 14749 27965 14783 27999
rect 14783 27965 14792 27999
rect 14740 27956 14792 27965
rect 16304 27956 16356 28008
rect 18144 27999 18196 28008
rect 18144 27965 18153 27999
rect 18153 27965 18187 27999
rect 18187 27965 18196 27999
rect 18144 27956 18196 27965
rect 19248 27956 19300 28008
rect 19340 27956 19392 28008
rect 25964 27956 26016 28008
rect 25504 27888 25556 27940
rect 30104 27956 30156 28008
rect 31024 27956 31076 28008
rect 31300 27956 31352 28008
rect 31852 27956 31904 28008
rect 30472 27888 30524 27940
rect 31760 27888 31812 27940
rect 2136 27820 2188 27872
rect 3148 27820 3200 27872
rect 4620 27820 4672 27872
rect 5448 27863 5500 27872
rect 5448 27829 5457 27863
rect 5457 27829 5491 27863
rect 5491 27829 5500 27863
rect 5448 27820 5500 27829
rect 6092 27820 6144 27872
rect 6276 27820 6328 27872
rect 10784 27820 10836 27872
rect 13452 27863 13504 27872
rect 13452 27829 13461 27863
rect 13461 27829 13495 27863
rect 13495 27829 13504 27863
rect 13452 27820 13504 27829
rect 15200 27820 15252 27872
rect 16120 27820 16172 27872
rect 16672 27863 16724 27872
rect 16672 27829 16681 27863
rect 16681 27829 16715 27863
rect 16715 27829 16724 27863
rect 16672 27820 16724 27829
rect 25872 27820 25924 27872
rect 30656 27820 30708 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2136 27659 2188 27668
rect 2136 27625 2166 27659
rect 2166 27625 2188 27659
rect 2136 27616 2188 27625
rect 3608 27659 3660 27668
rect 3608 27625 3617 27659
rect 3617 27625 3651 27659
rect 3651 27625 3660 27659
rect 3608 27616 3660 27625
rect 4620 27616 4672 27668
rect 5724 27616 5776 27668
rect 6828 27616 6880 27668
rect 9036 27616 9088 27668
rect 18144 27616 18196 27668
rect 3424 27548 3476 27600
rect 4068 27548 4120 27600
rect 6552 27548 6604 27600
rect 3148 27480 3200 27532
rect 6092 27480 6144 27532
rect 8208 27480 8260 27532
rect 10600 27480 10652 27532
rect 16304 27591 16356 27600
rect 16304 27557 16313 27591
rect 16313 27557 16347 27591
rect 16347 27557 16356 27591
rect 16304 27548 16356 27557
rect 16396 27548 16448 27600
rect 19340 27616 19392 27668
rect 19524 27659 19576 27668
rect 19524 27625 19554 27659
rect 19554 27625 19576 27659
rect 19524 27616 19576 27625
rect 19892 27616 19944 27668
rect 11796 27480 11848 27532
rect 12808 27480 12860 27532
rect 14832 27480 14884 27532
rect 1400 27412 1452 27464
rect 1860 27455 1912 27464
rect 1860 27421 1869 27455
rect 1869 27421 1903 27455
rect 1903 27421 1912 27455
rect 1860 27412 1912 27421
rect 3608 27412 3660 27464
rect 5448 27455 5500 27464
rect 5448 27421 5457 27455
rect 5457 27421 5491 27455
rect 5491 27421 5500 27455
rect 5448 27412 5500 27421
rect 5540 27412 5592 27464
rect 5816 27412 5868 27464
rect 2872 27344 2924 27396
rect 9128 27412 9180 27464
rect 5356 27276 5408 27328
rect 6184 27319 6236 27328
rect 6184 27285 6193 27319
rect 6193 27285 6227 27319
rect 6227 27285 6236 27319
rect 6184 27276 6236 27285
rect 6460 27344 6512 27396
rect 9588 27412 9640 27464
rect 10048 27412 10100 27464
rect 10140 27455 10192 27464
rect 10140 27421 10149 27455
rect 10149 27421 10183 27455
rect 10183 27421 10192 27455
rect 10140 27412 10192 27421
rect 10324 27455 10376 27464
rect 10324 27421 10333 27455
rect 10333 27421 10367 27455
rect 10367 27421 10376 27455
rect 10324 27412 10376 27421
rect 16672 27480 16724 27532
rect 25136 27616 25188 27668
rect 25504 27616 25556 27668
rect 32128 27616 32180 27668
rect 33232 27616 33284 27668
rect 33968 27659 34020 27668
rect 33968 27625 33977 27659
rect 33977 27625 34011 27659
rect 34011 27625 34020 27659
rect 33968 27616 34020 27625
rect 16396 27412 16448 27464
rect 17960 27480 18012 27532
rect 18880 27480 18932 27532
rect 19248 27523 19300 27532
rect 19248 27489 19257 27523
rect 19257 27489 19291 27523
rect 19291 27489 19300 27523
rect 19248 27480 19300 27489
rect 22652 27523 22704 27532
rect 22652 27489 22661 27523
rect 22661 27489 22695 27523
rect 22695 27489 22704 27523
rect 22652 27480 22704 27489
rect 24860 27523 24912 27532
rect 24860 27489 24869 27523
rect 24869 27489 24903 27523
rect 24903 27489 24912 27523
rect 24860 27480 24912 27489
rect 26148 27480 26200 27532
rect 30472 27480 30524 27532
rect 10508 27344 10560 27396
rect 10876 27344 10928 27396
rect 11060 27344 11112 27396
rect 12440 27387 12492 27396
rect 12440 27353 12449 27387
rect 12449 27353 12483 27387
rect 12483 27353 12492 27387
rect 12440 27344 12492 27353
rect 13728 27344 13780 27396
rect 6920 27276 6972 27328
rect 8116 27276 8168 27328
rect 10968 27276 11020 27328
rect 13360 27276 13412 27328
rect 14096 27319 14148 27328
rect 14096 27285 14105 27319
rect 14105 27285 14139 27319
rect 14139 27285 14148 27319
rect 14096 27276 14148 27285
rect 15108 27344 15160 27396
rect 15568 27387 15620 27396
rect 15568 27353 15577 27387
rect 15577 27353 15611 27387
rect 15611 27353 15620 27387
rect 15568 27344 15620 27353
rect 16856 27344 16908 27396
rect 17316 27344 17368 27396
rect 20812 27344 20864 27396
rect 20444 27276 20496 27328
rect 24768 27412 24820 27464
rect 26976 27412 27028 27464
rect 31300 27455 31352 27464
rect 31300 27421 31309 27455
rect 31309 27421 31343 27455
rect 31343 27421 31352 27455
rect 31300 27412 31352 27421
rect 22192 27344 22244 27396
rect 23296 27344 23348 27396
rect 25136 27387 25188 27396
rect 25136 27353 25145 27387
rect 25145 27353 25179 27387
rect 25179 27353 25188 27387
rect 25136 27344 25188 27353
rect 27528 27344 27580 27396
rect 30564 27344 30616 27396
rect 30748 27344 30800 27396
rect 33140 27344 33192 27396
rect 22100 27319 22152 27328
rect 22100 27285 22109 27319
rect 22109 27285 22143 27319
rect 22143 27285 22152 27319
rect 22100 27276 22152 27285
rect 22468 27319 22520 27328
rect 22468 27285 22477 27319
rect 22477 27285 22511 27319
rect 22511 27285 22520 27319
rect 22468 27276 22520 27285
rect 25320 27276 25372 27328
rect 25964 27276 26016 27328
rect 27712 27319 27764 27328
rect 27712 27285 27721 27319
rect 27721 27285 27755 27319
rect 27755 27285 27764 27319
rect 27712 27276 27764 27285
rect 28172 27319 28224 27328
rect 28172 27285 28181 27319
rect 28181 27285 28215 27319
rect 28215 27285 28224 27319
rect 28172 27276 28224 27285
rect 28448 27276 28500 27328
rect 29184 27276 29236 27328
rect 31024 27276 31076 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 5540 27115 5592 27124
rect 5540 27081 5565 27115
rect 5565 27081 5592 27115
rect 5540 27072 5592 27081
rect 6184 27072 6236 27124
rect 10692 27072 10744 27124
rect 13360 27115 13412 27124
rect 13360 27081 13369 27115
rect 13369 27081 13403 27115
rect 13403 27081 13412 27115
rect 13360 27072 13412 27081
rect 15568 27072 15620 27124
rect 19432 27072 19484 27124
rect 20812 27072 20864 27124
rect 2964 27004 3016 27056
rect 5448 27004 5500 27056
rect 5816 27047 5868 27056
rect 5816 27013 5825 27047
rect 5825 27013 5859 27047
rect 5859 27013 5868 27047
rect 5816 27004 5868 27013
rect 4804 26936 4856 26988
rect 5264 26936 5316 26988
rect 6736 27047 6788 27056
rect 6736 27013 6745 27047
rect 6745 27013 6779 27047
rect 6779 27013 6788 27047
rect 6736 27004 6788 27013
rect 6828 27004 6880 27056
rect 1676 26911 1728 26920
rect 1676 26877 1685 26911
rect 1685 26877 1719 26911
rect 1719 26877 1728 26911
rect 1676 26868 1728 26877
rect 1860 26732 1912 26784
rect 4712 26868 4764 26920
rect 5908 26868 5960 26920
rect 6460 26800 6512 26852
rect 3148 26775 3200 26784
rect 3148 26741 3157 26775
rect 3157 26741 3191 26775
rect 3191 26741 3200 26775
rect 3148 26732 3200 26741
rect 4620 26732 4672 26784
rect 5356 26732 5408 26784
rect 5632 26732 5684 26784
rect 6000 26775 6052 26784
rect 6000 26741 6009 26775
rect 6009 26741 6043 26775
rect 6043 26741 6052 26775
rect 6000 26732 6052 26741
rect 6092 26732 6144 26784
rect 6828 26868 6880 26920
rect 8392 26979 8444 26988
rect 8392 26945 8401 26979
rect 8401 26945 8435 26979
rect 8435 26945 8444 26979
rect 8392 26936 8444 26945
rect 8760 27047 8812 27056
rect 8760 27013 8769 27047
rect 8769 27013 8803 27047
rect 8803 27013 8812 27047
rect 8760 27004 8812 27013
rect 9588 27004 9640 27056
rect 9496 26936 9548 26988
rect 10048 27004 10100 27056
rect 10416 26936 10468 26988
rect 10968 27004 11020 27056
rect 14740 27004 14792 27056
rect 20444 27004 20496 27056
rect 20720 27004 20772 27056
rect 21824 27072 21876 27124
rect 22468 27072 22520 27124
rect 24952 27072 25004 27124
rect 25688 27072 25740 27124
rect 30932 27072 30984 27124
rect 31024 27072 31076 27124
rect 23848 27004 23900 27056
rect 25320 27047 25372 27056
rect 25320 27013 25329 27047
rect 25329 27013 25363 27047
rect 25363 27013 25372 27047
rect 25320 27004 25372 27013
rect 9864 26868 9916 26920
rect 10140 26868 10192 26920
rect 7380 26843 7432 26852
rect 7380 26809 7389 26843
rect 7389 26809 7423 26843
rect 7423 26809 7432 26843
rect 7380 26800 7432 26809
rect 8116 26800 8168 26852
rect 13268 26911 13320 26920
rect 13268 26877 13277 26911
rect 13277 26877 13311 26911
rect 13311 26877 13320 26911
rect 13268 26868 13320 26877
rect 16396 26979 16448 26988
rect 16396 26945 16405 26979
rect 16405 26945 16439 26979
rect 16439 26945 16448 26979
rect 16396 26936 16448 26945
rect 14096 26868 14148 26920
rect 14924 26868 14976 26920
rect 17040 26868 17092 26920
rect 17776 26911 17828 26920
rect 17776 26877 17785 26911
rect 17785 26877 17819 26911
rect 17819 26877 17828 26911
rect 17776 26868 17828 26877
rect 19248 26979 19300 26988
rect 19248 26945 19257 26979
rect 19257 26945 19291 26979
rect 19291 26945 19300 26979
rect 26148 27004 26200 27056
rect 27436 27004 27488 27056
rect 28172 27004 28224 27056
rect 30380 27004 30432 27056
rect 30564 27004 30616 27056
rect 30656 27047 30708 27056
rect 30656 27013 30665 27047
rect 30665 27013 30699 27047
rect 30699 27013 30708 27047
rect 30656 27004 30708 27013
rect 32128 27047 32180 27056
rect 32128 27013 32137 27047
rect 32137 27013 32171 27047
rect 32171 27013 32180 27047
rect 32128 27004 32180 27013
rect 19248 26936 19300 26945
rect 25688 26979 25740 26988
rect 25688 26945 25697 26979
rect 25697 26945 25731 26979
rect 25731 26945 25740 26979
rect 25688 26936 25740 26945
rect 18788 26911 18840 26920
rect 10876 26843 10928 26852
rect 10876 26809 10885 26843
rect 10885 26809 10919 26843
rect 10919 26809 10928 26843
rect 10876 26800 10928 26809
rect 16488 26800 16540 26852
rect 18788 26877 18797 26911
rect 18797 26877 18831 26911
rect 18831 26877 18840 26911
rect 18788 26868 18840 26877
rect 18880 26911 18932 26920
rect 18880 26877 18889 26911
rect 18889 26877 18923 26911
rect 18923 26877 18932 26911
rect 18880 26868 18932 26877
rect 22100 26868 22152 26920
rect 22836 26868 22888 26920
rect 24860 26868 24912 26920
rect 26516 26868 26568 26920
rect 26976 26911 27028 26920
rect 26976 26877 26985 26911
rect 26985 26877 27019 26911
rect 27019 26877 27028 26911
rect 26976 26868 27028 26877
rect 29000 26868 29052 26920
rect 29184 26911 29236 26920
rect 29184 26877 29193 26911
rect 29193 26877 29227 26911
rect 29227 26877 29236 26911
rect 29184 26868 29236 26877
rect 30012 26868 30064 26920
rect 31300 26936 31352 26988
rect 31392 26936 31444 26988
rect 33232 27115 33284 27124
rect 33232 27081 33241 27115
rect 33241 27081 33275 27115
rect 33275 27081 33284 27115
rect 33232 27072 33284 27081
rect 33968 27072 34020 27124
rect 7104 26775 7156 26784
rect 7104 26741 7113 26775
rect 7113 26741 7147 26775
rect 7147 26741 7156 26775
rect 7104 26732 7156 26741
rect 8944 26732 8996 26784
rect 10784 26732 10836 26784
rect 17224 26732 17276 26784
rect 17960 26732 18012 26784
rect 21824 26732 21876 26784
rect 22284 26732 22336 26784
rect 23296 26732 23348 26784
rect 30104 26732 30156 26784
rect 31484 26868 31536 26920
rect 33692 26911 33744 26920
rect 33692 26877 33701 26911
rect 33701 26877 33735 26911
rect 33735 26877 33744 26911
rect 33692 26868 33744 26877
rect 33876 26911 33928 26920
rect 33876 26877 33885 26911
rect 33885 26877 33919 26911
rect 33919 26877 33928 26911
rect 33876 26868 33928 26877
rect 33140 26800 33192 26852
rect 34060 26800 34112 26852
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 1676 26528 1728 26580
rect 4620 26528 4672 26580
rect 5908 26571 5960 26580
rect 5908 26537 5917 26571
rect 5917 26537 5951 26571
rect 5951 26537 5960 26571
rect 5908 26528 5960 26537
rect 6368 26571 6420 26580
rect 6368 26537 6377 26571
rect 6377 26537 6411 26571
rect 6411 26537 6420 26571
rect 6368 26528 6420 26537
rect 8208 26528 8260 26580
rect 8944 26528 8996 26580
rect 5816 26460 5868 26512
rect 9128 26460 9180 26512
rect 9220 26503 9272 26512
rect 9220 26469 9229 26503
rect 9229 26469 9263 26503
rect 9263 26469 9272 26503
rect 9220 26460 9272 26469
rect 3148 26392 3200 26444
rect 4528 26392 4580 26444
rect 6276 26392 6328 26444
rect 6552 26392 6604 26444
rect 7380 26392 7432 26444
rect 10692 26528 10744 26580
rect 12440 26528 12492 26580
rect 17776 26528 17828 26580
rect 22836 26571 22888 26580
rect 22836 26537 22845 26571
rect 22845 26537 22879 26571
rect 22879 26537 22888 26571
rect 22836 26528 22888 26537
rect 25228 26528 25280 26580
rect 27712 26528 27764 26580
rect 31484 26571 31536 26580
rect 31484 26537 31493 26571
rect 31493 26537 31527 26571
rect 31527 26537 31536 26571
rect 31484 26528 31536 26537
rect 13268 26460 13320 26512
rect 5724 26324 5776 26376
rect 8944 26367 8996 26376
rect 8944 26333 8953 26367
rect 8953 26333 8987 26367
rect 8987 26333 8996 26367
rect 8944 26324 8996 26333
rect 9680 26324 9732 26376
rect 13452 26435 13504 26444
rect 13452 26401 13461 26435
rect 13461 26401 13495 26435
rect 13495 26401 13504 26435
rect 13452 26392 13504 26401
rect 16488 26460 16540 26512
rect 14096 26392 14148 26444
rect 14740 26435 14792 26444
rect 14740 26401 14749 26435
rect 14749 26401 14783 26435
rect 14783 26401 14792 26435
rect 14740 26392 14792 26401
rect 16396 26392 16448 26444
rect 19248 26392 19300 26444
rect 10140 26367 10192 26376
rect 10140 26333 10149 26367
rect 10149 26333 10183 26367
rect 10183 26333 10192 26367
rect 10140 26324 10192 26333
rect 10324 26367 10376 26376
rect 10324 26333 10333 26367
rect 10333 26333 10367 26367
rect 10367 26333 10376 26367
rect 10324 26324 10376 26333
rect 13360 26367 13412 26376
rect 13360 26333 13369 26367
rect 13369 26333 13403 26367
rect 13403 26333 13412 26367
rect 13360 26324 13412 26333
rect 14924 26367 14976 26376
rect 14924 26333 14933 26367
rect 14933 26333 14967 26367
rect 14967 26333 14976 26367
rect 14924 26324 14976 26333
rect 22284 26435 22336 26444
rect 22284 26401 22293 26435
rect 22293 26401 22327 26435
rect 22327 26401 22336 26435
rect 22284 26392 22336 26401
rect 22652 26392 22704 26444
rect 23296 26435 23348 26444
rect 23296 26401 23305 26435
rect 23305 26401 23339 26435
rect 23339 26401 23348 26435
rect 23296 26392 23348 26401
rect 25504 26392 25556 26444
rect 25872 26435 25924 26444
rect 25872 26401 25881 26435
rect 25881 26401 25915 26435
rect 25915 26401 25924 26435
rect 25872 26392 25924 26401
rect 26148 26435 26200 26444
rect 26148 26401 26157 26435
rect 26157 26401 26191 26435
rect 26191 26401 26200 26435
rect 26148 26392 26200 26401
rect 28448 26435 28500 26444
rect 28448 26401 28457 26435
rect 28457 26401 28491 26435
rect 28491 26401 28500 26435
rect 28448 26392 28500 26401
rect 29000 26392 29052 26444
rect 30104 26392 30156 26444
rect 31024 26392 31076 26444
rect 22192 26367 22244 26376
rect 22192 26333 22201 26367
rect 22201 26333 22235 26367
rect 22235 26333 22244 26367
rect 22192 26324 22244 26333
rect 23848 26324 23900 26376
rect 33232 26392 33284 26444
rect 33876 26392 33928 26444
rect 33692 26324 33744 26376
rect 2780 26256 2832 26308
rect 6000 26256 6052 26308
rect 7656 26256 7708 26308
rect 10692 26256 10744 26308
rect 2228 26188 2280 26240
rect 4620 26188 4672 26240
rect 6828 26231 6880 26240
rect 6828 26197 6837 26231
rect 6837 26197 6871 26231
rect 6871 26197 6880 26231
rect 6828 26188 6880 26197
rect 10416 26188 10468 26240
rect 10876 26188 10928 26240
rect 11060 26256 11112 26308
rect 12348 26256 12400 26308
rect 13544 26256 13596 26308
rect 17408 26299 17460 26308
rect 17408 26265 17417 26299
rect 17417 26265 17451 26299
rect 17451 26265 17460 26299
rect 17408 26256 17460 26265
rect 12072 26231 12124 26240
rect 12072 26197 12081 26231
rect 12081 26197 12115 26231
rect 12115 26197 12124 26231
rect 12072 26188 12124 26197
rect 14096 26231 14148 26240
rect 14096 26197 14105 26231
rect 14105 26197 14139 26231
rect 14139 26197 14148 26231
rect 14096 26188 14148 26197
rect 14464 26231 14516 26240
rect 14464 26197 14473 26231
rect 14473 26197 14507 26231
rect 14507 26197 14516 26231
rect 14464 26188 14516 26197
rect 18328 26188 18380 26240
rect 19248 26256 19300 26308
rect 20720 26256 20772 26308
rect 26700 26299 26752 26308
rect 26700 26265 26709 26299
rect 26709 26265 26743 26299
rect 26743 26265 26752 26299
rect 26700 26256 26752 26265
rect 27436 26256 27488 26308
rect 30012 26299 30064 26308
rect 30012 26265 30021 26299
rect 30021 26265 30055 26299
rect 30055 26265 30064 26299
rect 30012 26256 30064 26265
rect 32128 26256 32180 26308
rect 30380 26188 30432 26240
rect 32404 26188 32456 26240
rect 33416 26231 33468 26240
rect 33416 26197 33425 26231
rect 33425 26197 33459 26231
rect 33459 26197 33468 26231
rect 33416 26188 33468 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 3700 26027 3752 26036
rect 3700 25993 3709 26027
rect 3709 25993 3743 26027
rect 3743 25993 3752 26027
rect 3700 25984 3752 25993
rect 4712 26027 4764 26036
rect 4712 25993 4721 26027
rect 4721 25993 4755 26027
rect 4755 25993 4764 26027
rect 4712 25984 4764 25993
rect 9680 26027 9732 26036
rect 9680 25993 9689 26027
rect 9689 25993 9723 26027
rect 9723 25993 9732 26027
rect 9680 25984 9732 25993
rect 10140 25984 10192 26036
rect 14464 25984 14516 26036
rect 17040 26027 17092 26036
rect 17040 25993 17049 26027
rect 17049 25993 17083 26027
rect 17083 25993 17092 26027
rect 17040 25984 17092 25993
rect 17408 26027 17460 26036
rect 17408 25993 17417 26027
rect 17417 25993 17451 26027
rect 17451 25993 17460 26027
rect 17408 25984 17460 25993
rect 2688 25916 2740 25968
rect 2780 25780 2832 25832
rect 3792 25848 3844 25900
rect 7656 25916 7708 25968
rect 6460 25848 6512 25900
rect 7012 25848 7064 25900
rect 8208 25916 8260 25968
rect 8668 25916 8720 25968
rect 10784 25916 10836 25968
rect 13544 25916 13596 25968
rect 4068 25780 4120 25832
rect 5724 25780 5776 25832
rect 6736 25823 6788 25832
rect 6736 25789 6745 25823
rect 6745 25789 6779 25823
rect 6779 25789 6788 25823
rect 6736 25780 6788 25789
rect 6460 25712 6512 25764
rect 9220 25780 9272 25832
rect 9496 25780 9548 25832
rect 10048 25823 10100 25832
rect 10048 25789 10057 25823
rect 10057 25789 10091 25823
rect 10091 25789 10100 25823
rect 10048 25780 10100 25789
rect 10508 25712 10560 25764
rect 10876 25780 10928 25832
rect 5816 25644 5868 25696
rect 10048 25644 10100 25696
rect 12072 25848 12124 25900
rect 12808 25891 12860 25900
rect 12808 25857 12817 25891
rect 12817 25857 12851 25891
rect 12851 25857 12860 25891
rect 12808 25848 12860 25857
rect 18880 25984 18932 26036
rect 17960 25959 18012 25968
rect 17960 25925 17969 25959
rect 17969 25925 18003 25959
rect 18003 25925 18012 25959
rect 17960 25916 18012 25925
rect 19248 25916 19300 25968
rect 24952 25984 25004 26036
rect 26148 25984 26200 26036
rect 25780 25959 25832 25968
rect 25780 25925 25789 25959
rect 25789 25925 25823 25959
rect 25823 25925 25832 25959
rect 25780 25916 25832 25925
rect 20352 25848 20404 25900
rect 26516 25916 26568 25968
rect 14096 25780 14148 25832
rect 16856 25823 16908 25832
rect 16856 25789 16865 25823
rect 16865 25789 16899 25823
rect 16899 25789 16908 25823
rect 16856 25780 16908 25789
rect 16948 25823 17000 25832
rect 16948 25789 16957 25823
rect 16957 25789 16991 25823
rect 16991 25789 17000 25823
rect 16948 25780 17000 25789
rect 18512 25780 18564 25832
rect 28080 25891 28132 25900
rect 28080 25857 28089 25891
rect 28089 25857 28123 25891
rect 28123 25857 28132 25891
rect 28080 25848 28132 25857
rect 28264 25891 28316 25900
rect 28264 25857 28273 25891
rect 28273 25857 28307 25891
rect 28307 25857 28316 25891
rect 28264 25848 28316 25857
rect 31484 25984 31536 26036
rect 33692 25984 33744 26036
rect 30012 25916 30064 25968
rect 30380 25916 30432 25968
rect 32404 25959 32456 25968
rect 32404 25925 32413 25959
rect 32413 25925 32447 25959
rect 32447 25925 32456 25959
rect 32404 25916 32456 25925
rect 25136 25712 25188 25764
rect 25504 25823 25556 25832
rect 25504 25789 25513 25823
rect 25513 25789 25547 25823
rect 25547 25789 25556 25823
rect 25504 25780 25556 25789
rect 26240 25780 26292 25832
rect 26700 25780 26752 25832
rect 27804 25780 27856 25832
rect 28356 25823 28408 25832
rect 28356 25789 28365 25823
rect 28365 25789 28399 25823
rect 28399 25789 28408 25823
rect 28356 25780 28408 25789
rect 25964 25712 26016 25764
rect 19432 25687 19484 25696
rect 19432 25653 19441 25687
rect 19441 25653 19475 25687
rect 19475 25653 19484 25687
rect 19432 25644 19484 25653
rect 20996 25644 21048 25696
rect 29644 25891 29696 25900
rect 29644 25857 29653 25891
rect 29653 25857 29687 25891
rect 29687 25857 29696 25891
rect 29644 25848 29696 25857
rect 33508 25848 33560 25900
rect 34060 25848 34112 25900
rect 29552 25780 29604 25832
rect 30196 25823 30248 25832
rect 30196 25789 30205 25823
rect 30205 25789 30239 25823
rect 30239 25789 30248 25823
rect 30196 25780 30248 25789
rect 31116 25780 31168 25832
rect 32128 25823 32180 25832
rect 32128 25789 32137 25823
rect 32137 25789 32171 25823
rect 32171 25789 32180 25823
rect 32128 25780 32180 25789
rect 30656 25644 30708 25696
rect 31760 25644 31812 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 848 25372 900 25424
rect 2228 25347 2280 25356
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 2228 25313 2237 25347
rect 2237 25313 2271 25347
rect 2271 25313 2280 25347
rect 2228 25304 2280 25313
rect 2136 25279 2188 25288
rect 2136 25245 2145 25279
rect 2145 25245 2179 25279
rect 2179 25245 2188 25279
rect 2136 25236 2188 25245
rect 2780 25440 2832 25492
rect 3516 25440 3568 25492
rect 5356 25440 5408 25492
rect 5908 25483 5960 25492
rect 5908 25449 5917 25483
rect 5917 25449 5951 25483
rect 5951 25449 5960 25483
rect 5908 25440 5960 25449
rect 6368 25440 6420 25492
rect 2688 25372 2740 25424
rect 6736 25440 6788 25492
rect 10140 25483 10192 25492
rect 10140 25449 10149 25483
rect 10149 25449 10183 25483
rect 10183 25449 10192 25483
rect 10140 25440 10192 25449
rect 10508 25440 10560 25492
rect 10692 25440 10744 25492
rect 16948 25440 17000 25492
rect 18788 25440 18840 25492
rect 2780 25347 2832 25356
rect 2780 25313 2789 25347
rect 2789 25313 2823 25347
rect 2823 25313 2832 25347
rect 2780 25304 2832 25313
rect 3148 25304 3200 25356
rect 3792 25347 3844 25356
rect 3792 25313 3801 25347
rect 3801 25313 3835 25347
rect 3835 25313 3844 25347
rect 3792 25304 3844 25313
rect 6828 25372 6880 25424
rect 6092 25304 6144 25356
rect 14464 25372 14516 25424
rect 10232 25347 10284 25356
rect 10232 25313 10241 25347
rect 10241 25313 10275 25347
rect 10275 25313 10284 25347
rect 10232 25304 10284 25313
rect 14740 25347 14792 25356
rect 14740 25313 14749 25347
rect 14749 25313 14783 25347
rect 14783 25313 14792 25347
rect 14740 25304 14792 25313
rect 17224 25347 17276 25356
rect 17224 25313 17233 25347
rect 17233 25313 17267 25347
rect 17267 25313 17276 25347
rect 17224 25304 17276 25313
rect 5724 25279 5776 25288
rect 5724 25245 5733 25279
rect 5733 25245 5767 25279
rect 5767 25245 5776 25279
rect 5724 25236 5776 25245
rect 5908 25279 5960 25288
rect 5908 25245 5917 25279
rect 5917 25245 5951 25279
rect 5951 25245 5960 25279
rect 5908 25236 5960 25245
rect 6368 25279 6420 25288
rect 6368 25245 6377 25279
rect 6377 25245 6411 25279
rect 6411 25245 6420 25279
rect 6368 25236 6420 25245
rect 6552 25236 6604 25288
rect 6736 25236 6788 25288
rect 4344 25168 4396 25220
rect 4528 25168 4580 25220
rect 5448 25168 5500 25220
rect 1860 25100 1912 25152
rect 3332 25100 3384 25152
rect 6920 25168 6972 25220
rect 10048 25279 10100 25288
rect 10048 25245 10057 25279
rect 10057 25245 10091 25279
rect 10091 25245 10100 25279
rect 10048 25236 10100 25245
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 14464 25236 14516 25288
rect 14924 25279 14976 25288
rect 14924 25245 14933 25279
rect 14933 25245 14967 25279
rect 14967 25245 14976 25279
rect 14924 25236 14976 25245
rect 19248 25236 19300 25288
rect 20444 25236 20496 25288
rect 22284 25304 22336 25356
rect 21824 25279 21876 25288
rect 21824 25245 21833 25279
rect 21833 25245 21867 25279
rect 21867 25245 21876 25279
rect 21824 25236 21876 25245
rect 22836 25236 22888 25288
rect 24952 25347 25004 25356
rect 24952 25313 24961 25347
rect 24961 25313 24995 25347
rect 24995 25313 25004 25347
rect 24952 25304 25004 25313
rect 29644 25304 29696 25356
rect 30564 25304 30616 25356
rect 23388 25236 23440 25288
rect 27436 25236 27488 25288
rect 9956 25168 10008 25220
rect 10232 25100 10284 25152
rect 10600 25211 10652 25220
rect 10600 25177 10625 25211
rect 10625 25177 10652 25211
rect 10600 25168 10652 25177
rect 13820 25168 13872 25220
rect 15200 25211 15252 25220
rect 15200 25177 15209 25211
rect 15209 25177 15243 25211
rect 15243 25177 15252 25211
rect 15200 25168 15252 25177
rect 15844 25168 15896 25220
rect 18512 25168 18564 25220
rect 20352 25168 20404 25220
rect 20812 25168 20864 25220
rect 22100 25168 22152 25220
rect 25228 25211 25280 25220
rect 25228 25177 25237 25211
rect 25237 25177 25271 25211
rect 25271 25177 25280 25211
rect 25228 25168 25280 25177
rect 26608 25168 26660 25220
rect 30196 25236 30248 25288
rect 32128 25236 32180 25288
rect 33416 25304 33468 25356
rect 34428 25304 34480 25356
rect 33784 25279 33836 25288
rect 33784 25245 33793 25279
rect 33793 25245 33827 25279
rect 33827 25245 33836 25279
rect 33784 25236 33836 25245
rect 14004 25100 14056 25152
rect 27436 25100 27488 25152
rect 30472 25168 30524 25220
rect 31392 25168 31444 25220
rect 33324 25211 33376 25220
rect 33324 25177 33333 25211
rect 33333 25177 33367 25211
rect 33367 25177 33376 25211
rect 33324 25168 33376 25177
rect 34520 25168 34572 25220
rect 35440 25100 35492 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 1584 24896 1636 24948
rect 2136 24896 2188 24948
rect 2688 24896 2740 24948
rect 2964 24828 3016 24880
rect 3148 24803 3200 24812
rect 3148 24769 3157 24803
rect 3157 24769 3191 24803
rect 3191 24769 3200 24803
rect 3148 24760 3200 24769
rect 4344 24939 4396 24948
rect 4344 24905 4353 24939
rect 4353 24905 4387 24939
rect 4387 24905 4396 24939
rect 4344 24896 4396 24905
rect 5724 24896 5776 24948
rect 6092 24896 6144 24948
rect 14004 24939 14056 24948
rect 14004 24905 14013 24939
rect 14013 24905 14047 24939
rect 14047 24905 14056 24939
rect 14004 24896 14056 24905
rect 15200 24896 15252 24948
rect 16948 24896 17000 24948
rect 3332 24692 3384 24744
rect 4528 24828 4580 24880
rect 4160 24803 4212 24812
rect 4160 24769 4169 24803
rect 4169 24769 4203 24803
rect 4203 24769 4212 24803
rect 4160 24760 4212 24769
rect 4804 24803 4856 24812
rect 4804 24769 4813 24803
rect 4813 24769 4847 24803
rect 4847 24769 4856 24803
rect 5448 24828 5500 24880
rect 6368 24828 6420 24880
rect 4804 24760 4856 24769
rect 5356 24803 5408 24812
rect 5356 24769 5365 24803
rect 5365 24769 5399 24803
rect 5399 24769 5408 24803
rect 5356 24760 5408 24769
rect 5908 24760 5960 24812
rect 6736 24760 6788 24812
rect 7012 24828 7064 24880
rect 8668 24828 8720 24880
rect 19248 24828 19300 24880
rect 11060 24760 11112 24812
rect 13912 24803 13964 24812
rect 13912 24769 13921 24803
rect 13921 24769 13955 24803
rect 13955 24769 13964 24803
rect 13912 24760 13964 24769
rect 18512 24803 18564 24812
rect 18512 24769 18521 24803
rect 18521 24769 18555 24803
rect 18555 24769 18564 24803
rect 18512 24760 18564 24769
rect 20444 24760 20496 24812
rect 22928 24896 22980 24948
rect 28356 24896 28408 24948
rect 28724 24896 28776 24948
rect 34428 24939 34480 24948
rect 34428 24905 34437 24939
rect 34437 24905 34471 24939
rect 34471 24905 34480 24939
rect 34428 24896 34480 24905
rect 22100 24871 22152 24880
rect 22100 24837 22109 24871
rect 22109 24837 22143 24871
rect 22143 24837 22152 24871
rect 22100 24828 22152 24837
rect 22560 24828 22612 24880
rect 20996 24803 21048 24812
rect 20996 24769 21005 24803
rect 21005 24769 21039 24803
rect 21039 24769 21048 24803
rect 20996 24760 21048 24769
rect 25504 24828 25556 24880
rect 7104 24735 7156 24744
rect 7104 24701 7113 24735
rect 7113 24701 7147 24735
rect 7147 24701 7156 24735
rect 7104 24692 7156 24701
rect 8300 24692 8352 24744
rect 13820 24692 13872 24744
rect 14740 24692 14792 24744
rect 16120 24735 16172 24744
rect 16120 24701 16129 24735
rect 16129 24701 16163 24735
rect 16163 24701 16172 24735
rect 16120 24692 16172 24701
rect 16304 24735 16356 24744
rect 16304 24701 16313 24735
rect 16313 24701 16347 24735
rect 16347 24701 16356 24735
rect 16304 24692 16356 24701
rect 16856 24692 16908 24744
rect 5724 24624 5776 24676
rect 19892 24624 19944 24676
rect 3056 24556 3108 24608
rect 3700 24599 3752 24608
rect 3700 24565 3709 24599
rect 3709 24565 3743 24599
rect 3743 24565 3752 24599
rect 3700 24556 3752 24565
rect 6552 24556 6604 24608
rect 6736 24556 6788 24608
rect 13084 24556 13136 24608
rect 20352 24556 20404 24608
rect 22560 24692 22612 24744
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 27528 24828 27580 24880
rect 29552 24828 29604 24880
rect 33508 24828 33560 24880
rect 30380 24760 30432 24812
rect 31208 24803 31260 24812
rect 31208 24769 31217 24803
rect 31217 24769 31251 24803
rect 31251 24769 31260 24803
rect 31208 24760 31260 24769
rect 23388 24692 23440 24744
rect 23664 24735 23716 24744
rect 23664 24701 23673 24735
rect 23673 24701 23707 24735
rect 23707 24701 23716 24735
rect 23664 24692 23716 24701
rect 23940 24735 23992 24744
rect 23940 24701 23949 24735
rect 23949 24701 23983 24735
rect 23983 24701 23992 24735
rect 23940 24692 23992 24701
rect 25044 24624 25096 24676
rect 23204 24556 23256 24608
rect 26056 24735 26108 24744
rect 26056 24701 26065 24735
rect 26065 24701 26099 24735
rect 26099 24701 26108 24735
rect 26056 24692 26108 24701
rect 26240 24692 26292 24744
rect 27804 24692 27856 24744
rect 29368 24692 29420 24744
rect 28632 24556 28684 24608
rect 32036 24692 32088 24744
rect 32128 24692 32180 24744
rect 33324 24692 33376 24744
rect 30840 24599 30892 24608
rect 30840 24565 30849 24599
rect 30849 24565 30883 24599
rect 30883 24565 30892 24599
rect 30840 24556 30892 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 7104 24352 7156 24404
rect 13912 24395 13964 24404
rect 13912 24361 13921 24395
rect 13921 24361 13955 24395
rect 13955 24361 13964 24395
rect 13912 24352 13964 24361
rect 16120 24352 16172 24404
rect 22284 24395 22336 24404
rect 22284 24361 22293 24395
rect 22293 24361 22327 24395
rect 22327 24361 22336 24395
rect 22284 24352 22336 24361
rect 25872 24352 25924 24404
rect 28264 24352 28316 24404
rect 31208 24352 31260 24404
rect 3148 24216 3200 24268
rect 4068 24216 4120 24268
rect 2964 24148 3016 24200
rect 6920 24148 6972 24200
rect 1860 24123 1912 24132
rect 1860 24089 1869 24123
rect 1869 24089 1903 24123
rect 1903 24089 1912 24123
rect 1860 24080 1912 24089
rect 6736 24080 6788 24132
rect 11796 24216 11848 24268
rect 12164 24259 12216 24268
rect 12164 24225 12173 24259
rect 12173 24225 12207 24259
rect 12207 24225 12216 24259
rect 12164 24216 12216 24225
rect 13084 24216 13136 24268
rect 18512 24216 18564 24268
rect 7748 24191 7800 24200
rect 7748 24157 7757 24191
rect 7757 24157 7791 24191
rect 7791 24157 7800 24191
rect 7748 24148 7800 24157
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 15844 24148 15896 24200
rect 20444 24284 20496 24336
rect 31116 24284 31168 24336
rect 20352 24216 20404 24268
rect 20812 24259 20864 24268
rect 20812 24225 20821 24259
rect 20821 24225 20855 24259
rect 20855 24225 20864 24259
rect 20812 24216 20864 24225
rect 23664 24216 23716 24268
rect 25044 24216 25096 24268
rect 28632 24259 28684 24268
rect 28632 24225 28641 24259
rect 28641 24225 28675 24259
rect 28675 24225 28684 24259
rect 28632 24216 28684 24225
rect 29368 24259 29420 24268
rect 29368 24225 29377 24259
rect 29377 24225 29411 24259
rect 29411 24225 29420 24259
rect 29368 24216 29420 24225
rect 30840 24216 30892 24268
rect 34520 24395 34572 24404
rect 34520 24361 34529 24395
rect 34529 24361 34563 24395
rect 34563 24361 34572 24395
rect 34520 24352 34572 24361
rect 32036 24259 32088 24268
rect 32036 24225 32045 24259
rect 32045 24225 32079 24259
rect 32079 24225 32088 24259
rect 32036 24216 32088 24225
rect 32128 24216 32180 24268
rect 19892 24191 19944 24200
rect 19892 24157 19901 24191
rect 19901 24157 19935 24191
rect 19935 24157 19944 24191
rect 19892 24148 19944 24157
rect 20076 24148 20128 24200
rect 22560 24148 22612 24200
rect 13820 24080 13872 24132
rect 14740 24123 14792 24132
rect 14740 24089 14749 24123
rect 14749 24089 14783 24123
rect 14783 24089 14792 24123
rect 14740 24080 14792 24089
rect 17776 24080 17828 24132
rect 24124 24123 24176 24132
rect 24124 24089 24133 24123
rect 24133 24089 24167 24123
rect 24167 24089 24176 24123
rect 24124 24080 24176 24089
rect 26240 24191 26292 24200
rect 26240 24157 26249 24191
rect 26249 24157 26283 24191
rect 26283 24157 26292 24191
rect 26240 24148 26292 24157
rect 27528 24148 27580 24200
rect 16396 24055 16448 24064
rect 16396 24021 16405 24055
rect 16405 24021 16439 24055
rect 16439 24021 16448 24055
rect 16396 24012 16448 24021
rect 19984 24012 20036 24064
rect 22928 24012 22980 24064
rect 26516 24123 26568 24132
rect 26516 24089 26525 24123
rect 26525 24089 26559 24123
rect 26559 24089 26568 24123
rect 26516 24080 26568 24089
rect 28724 24191 28776 24200
rect 28724 24157 28733 24191
rect 28733 24157 28767 24191
rect 28767 24157 28776 24191
rect 28724 24148 28776 24157
rect 28908 24191 28960 24200
rect 28908 24157 28917 24191
rect 28917 24157 28951 24191
rect 28951 24157 28960 24191
rect 28908 24148 28960 24157
rect 29552 24191 29604 24200
rect 29552 24157 29561 24191
rect 29561 24157 29595 24191
rect 29595 24157 29604 24191
rect 29552 24148 29604 24157
rect 31760 24191 31812 24200
rect 31760 24157 31769 24191
rect 31769 24157 31803 24191
rect 31803 24157 31812 24191
rect 31760 24148 31812 24157
rect 30380 24080 30432 24132
rect 33048 24123 33100 24132
rect 33048 24089 33057 24123
rect 33057 24089 33091 24123
rect 33091 24089 33100 24123
rect 33048 24080 33100 24089
rect 33508 24080 33560 24132
rect 33232 24012 33284 24064
rect 34060 24012 34112 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 3700 23740 3752 23792
rect 5632 23808 5684 23860
rect 7748 23808 7800 23860
rect 5080 23740 5132 23792
rect 5356 23740 5408 23792
rect 848 23672 900 23724
rect 2136 23672 2188 23724
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 6920 23672 6972 23724
rect 8024 23672 8076 23724
rect 8576 23672 8628 23724
rect 8760 23715 8812 23724
rect 8760 23681 8769 23715
rect 8769 23681 8803 23715
rect 8803 23681 8812 23715
rect 9220 23740 9272 23792
rect 9496 23851 9548 23860
rect 9496 23817 9505 23851
rect 9505 23817 9539 23851
rect 9539 23817 9548 23851
rect 9496 23808 9548 23817
rect 10140 23851 10192 23860
rect 10140 23817 10149 23851
rect 10149 23817 10183 23851
rect 10183 23817 10192 23851
rect 10140 23808 10192 23817
rect 10692 23808 10744 23860
rect 13912 23808 13964 23860
rect 14740 23808 14792 23860
rect 16120 23808 16172 23860
rect 17776 23851 17828 23860
rect 17776 23817 17785 23851
rect 17785 23817 17819 23851
rect 17819 23817 17828 23851
rect 17776 23808 17828 23817
rect 18696 23808 18748 23860
rect 20076 23808 20128 23860
rect 25228 23808 25280 23860
rect 25872 23808 25924 23860
rect 26516 23808 26568 23860
rect 28264 23808 28316 23860
rect 33048 23808 33100 23860
rect 34520 23808 34572 23860
rect 10232 23783 10284 23792
rect 10232 23749 10241 23783
rect 10241 23749 10275 23783
rect 10275 23749 10284 23783
rect 10232 23740 10284 23749
rect 8760 23672 8812 23681
rect 9772 23672 9824 23724
rect 16396 23740 16448 23792
rect 19248 23740 19300 23792
rect 19984 23783 20036 23792
rect 19984 23749 19993 23783
rect 19993 23749 20027 23783
rect 20027 23749 20036 23783
rect 19984 23740 20036 23749
rect 23940 23783 23992 23792
rect 23940 23749 23949 23783
rect 23949 23749 23983 23783
rect 23983 23749 23992 23783
rect 23940 23740 23992 23749
rect 27436 23783 27488 23792
rect 27436 23749 27445 23783
rect 27445 23749 27479 23783
rect 27479 23749 27488 23783
rect 27436 23740 27488 23749
rect 30472 23740 30524 23792
rect 10508 23672 10560 23724
rect 13912 23672 13964 23724
rect 10876 23604 10928 23656
rect 15384 23604 15436 23656
rect 16304 23604 16356 23656
rect 17132 23647 17184 23656
rect 17132 23613 17141 23647
rect 17141 23613 17175 23647
rect 17175 23613 17184 23647
rect 17132 23604 17184 23613
rect 17316 23647 17368 23656
rect 17316 23613 17325 23647
rect 17325 23613 17359 23647
rect 17359 23613 17368 23647
rect 17316 23604 17368 23613
rect 19616 23604 19668 23656
rect 20352 23672 20404 23724
rect 23204 23715 23256 23724
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 23388 23672 23440 23724
rect 23480 23715 23532 23724
rect 23480 23681 23489 23715
rect 23489 23681 23523 23715
rect 23523 23681 23532 23715
rect 23480 23672 23532 23681
rect 24124 23672 24176 23724
rect 26516 23672 26568 23724
rect 30564 23715 30616 23724
rect 30564 23681 30573 23715
rect 30573 23681 30607 23715
rect 30607 23681 30616 23715
rect 30564 23672 30616 23681
rect 30748 23715 30800 23724
rect 30748 23681 30757 23715
rect 30757 23681 30791 23715
rect 30791 23681 30800 23715
rect 30748 23672 30800 23681
rect 31760 23740 31812 23792
rect 23756 23604 23808 23656
rect 5816 23536 5868 23588
rect 26056 23604 26108 23656
rect 27528 23647 27580 23656
rect 27528 23613 27537 23647
rect 27537 23613 27571 23647
rect 27571 23613 27580 23647
rect 27528 23604 27580 23613
rect 30196 23604 30248 23656
rect 30656 23604 30708 23656
rect 32404 23604 32456 23656
rect 33876 23715 33928 23724
rect 33876 23681 33885 23715
rect 33885 23681 33919 23715
rect 33919 23681 33928 23715
rect 33876 23672 33928 23681
rect 34060 23672 34112 23724
rect 33232 23647 33284 23656
rect 33232 23613 33241 23647
rect 33241 23613 33275 23647
rect 33275 23613 33284 23647
rect 33232 23604 33284 23613
rect 34428 23604 34480 23656
rect 27620 23536 27672 23588
rect 28080 23536 28132 23588
rect 28908 23536 28960 23588
rect 5264 23468 5316 23520
rect 5540 23468 5592 23520
rect 6184 23468 6236 23520
rect 8668 23468 8720 23520
rect 9128 23468 9180 23520
rect 9680 23511 9732 23520
rect 9680 23477 9689 23511
rect 9689 23477 9723 23511
rect 9723 23477 9732 23511
rect 9680 23468 9732 23477
rect 10416 23511 10468 23520
rect 10416 23477 10425 23511
rect 10425 23477 10459 23511
rect 10459 23477 10468 23511
rect 10416 23468 10468 23477
rect 10600 23511 10652 23520
rect 10600 23477 10609 23511
rect 10609 23477 10643 23511
rect 10643 23477 10652 23511
rect 10600 23468 10652 23477
rect 12440 23468 12492 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 5080 23264 5132 23316
rect 6368 23264 6420 23316
rect 8760 23307 8812 23316
rect 8760 23273 8769 23307
rect 8769 23273 8803 23307
rect 8803 23273 8812 23307
rect 8760 23264 8812 23273
rect 9220 23264 9272 23316
rect 9680 23264 9732 23316
rect 10416 23264 10468 23316
rect 13912 23307 13964 23316
rect 13912 23273 13921 23307
rect 13921 23273 13955 23307
rect 13955 23273 13964 23307
rect 13912 23264 13964 23273
rect 9496 23196 9548 23248
rect 9772 23196 9824 23248
rect 3148 23128 3200 23180
rect 5264 23171 5316 23180
rect 5264 23137 5273 23171
rect 5273 23137 5307 23171
rect 5307 23137 5316 23171
rect 5264 23128 5316 23137
rect 10324 23171 10376 23180
rect 10324 23137 10333 23171
rect 10333 23137 10367 23171
rect 10367 23137 10376 23171
rect 10324 23128 10376 23137
rect 12164 23171 12216 23180
rect 12164 23137 12173 23171
rect 12173 23137 12207 23171
rect 12207 23137 12216 23171
rect 12164 23128 12216 23137
rect 12440 23171 12492 23180
rect 12440 23137 12449 23171
rect 12449 23137 12483 23171
rect 12483 23137 12492 23171
rect 12440 23128 12492 23137
rect 14648 23171 14700 23180
rect 14648 23137 14657 23171
rect 14657 23137 14691 23171
rect 14691 23137 14700 23171
rect 14648 23128 14700 23137
rect 2780 23103 2832 23112
rect 2780 23069 2789 23103
rect 2789 23069 2823 23103
rect 2823 23069 2832 23103
rect 2780 23060 2832 23069
rect 3700 23060 3752 23112
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 4068 23060 4120 23112
rect 4804 22992 4856 23044
rect 8300 23060 8352 23112
rect 5540 22992 5592 23044
rect 2688 22924 2740 22976
rect 3424 22924 3476 22976
rect 5264 22924 5316 22976
rect 7288 23035 7340 23044
rect 7288 23001 7297 23035
rect 7297 23001 7331 23035
rect 7331 23001 7340 23035
rect 7288 22992 7340 23001
rect 9128 23060 9180 23112
rect 9496 23035 9548 23044
rect 9496 23001 9505 23035
rect 9505 23001 9539 23035
rect 9539 23001 9548 23035
rect 9496 22992 9548 23001
rect 9680 23103 9732 23112
rect 9680 23069 9689 23103
rect 9689 23069 9723 23103
rect 9723 23069 9732 23103
rect 9680 23060 9732 23069
rect 9772 23103 9824 23112
rect 9772 23069 9781 23103
rect 9781 23069 9815 23103
rect 9815 23069 9824 23103
rect 9772 23060 9824 23069
rect 9864 23103 9916 23112
rect 9864 23069 9873 23103
rect 9873 23069 9907 23103
rect 9907 23069 9916 23103
rect 9864 23060 9916 23069
rect 15292 23103 15344 23112
rect 15292 23069 15301 23103
rect 15301 23069 15335 23103
rect 15335 23069 15344 23103
rect 15292 23060 15344 23069
rect 23480 23264 23532 23316
rect 30656 23264 30708 23316
rect 34428 23307 34480 23316
rect 34428 23273 34437 23307
rect 34437 23273 34471 23307
rect 34471 23273 34480 23307
rect 34428 23264 34480 23273
rect 18696 23103 18748 23112
rect 18696 23069 18705 23103
rect 18705 23069 18739 23103
rect 18739 23069 18748 23103
rect 18696 23060 18748 23069
rect 27528 23196 27580 23248
rect 21364 23128 21416 23180
rect 10048 22992 10100 23044
rect 11060 22992 11112 23044
rect 13820 22992 13872 23044
rect 10876 22924 10928 22976
rect 14004 22924 14056 22976
rect 14556 22924 14608 22976
rect 15568 23035 15620 23044
rect 15568 23001 15577 23035
rect 15577 23001 15611 23035
rect 15611 23001 15620 23035
rect 15568 22992 15620 23001
rect 16856 22992 16908 23044
rect 15844 22924 15896 22976
rect 17040 22967 17092 22976
rect 17040 22933 17049 22967
rect 17049 22933 17083 22967
rect 17083 22933 17092 22967
rect 17040 22924 17092 22933
rect 18052 23035 18104 23044
rect 18052 23001 18061 23035
rect 18061 23001 18095 23035
rect 18095 23001 18104 23035
rect 18052 22992 18104 23001
rect 19984 23035 20036 23044
rect 19984 23001 19993 23035
rect 19993 23001 20027 23035
rect 20027 23001 20036 23035
rect 19984 22992 20036 23001
rect 20536 23060 20588 23112
rect 22928 23171 22980 23180
rect 22928 23137 22937 23171
rect 22937 23137 22971 23171
rect 22971 23137 22980 23171
rect 22928 23128 22980 23137
rect 23664 23128 23716 23180
rect 26240 23128 26292 23180
rect 26976 23128 27028 23180
rect 30196 23171 30248 23180
rect 30196 23137 30205 23171
rect 30205 23137 30239 23171
rect 30239 23137 30248 23171
rect 30196 23128 30248 23137
rect 32128 23128 32180 23180
rect 21180 23035 21232 23044
rect 21180 23001 21189 23035
rect 21189 23001 21223 23035
rect 21223 23001 21232 23035
rect 21180 22992 21232 23001
rect 22468 23060 22520 23112
rect 27620 23060 27672 23112
rect 28632 23103 28684 23112
rect 18144 22924 18196 22976
rect 22192 22924 22244 22976
rect 23572 22992 23624 23044
rect 23940 22924 23992 22976
rect 26148 22992 26200 23044
rect 27252 22992 27304 23044
rect 26240 22924 26292 22976
rect 26884 22924 26936 22976
rect 28632 23069 28641 23103
rect 28641 23069 28675 23103
rect 28675 23069 28684 23103
rect 28632 23060 28684 23069
rect 29000 23060 29052 23112
rect 29552 23060 29604 23112
rect 33232 22992 33284 23044
rect 27896 22924 27948 22976
rect 29368 22924 29420 22976
rect 31484 22924 31536 22976
rect 33416 22992 33468 23044
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 1124 22720 1176 22772
rect 2688 22695 2740 22704
rect 2688 22661 2697 22695
rect 2697 22661 2731 22695
rect 2731 22661 2740 22695
rect 2688 22652 2740 22661
rect 3424 22695 3476 22704
rect 3424 22661 3433 22695
rect 3433 22661 3467 22695
rect 3467 22661 3476 22695
rect 3424 22652 3476 22661
rect 3700 22652 3752 22704
rect 4804 22652 4856 22704
rect 5540 22695 5592 22704
rect 5540 22661 5549 22695
rect 5549 22661 5583 22695
rect 5583 22661 5592 22695
rect 5540 22652 5592 22661
rect 5632 22652 5684 22704
rect 6276 22652 6328 22704
rect 7288 22720 7340 22772
rect 8576 22763 8628 22772
rect 8576 22729 8585 22763
rect 8585 22729 8619 22763
rect 8619 22729 8628 22763
rect 8576 22720 8628 22729
rect 8668 22763 8720 22772
rect 8668 22729 8677 22763
rect 8677 22729 8711 22763
rect 8711 22729 8720 22763
rect 8668 22720 8720 22729
rect 3148 22627 3200 22636
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 2780 22559 2832 22568
rect 2780 22525 2789 22559
rect 2789 22525 2823 22559
rect 2823 22525 2832 22559
rect 2780 22516 2832 22525
rect 4068 22516 4120 22568
rect 4804 22516 4856 22568
rect 5264 22516 5316 22568
rect 6920 22584 6972 22636
rect 9128 22652 9180 22704
rect 10048 22763 10100 22772
rect 10048 22729 10057 22763
rect 10057 22729 10091 22763
rect 10091 22729 10100 22763
rect 10048 22720 10100 22729
rect 10508 22763 10560 22772
rect 10508 22729 10517 22763
rect 10517 22729 10551 22763
rect 10551 22729 10560 22763
rect 10508 22720 10560 22729
rect 9404 22584 9456 22636
rect 5724 22491 5776 22500
rect 5724 22457 5733 22491
rect 5733 22457 5767 22491
rect 5767 22457 5776 22491
rect 5724 22448 5776 22457
rect 1676 22380 1728 22432
rect 4896 22423 4948 22432
rect 4896 22389 4905 22423
rect 4905 22389 4939 22423
rect 4939 22389 4948 22423
rect 4896 22380 4948 22389
rect 5448 22380 5500 22432
rect 6552 22516 6604 22568
rect 10416 22584 10468 22636
rect 10508 22627 10560 22636
rect 10508 22593 10517 22627
rect 10517 22593 10551 22627
rect 10551 22593 10560 22627
rect 10508 22584 10560 22593
rect 10784 22652 10836 22704
rect 10692 22627 10744 22636
rect 10692 22593 10701 22627
rect 10701 22593 10735 22627
rect 10735 22593 10744 22627
rect 10692 22584 10744 22593
rect 10876 22627 10928 22636
rect 10876 22593 10885 22627
rect 10885 22593 10919 22627
rect 10919 22593 10928 22627
rect 10876 22584 10928 22593
rect 12164 22584 12216 22636
rect 14096 22720 14148 22772
rect 14464 22720 14516 22772
rect 15292 22720 15344 22772
rect 17316 22720 17368 22772
rect 19616 22720 19668 22772
rect 20628 22720 20680 22772
rect 13820 22652 13872 22704
rect 15844 22652 15896 22704
rect 16856 22652 16908 22704
rect 18052 22695 18104 22704
rect 18052 22661 18061 22695
rect 18061 22661 18095 22695
rect 18095 22661 18104 22695
rect 18052 22652 18104 22661
rect 18144 22652 18196 22704
rect 19984 22652 20036 22704
rect 14096 22627 14148 22636
rect 14096 22593 14105 22627
rect 14105 22593 14139 22627
rect 14139 22593 14148 22627
rect 14096 22584 14148 22593
rect 17040 22584 17092 22636
rect 19616 22627 19668 22636
rect 14004 22516 14056 22568
rect 14372 22559 14424 22568
rect 14372 22525 14381 22559
rect 14381 22525 14415 22559
rect 14415 22525 14424 22559
rect 14372 22516 14424 22525
rect 17132 22516 17184 22568
rect 19616 22593 19625 22627
rect 19625 22593 19659 22627
rect 19659 22593 19668 22627
rect 19616 22584 19668 22593
rect 23572 22720 23624 22772
rect 23940 22720 23992 22772
rect 27068 22720 27120 22772
rect 22192 22695 22244 22704
rect 22192 22661 22201 22695
rect 22201 22661 22235 22695
rect 22235 22661 22244 22695
rect 22192 22652 22244 22661
rect 22652 22652 22704 22704
rect 26148 22652 26200 22704
rect 27252 22695 27304 22704
rect 27252 22661 27261 22695
rect 27261 22661 27295 22695
rect 27295 22661 27304 22695
rect 27252 22652 27304 22661
rect 28632 22720 28684 22772
rect 30748 22763 30800 22772
rect 30748 22729 30757 22763
rect 30757 22729 30791 22763
rect 30791 22729 30800 22763
rect 30748 22720 30800 22729
rect 33876 22763 33928 22772
rect 33876 22729 33885 22763
rect 33885 22729 33919 22763
rect 33919 22729 33928 22763
rect 33876 22720 33928 22729
rect 31484 22652 31536 22704
rect 32404 22695 32456 22704
rect 32404 22661 32413 22695
rect 32413 22661 32447 22695
rect 32447 22661 32456 22695
rect 32404 22652 32456 22661
rect 33416 22652 33468 22704
rect 20536 22516 20588 22568
rect 23664 22584 23716 22636
rect 25412 22584 25464 22636
rect 25964 22627 26016 22636
rect 25964 22593 25973 22627
rect 25973 22593 26007 22627
rect 26007 22593 26016 22627
rect 25964 22584 26016 22593
rect 29000 22627 29052 22636
rect 29000 22593 29009 22627
rect 29009 22593 29043 22627
rect 29043 22593 29052 22627
rect 29000 22584 29052 22593
rect 32128 22627 32180 22636
rect 32128 22593 32137 22627
rect 32137 22593 32171 22627
rect 32171 22593 32180 22627
rect 32128 22584 32180 22593
rect 22560 22516 22612 22568
rect 24032 22559 24084 22568
rect 24032 22525 24041 22559
rect 24041 22525 24075 22559
rect 24075 22525 24084 22559
rect 24032 22516 24084 22525
rect 21364 22491 21416 22500
rect 21364 22457 21373 22491
rect 21373 22457 21407 22491
rect 21407 22457 21416 22491
rect 21364 22448 21416 22457
rect 25044 22448 25096 22500
rect 7288 22380 7340 22432
rect 7656 22423 7708 22432
rect 7656 22389 7665 22423
rect 7665 22389 7699 22423
rect 7699 22389 7708 22423
rect 7656 22380 7708 22389
rect 8208 22380 8260 22432
rect 8392 22380 8444 22432
rect 9772 22380 9824 22432
rect 10784 22380 10836 22432
rect 14556 22380 14608 22432
rect 15016 22380 15068 22432
rect 15844 22423 15896 22432
rect 15844 22389 15853 22423
rect 15853 22389 15887 22423
rect 15887 22389 15896 22423
rect 15844 22380 15896 22389
rect 16856 22423 16908 22432
rect 16856 22389 16865 22423
rect 16865 22389 16899 22423
rect 16899 22389 16908 22423
rect 16856 22380 16908 22389
rect 25504 22423 25556 22432
rect 25504 22389 25513 22423
rect 25513 22389 25547 22423
rect 25547 22389 25556 22423
rect 26148 22559 26200 22568
rect 26148 22525 26157 22559
rect 26157 22525 26191 22559
rect 26191 22525 26200 22559
rect 26148 22516 26200 22525
rect 26424 22516 26476 22568
rect 26976 22559 27028 22568
rect 26976 22525 26985 22559
rect 26985 22525 27019 22559
rect 27019 22525 27028 22559
rect 26976 22516 27028 22525
rect 29276 22559 29328 22568
rect 29276 22525 29285 22559
rect 29285 22525 29319 22559
rect 29319 22525 29328 22559
rect 29276 22516 29328 22525
rect 25504 22380 25556 22389
rect 27068 22380 27120 22432
rect 30012 22380 30064 22432
rect 30472 22380 30524 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1676 22219 1728 22228
rect 1676 22185 1706 22219
rect 1706 22185 1728 22219
rect 1676 22176 1728 22185
rect 3976 22176 4028 22228
rect 5448 22176 5500 22228
rect 2780 22108 2832 22160
rect 6276 22219 6328 22228
rect 6276 22185 6285 22219
rect 6285 22185 6319 22219
rect 6319 22185 6328 22219
rect 6276 22176 6328 22185
rect 10600 22176 10652 22228
rect 14372 22176 14424 22228
rect 15568 22219 15620 22228
rect 15568 22185 15577 22219
rect 15577 22185 15611 22219
rect 15611 22185 15620 22219
rect 15568 22176 15620 22185
rect 16856 22176 16908 22228
rect 21180 22176 21232 22228
rect 22468 22219 22520 22228
rect 22468 22185 22477 22219
rect 22477 22185 22511 22219
rect 22511 22185 22520 22219
rect 22468 22176 22520 22185
rect 25044 22176 25096 22228
rect 25964 22176 26016 22228
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 4896 22040 4948 22092
rect 9680 22108 9732 22160
rect 10508 22108 10560 22160
rect 5816 22040 5868 22092
rect 6828 22040 6880 22092
rect 7104 22040 7156 22092
rect 15016 22083 15068 22092
rect 15016 22049 15025 22083
rect 15025 22049 15059 22083
rect 15059 22049 15068 22083
rect 15016 22040 15068 22049
rect 15384 22108 15436 22160
rect 2964 21904 3016 21956
rect 3884 21904 3936 21956
rect 4344 21947 4396 21956
rect 4344 21913 4353 21947
rect 4353 21913 4387 21947
rect 4387 21913 4396 21947
rect 4344 21904 4396 21913
rect 4160 21836 4212 21888
rect 4712 21836 4764 21888
rect 6828 21904 6880 21956
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 8208 21972 8260 22024
rect 10048 21972 10100 22024
rect 15844 22040 15896 22092
rect 17224 22040 17276 22092
rect 20628 22040 20680 22092
rect 23664 22040 23716 22092
rect 25412 22040 25464 22092
rect 26240 22219 26292 22228
rect 26240 22185 26249 22219
rect 26249 22185 26283 22219
rect 26283 22185 26292 22219
rect 26240 22176 26292 22185
rect 27896 22219 27948 22228
rect 27896 22185 27926 22219
rect 27926 22185 27948 22219
rect 27896 22176 27948 22185
rect 29368 22219 29420 22228
rect 29368 22185 29377 22219
rect 29377 22185 29411 22219
rect 29411 22185 29420 22219
rect 29368 22176 29420 22185
rect 26424 22108 26476 22160
rect 15292 21972 15344 22024
rect 11060 21904 11112 21956
rect 16948 21904 17000 21956
rect 18144 21904 18196 21956
rect 22560 21904 22612 21956
rect 5540 21836 5592 21888
rect 6000 21836 6052 21888
rect 6184 21836 6236 21888
rect 6460 21879 6512 21888
rect 6460 21845 6469 21879
rect 6469 21845 6503 21879
rect 6503 21845 6512 21879
rect 6460 21836 6512 21845
rect 7104 21879 7156 21888
rect 7104 21845 7113 21879
rect 7113 21845 7147 21879
rect 7147 21845 7156 21879
rect 7104 21836 7156 21845
rect 23572 22015 23624 22024
rect 23572 21981 23581 22015
rect 23581 21981 23615 22015
rect 23615 21981 23624 22015
rect 23572 21972 23624 21981
rect 23756 22015 23808 22024
rect 23756 21981 23765 22015
rect 23765 21981 23799 22015
rect 23799 21981 23808 22015
rect 23756 21972 23808 21981
rect 24032 21972 24084 22024
rect 26976 22040 27028 22092
rect 29276 22040 29328 22092
rect 26884 21972 26936 22024
rect 30012 22015 30064 22024
rect 30012 21981 30021 22015
rect 30021 21981 30055 22015
rect 30055 21981 30064 22015
rect 30012 21972 30064 21981
rect 30748 22040 30800 22092
rect 26148 21904 26200 21956
rect 27988 21904 28040 21956
rect 25504 21836 25556 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 5540 21632 5592 21684
rect 8024 21632 8076 21684
rect 9680 21632 9732 21684
rect 9956 21675 10008 21684
rect 9956 21641 9965 21675
rect 9965 21641 9999 21675
rect 9999 21641 10008 21675
rect 9956 21632 10008 21641
rect 10416 21632 10468 21684
rect 2964 21564 3016 21616
rect 3700 21564 3752 21616
rect 8760 21564 8812 21616
rect 6460 21496 6512 21548
rect 6920 21496 6972 21548
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 9588 21564 9640 21616
rect 1400 21428 1452 21480
rect 3424 21471 3476 21480
rect 3424 21437 3433 21471
rect 3433 21437 3467 21471
rect 3467 21437 3476 21471
rect 3424 21428 3476 21437
rect 9128 21428 9180 21480
rect 8208 21360 8260 21412
rect 9312 21360 9364 21412
rect 28356 21496 28408 21548
rect 29552 21496 29604 21548
rect 9956 21428 10008 21480
rect 10784 21471 10836 21480
rect 10784 21437 10793 21471
rect 10793 21437 10827 21471
rect 10827 21437 10836 21471
rect 10784 21428 10836 21437
rect 28724 21471 28776 21480
rect 28724 21437 28733 21471
rect 28733 21437 28767 21471
rect 28767 21437 28776 21471
rect 28724 21428 28776 21437
rect 30564 21428 30616 21480
rect 31576 21471 31628 21480
rect 31576 21437 31585 21471
rect 31585 21437 31619 21471
rect 31619 21437 31628 21471
rect 31576 21428 31628 21437
rect 32772 21471 32824 21480
rect 32772 21437 32781 21471
rect 32781 21437 32815 21471
rect 32815 21437 32824 21471
rect 32772 21428 32824 21437
rect 3884 21292 3936 21344
rect 4712 21292 4764 21344
rect 6092 21292 6144 21344
rect 7472 21292 7524 21344
rect 8024 21292 8076 21344
rect 9036 21292 9088 21344
rect 10324 21292 10376 21344
rect 27620 21292 27672 21344
rect 31024 21292 31076 21344
rect 31116 21335 31168 21344
rect 31116 21301 31125 21335
rect 31125 21301 31159 21335
rect 31159 21301 31168 21335
rect 31116 21292 31168 21301
rect 31668 21292 31720 21344
rect 32956 21292 33008 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3424 21088 3476 21140
rect 5540 21088 5592 21140
rect 7012 21088 7064 21140
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 4620 20952 4672 21004
rect 6092 20995 6144 21004
rect 6092 20961 6101 20995
rect 6101 20961 6135 20995
rect 6135 20961 6144 20995
rect 6092 20952 6144 20961
rect 6920 20995 6972 21004
rect 6920 20961 6929 20995
rect 6929 20961 6963 20995
rect 6963 20961 6972 20995
rect 6920 20952 6972 20961
rect 7012 20995 7064 21004
rect 7012 20961 7021 20995
rect 7021 20961 7055 20995
rect 7055 20961 7064 20995
rect 7012 20952 7064 20961
rect 8300 21088 8352 21140
rect 7932 21020 7984 21072
rect 3884 20927 3936 20936
rect 3884 20893 3893 20927
rect 3893 20893 3927 20927
rect 3927 20893 3936 20927
rect 3884 20884 3936 20893
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 6368 20927 6420 20936
rect 6368 20893 6377 20927
rect 6377 20893 6411 20927
rect 6411 20893 6420 20927
rect 6368 20884 6420 20893
rect 7104 20884 7156 20936
rect 7472 20927 7524 20936
rect 7472 20893 7481 20927
rect 7481 20893 7515 20927
rect 7515 20893 7524 20927
rect 7472 20884 7524 20893
rect 8208 20952 8260 21004
rect 7932 20884 7984 20936
rect 8024 20927 8076 20936
rect 8024 20893 8033 20927
rect 8033 20893 8067 20927
rect 8067 20893 8076 20927
rect 8024 20884 8076 20893
rect 8300 20927 8352 20936
rect 8300 20893 8309 20927
rect 8309 20893 8343 20927
rect 8343 20893 8352 20927
rect 8300 20884 8352 20893
rect 9128 21020 9180 21072
rect 9956 21131 10008 21140
rect 9956 21097 9965 21131
rect 9965 21097 9999 21131
rect 9999 21097 10008 21131
rect 9956 21088 10008 21097
rect 8760 20952 8812 21004
rect 9864 21020 9916 21072
rect 10416 21088 10468 21140
rect 10784 21088 10836 21140
rect 29552 21131 29604 21140
rect 29552 21097 29561 21131
rect 29561 21097 29595 21131
rect 29595 21097 29604 21131
rect 29552 21088 29604 21097
rect 31576 21088 31628 21140
rect 32772 21088 32824 21140
rect 9312 20995 9364 21004
rect 9312 20961 9321 20995
rect 9321 20961 9355 20995
rect 9355 20961 9364 20995
rect 9312 20952 9364 20961
rect 9588 20884 9640 20936
rect 9680 20884 9732 20936
rect 10048 20995 10100 21004
rect 10048 20961 10057 20995
rect 10057 20961 10091 20995
rect 10091 20961 10100 20995
rect 10048 20952 10100 20961
rect 10324 20995 10376 21004
rect 10324 20961 10333 20995
rect 10333 20961 10367 20995
rect 10367 20961 10376 20995
rect 10324 20952 10376 20961
rect 23572 21020 23624 21072
rect 16856 20927 16908 20936
rect 16856 20893 16865 20927
rect 16865 20893 16899 20927
rect 16899 20893 16908 20927
rect 16856 20884 16908 20893
rect 23664 20952 23716 21004
rect 27620 20995 27672 21004
rect 27620 20961 27629 20995
rect 27629 20961 27663 20995
rect 27663 20961 27672 20995
rect 27620 20952 27672 20961
rect 27988 20952 28040 21004
rect 1676 20859 1728 20868
rect 1676 20825 1685 20859
rect 1685 20825 1719 20859
rect 1719 20825 1728 20859
rect 1676 20816 1728 20825
rect 2964 20816 3016 20868
rect 4804 20816 4856 20868
rect 10048 20816 10100 20868
rect 11060 20816 11112 20868
rect 16028 20816 16080 20868
rect 3148 20791 3200 20800
rect 3148 20757 3157 20791
rect 3157 20757 3191 20791
rect 3191 20757 3200 20791
rect 3148 20748 3200 20757
rect 6644 20748 6696 20800
rect 7840 20748 7892 20800
rect 8300 20748 8352 20800
rect 8944 20748 8996 20800
rect 9128 20791 9180 20800
rect 9128 20757 9137 20791
rect 9137 20757 9171 20791
rect 9171 20757 9180 20791
rect 9128 20748 9180 20757
rect 9772 20748 9824 20800
rect 16120 20748 16172 20800
rect 16580 20816 16632 20868
rect 17132 20859 17184 20868
rect 17132 20825 17141 20859
rect 17141 20825 17175 20859
rect 17175 20825 17184 20859
rect 17132 20816 17184 20825
rect 18144 20816 18196 20868
rect 22100 20859 22152 20868
rect 22100 20825 22109 20859
rect 22109 20825 22143 20859
rect 22143 20825 22152 20859
rect 22100 20816 22152 20825
rect 22836 20927 22888 20936
rect 22836 20893 22845 20927
rect 22845 20893 22879 20927
rect 22879 20893 22888 20927
rect 22836 20884 22888 20893
rect 24952 20884 25004 20936
rect 26976 20884 27028 20936
rect 17960 20748 18012 20800
rect 18052 20748 18104 20800
rect 20720 20791 20772 20800
rect 20720 20757 20729 20791
rect 20729 20757 20763 20791
rect 20763 20757 20772 20791
rect 20720 20748 20772 20757
rect 20812 20748 20864 20800
rect 22836 20748 22888 20800
rect 27068 20816 27120 20868
rect 31024 20995 31076 21004
rect 31024 20961 31033 20995
rect 31033 20961 31067 20995
rect 31067 20961 31076 20995
rect 31024 20952 31076 20961
rect 31760 20952 31812 21004
rect 33416 20884 33468 20936
rect 25136 20748 25188 20800
rect 28356 20748 28408 20800
rect 30748 20816 30800 20868
rect 32864 20816 32916 20868
rect 32956 20859 33008 20868
rect 32956 20825 32965 20859
rect 32965 20825 32999 20859
rect 32999 20825 33008 20859
rect 32956 20816 33008 20825
rect 33508 20816 33560 20868
rect 33968 20927 34020 20936
rect 33968 20893 33977 20927
rect 33977 20893 34011 20927
rect 34011 20893 34020 20927
rect 33968 20884 34020 20893
rect 34152 20884 34204 20936
rect 34980 20859 35032 20868
rect 34980 20825 34989 20859
rect 34989 20825 35023 20859
rect 35023 20825 35032 20859
rect 34980 20816 35032 20825
rect 35440 20816 35492 20868
rect 33968 20748 34020 20800
rect 34428 20748 34480 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 4804 20544 4856 20596
rect 6828 20544 6880 20596
rect 6644 20519 6696 20528
rect 6644 20485 6653 20519
rect 6653 20485 6687 20519
rect 6687 20485 6696 20519
rect 6644 20476 6696 20485
rect 8208 20544 8260 20596
rect 8300 20544 8352 20596
rect 3148 20408 3200 20460
rect 8116 20408 8168 20460
rect 9588 20587 9640 20596
rect 9588 20553 9597 20587
rect 9597 20553 9631 20587
rect 9631 20553 9640 20587
rect 9588 20544 9640 20553
rect 10048 20544 10100 20596
rect 11060 20476 11112 20528
rect 16120 20587 16172 20596
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 1676 20340 1728 20392
rect 2964 20340 3016 20392
rect 6368 20383 6420 20392
rect 6368 20349 6377 20383
rect 6377 20349 6411 20383
rect 6411 20349 6420 20383
rect 6368 20340 6420 20349
rect 8760 20383 8812 20392
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 8760 20340 8812 20349
rect 8944 20408 8996 20460
rect 15936 20476 15988 20528
rect 17132 20476 17184 20528
rect 19248 20476 19300 20528
rect 22100 20519 22152 20528
rect 22100 20485 22109 20519
rect 22109 20485 22143 20519
rect 22143 20485 22152 20519
rect 22100 20476 22152 20485
rect 22836 20544 22888 20596
rect 23664 20587 23716 20596
rect 23664 20553 23673 20587
rect 23673 20553 23707 20587
rect 23707 20553 23716 20587
rect 23664 20544 23716 20553
rect 22560 20476 22612 20528
rect 26148 20544 26200 20596
rect 26976 20544 27028 20596
rect 15568 20408 15620 20460
rect 11060 20383 11112 20392
rect 11060 20349 11069 20383
rect 11069 20349 11103 20383
rect 11103 20349 11112 20383
rect 11060 20340 11112 20349
rect 13820 20383 13872 20392
rect 13820 20349 13829 20383
rect 13829 20349 13863 20383
rect 13863 20349 13872 20383
rect 13820 20340 13872 20349
rect 7748 20272 7800 20324
rect 9680 20272 9732 20324
rect 16304 20383 16356 20392
rect 16304 20349 16313 20383
rect 16313 20349 16347 20383
rect 16347 20349 16356 20383
rect 16304 20340 16356 20349
rect 18420 20408 18472 20460
rect 18052 20340 18104 20392
rect 19156 20272 19208 20324
rect 15568 20247 15620 20256
rect 15568 20213 15577 20247
rect 15577 20213 15611 20247
rect 15611 20213 15620 20247
rect 15568 20204 15620 20213
rect 19524 20204 19576 20256
rect 20720 20340 20772 20392
rect 20812 20340 20864 20392
rect 22560 20340 22612 20392
rect 25136 20519 25188 20528
rect 25136 20485 25145 20519
rect 25145 20485 25179 20519
rect 25179 20485 25188 20519
rect 25136 20476 25188 20485
rect 26516 20408 26568 20460
rect 23664 20340 23716 20392
rect 25412 20383 25464 20392
rect 25412 20349 25421 20383
rect 25421 20349 25455 20383
rect 25455 20349 25464 20383
rect 25412 20340 25464 20349
rect 22284 20204 22336 20256
rect 25044 20204 25096 20256
rect 27988 20476 28040 20528
rect 30564 20544 30616 20596
rect 32772 20544 32824 20596
rect 32864 20544 32916 20596
rect 30748 20476 30800 20528
rect 31116 20476 31168 20528
rect 33324 20476 33376 20528
rect 35440 20544 35492 20596
rect 33508 20476 33560 20528
rect 34980 20476 35032 20528
rect 34152 20408 34204 20460
rect 34428 20451 34480 20460
rect 34428 20417 34437 20451
rect 34437 20417 34471 20451
rect 34471 20417 34480 20451
rect 34428 20408 34480 20417
rect 34520 20451 34572 20460
rect 34520 20417 34529 20451
rect 34529 20417 34563 20451
rect 34563 20417 34572 20451
rect 34520 20408 34572 20417
rect 27712 20340 27764 20392
rect 31760 20340 31812 20392
rect 33232 20340 33284 20392
rect 28448 20204 28500 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 1952 20000 2004 20052
rect 4068 20000 4120 20052
rect 7840 20000 7892 20052
rect 8024 20000 8076 20052
rect 8116 20043 8168 20052
rect 8116 20009 8125 20043
rect 8125 20009 8159 20043
rect 8159 20009 8168 20043
rect 8116 20000 8168 20009
rect 11060 20000 11112 20052
rect 18420 20043 18472 20052
rect 18420 20009 18429 20043
rect 18429 20009 18463 20043
rect 18463 20009 18472 20043
rect 18420 20000 18472 20009
rect 24860 20000 24912 20052
rect 26516 20043 26568 20052
rect 26516 20009 26525 20043
rect 26525 20009 26559 20043
rect 26559 20009 26568 20043
rect 26516 20000 26568 20009
rect 9772 19907 9824 19916
rect 9772 19873 9781 19907
rect 9781 19873 9815 19907
rect 9815 19873 9824 19907
rect 9772 19864 9824 19873
rect 19524 19864 19576 19916
rect 25412 19864 25464 19916
rect 26976 19864 27028 19916
rect 2412 19839 2464 19848
rect 2412 19805 2421 19839
rect 2421 19805 2455 19839
rect 2455 19805 2464 19839
rect 2412 19796 2464 19805
rect 2596 19839 2648 19848
rect 2596 19805 2605 19839
rect 2605 19805 2639 19839
rect 2639 19805 2648 19839
rect 2596 19796 2648 19805
rect 1768 19728 1820 19780
rect 3148 19771 3200 19780
rect 3148 19737 3157 19771
rect 3157 19737 3191 19771
rect 3191 19737 3200 19771
rect 3148 19728 3200 19737
rect 3884 19728 3936 19780
rect 8208 19796 8260 19848
rect 9864 19796 9916 19848
rect 7932 19771 7984 19780
rect 7932 19737 7957 19771
rect 7957 19737 7984 19771
rect 22284 19839 22336 19848
rect 22284 19805 22293 19839
rect 22293 19805 22327 19839
rect 22327 19805 22336 19839
rect 22284 19796 22336 19805
rect 26148 19796 26200 19848
rect 27068 19839 27120 19848
rect 27068 19805 27077 19839
rect 27077 19805 27111 19839
rect 27111 19805 27120 19839
rect 27068 19796 27120 19805
rect 27712 19907 27764 19916
rect 27712 19873 27721 19907
rect 27721 19873 27755 19907
rect 27755 19873 27764 19907
rect 27712 19864 27764 19873
rect 28448 19907 28500 19916
rect 28448 19873 28457 19907
rect 28457 19873 28491 19907
rect 28491 19873 28500 19907
rect 28448 19864 28500 19873
rect 7932 19728 7984 19737
rect 16856 19728 16908 19780
rect 2320 19660 2372 19712
rect 2596 19660 2648 19712
rect 2964 19703 3016 19712
rect 2964 19669 2991 19703
rect 2991 19669 3016 19703
rect 2964 19660 3016 19669
rect 3976 19660 4028 19712
rect 19248 19728 19300 19780
rect 17776 19660 17828 19712
rect 19800 19728 19852 19780
rect 22560 19771 22612 19780
rect 22560 19737 22569 19771
rect 22569 19737 22603 19771
rect 22603 19737 22612 19771
rect 22560 19728 22612 19737
rect 20904 19660 20956 19712
rect 20996 19703 21048 19712
rect 20996 19669 21005 19703
rect 21005 19669 21039 19703
rect 21039 19669 21048 19703
rect 20996 19660 21048 19669
rect 25044 19771 25096 19780
rect 25044 19737 25053 19771
rect 25053 19737 25087 19771
rect 25087 19737 25096 19771
rect 25044 19728 25096 19737
rect 26608 19771 26660 19780
rect 26608 19737 26617 19771
rect 26617 19737 26651 19771
rect 26651 19737 26660 19771
rect 26608 19728 26660 19737
rect 25136 19660 25188 19712
rect 26056 19660 26108 19712
rect 28356 19839 28408 19848
rect 28356 19805 28365 19839
rect 28365 19805 28399 19839
rect 28399 19805 28408 19839
rect 28356 19796 28408 19805
rect 29092 19728 29144 19780
rect 30196 19839 30248 19848
rect 30196 19805 30205 19839
rect 30205 19805 30239 19839
rect 30239 19805 30248 19839
rect 30196 19796 30248 19805
rect 30288 19839 30340 19848
rect 30288 19805 30297 19839
rect 30297 19805 30331 19839
rect 30331 19805 30340 19839
rect 30288 19796 30340 19805
rect 31116 19839 31168 19848
rect 31116 19805 31125 19839
rect 31125 19805 31159 19839
rect 31159 19805 31168 19839
rect 31116 19796 31168 19805
rect 34520 19864 34572 19916
rect 31392 19839 31444 19848
rect 31392 19805 31401 19839
rect 31401 19805 31435 19839
rect 31435 19805 31444 19839
rect 31392 19796 31444 19805
rect 30380 19728 30432 19780
rect 35348 19839 35400 19848
rect 35348 19805 35357 19839
rect 35357 19805 35391 19839
rect 35391 19805 35400 19839
rect 35348 19796 35400 19805
rect 34704 19771 34756 19780
rect 34704 19737 34713 19771
rect 34713 19737 34747 19771
rect 34747 19737 34756 19771
rect 34704 19728 34756 19737
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 2412 19456 2464 19508
rect 1768 19431 1820 19440
rect 1768 19397 1777 19431
rect 1777 19397 1811 19431
rect 1811 19397 1820 19431
rect 1768 19388 1820 19397
rect 1952 19431 2004 19440
rect 1952 19397 1961 19431
rect 1961 19397 1995 19431
rect 1995 19397 2004 19431
rect 1952 19388 2004 19397
rect 2964 19456 3016 19508
rect 8024 19456 8076 19508
rect 3056 19388 3108 19440
rect 6828 19388 6880 19440
rect 6920 19388 6972 19440
rect 16120 19456 16172 19508
rect 9404 19388 9456 19440
rect 16028 19388 16080 19440
rect 16580 19388 16632 19440
rect 3976 19320 4028 19372
rect 4620 19320 4672 19372
rect 4804 19320 4856 19372
rect 6368 19320 6420 19372
rect 10048 19320 10100 19372
rect 13820 19320 13872 19372
rect 17132 19363 17184 19372
rect 17132 19329 17141 19363
rect 17141 19329 17175 19363
rect 17175 19329 17184 19363
rect 17132 19320 17184 19329
rect 1400 19252 1452 19304
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 15016 19252 15068 19304
rect 18052 19388 18104 19440
rect 18420 19456 18472 19508
rect 22560 19456 22612 19508
rect 24860 19456 24912 19508
rect 25136 19456 25188 19508
rect 26148 19456 26200 19508
rect 27988 19456 28040 19508
rect 30472 19456 30524 19508
rect 34152 19456 34204 19508
rect 34520 19456 34572 19508
rect 18328 19431 18380 19440
rect 18328 19397 18337 19431
rect 18337 19397 18371 19431
rect 18371 19397 18380 19431
rect 18328 19388 18380 19397
rect 19800 19388 19852 19440
rect 26608 19388 26660 19440
rect 17776 19320 17828 19372
rect 20720 19320 20772 19372
rect 20812 19363 20864 19372
rect 20812 19329 20821 19363
rect 20821 19329 20855 19363
rect 20855 19329 20864 19363
rect 20812 19320 20864 19329
rect 20996 19320 21048 19372
rect 29276 19320 29328 19372
rect 31116 19320 31168 19372
rect 31944 19320 31996 19372
rect 35440 19320 35492 19372
rect 18604 19252 18656 19304
rect 23756 19295 23808 19304
rect 23756 19261 23765 19295
rect 23765 19261 23799 19295
rect 23799 19261 23808 19295
rect 23756 19252 23808 19261
rect 23664 19184 23716 19236
rect 26056 19252 26108 19304
rect 26976 19252 27028 19304
rect 31300 19252 31352 19304
rect 31760 19252 31812 19304
rect 33140 19252 33192 19304
rect 34704 19252 34756 19304
rect 4068 19116 4120 19168
rect 4620 19116 4672 19168
rect 15844 19159 15896 19168
rect 15844 19125 15853 19159
rect 15853 19125 15887 19159
rect 15887 19125 15896 19159
rect 15844 19116 15896 19125
rect 27068 19116 27120 19168
rect 29460 19116 29512 19168
rect 33232 19116 33284 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 8760 18955 8812 18964
rect 8760 18921 8769 18955
rect 8769 18921 8803 18955
rect 8803 18921 8812 18955
rect 8760 18912 8812 18921
rect 18328 18912 18380 18964
rect 16304 18844 16356 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 4068 18819 4120 18828
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 4528 18776 4580 18828
rect 7748 18776 7800 18828
rect 15016 18819 15068 18828
rect 15016 18785 15025 18819
rect 15025 18785 15059 18819
rect 15059 18785 15068 18819
rect 15016 18776 15068 18785
rect 15844 18776 15896 18828
rect 20904 18844 20956 18896
rect 19524 18819 19576 18828
rect 19524 18785 19533 18819
rect 19533 18785 19567 18819
rect 19567 18785 19576 18819
rect 19524 18776 19576 18785
rect 22376 18776 22428 18828
rect 1676 18683 1728 18692
rect 1676 18649 1685 18683
rect 1685 18649 1719 18683
rect 1719 18649 1728 18683
rect 1676 18640 1728 18649
rect 3056 18640 3108 18692
rect 3884 18708 3936 18760
rect 4252 18683 4304 18692
rect 4252 18649 4286 18683
rect 4286 18649 4304 18683
rect 4252 18640 4304 18649
rect 4620 18640 4672 18692
rect 3148 18615 3200 18624
rect 3148 18581 3157 18615
rect 3157 18581 3191 18615
rect 3191 18581 3200 18615
rect 3148 18572 3200 18581
rect 4804 18572 4856 18624
rect 5264 18572 5316 18624
rect 5632 18572 5684 18624
rect 6736 18640 6788 18692
rect 6828 18572 6880 18624
rect 6920 18572 6972 18624
rect 9404 18640 9456 18692
rect 15568 18708 15620 18760
rect 16856 18708 16908 18760
rect 24124 18708 24176 18760
rect 24768 18751 24820 18760
rect 27068 18912 27120 18964
rect 30288 18912 30340 18964
rect 31300 18955 31352 18964
rect 31300 18921 31309 18955
rect 31309 18921 31343 18955
rect 31343 18921 31352 18955
rect 31300 18912 31352 18921
rect 35348 18887 35400 18896
rect 35348 18853 35357 18887
rect 35357 18853 35391 18887
rect 35391 18853 35400 18887
rect 35348 18844 35400 18853
rect 24768 18717 24803 18751
rect 24803 18717 24820 18751
rect 24768 18708 24820 18717
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 26976 18708 27028 18760
rect 30380 18776 30432 18828
rect 31852 18776 31904 18828
rect 33324 18776 33376 18828
rect 35256 18708 35308 18760
rect 16212 18640 16264 18692
rect 17224 18683 17276 18692
rect 17224 18649 17233 18683
rect 17233 18649 17267 18683
rect 17267 18649 17276 18683
rect 17224 18640 17276 18649
rect 17960 18640 18012 18692
rect 19800 18683 19852 18692
rect 19800 18649 19809 18683
rect 19809 18649 19843 18683
rect 19843 18649 19852 18683
rect 19800 18640 19852 18649
rect 20812 18640 20864 18692
rect 7932 18572 7984 18624
rect 14924 18572 14976 18624
rect 16488 18615 16540 18624
rect 16488 18581 16497 18615
rect 16497 18581 16531 18615
rect 16531 18581 16540 18615
rect 16488 18572 16540 18581
rect 20720 18572 20772 18624
rect 21272 18615 21324 18624
rect 21272 18581 21281 18615
rect 21281 18581 21315 18615
rect 21315 18581 21324 18615
rect 21272 18572 21324 18581
rect 25596 18572 25648 18624
rect 27068 18640 27120 18692
rect 26332 18572 26384 18624
rect 28264 18640 28316 18692
rect 30840 18640 30892 18692
rect 33600 18640 33652 18692
rect 34796 18683 34848 18692
rect 34796 18649 34805 18683
rect 34805 18649 34839 18683
rect 34839 18649 34848 18683
rect 34796 18640 34848 18649
rect 29092 18572 29144 18624
rect 33784 18615 33836 18624
rect 33784 18581 33793 18615
rect 33793 18581 33827 18615
rect 33827 18581 33836 18615
rect 33784 18572 33836 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 3976 18411 4028 18420
rect 3976 18377 3985 18411
rect 3985 18377 4019 18411
rect 4019 18377 4028 18411
rect 3976 18368 4028 18377
rect 4528 18368 4580 18420
rect 4896 18368 4948 18420
rect 10048 18368 10100 18420
rect 16488 18368 16540 18420
rect 17224 18368 17276 18420
rect 5264 18300 5316 18352
rect 7656 18300 7708 18352
rect 7932 18300 7984 18352
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 3148 18232 3200 18284
rect 14924 18343 14976 18352
rect 14924 18309 14933 18343
rect 14933 18309 14967 18343
rect 14967 18309 14976 18343
rect 14924 18300 14976 18309
rect 15660 18300 15712 18352
rect 18328 18343 18380 18352
rect 18328 18309 18337 18343
rect 18337 18309 18371 18343
rect 18371 18309 18380 18343
rect 18328 18300 18380 18309
rect 19064 18300 19116 18352
rect 19800 18300 19852 18352
rect 1676 18164 1728 18216
rect 2596 18164 2648 18216
rect 9864 18207 9916 18216
rect 9864 18173 9873 18207
rect 9873 18173 9907 18207
rect 9907 18173 9916 18207
rect 9864 18164 9916 18173
rect 1400 18071 1452 18080
rect 1400 18037 1409 18071
rect 1409 18037 1443 18071
rect 1443 18037 1452 18071
rect 1400 18028 1452 18037
rect 4252 18096 4304 18148
rect 5080 18096 5132 18148
rect 4620 18028 4672 18080
rect 9404 18028 9456 18080
rect 13820 18232 13872 18284
rect 14280 18232 14332 18284
rect 20996 18300 21048 18352
rect 18604 18207 18656 18216
rect 18604 18173 18613 18207
rect 18613 18173 18647 18207
rect 18647 18173 18656 18207
rect 18604 18164 18656 18173
rect 22284 18275 22336 18284
rect 22284 18241 22293 18275
rect 22293 18241 22327 18275
rect 22327 18241 22336 18275
rect 22284 18232 22336 18241
rect 21272 18164 21324 18216
rect 22560 18207 22612 18216
rect 22560 18173 22569 18207
rect 22569 18173 22603 18207
rect 22603 18173 22612 18207
rect 22560 18164 22612 18173
rect 23756 18164 23808 18216
rect 24124 18207 24176 18216
rect 24124 18173 24133 18207
rect 24133 18173 24167 18207
rect 24167 18173 24176 18207
rect 24124 18164 24176 18173
rect 25596 18343 25648 18352
rect 25596 18309 25605 18343
rect 25605 18309 25639 18343
rect 25639 18309 25648 18343
rect 25596 18300 25648 18309
rect 29000 18368 29052 18420
rect 30196 18368 30248 18420
rect 28264 18300 28316 18352
rect 30932 18232 30984 18284
rect 31944 18300 31996 18352
rect 35348 18368 35400 18420
rect 33600 18300 33652 18352
rect 25136 18164 25188 18216
rect 26976 18207 27028 18216
rect 26976 18173 26985 18207
rect 26985 18173 27019 18207
rect 27019 18173 27028 18207
rect 26976 18164 27028 18173
rect 27620 18164 27672 18216
rect 31208 18207 31260 18216
rect 31208 18173 31217 18207
rect 31217 18173 31251 18207
rect 31251 18173 31260 18207
rect 31208 18164 31260 18173
rect 31760 18164 31812 18216
rect 32128 18164 32180 18216
rect 22008 18096 22060 18148
rect 31576 18096 31628 18148
rect 33416 18164 33468 18216
rect 35256 18164 35308 18216
rect 11336 18071 11388 18080
rect 11336 18037 11345 18071
rect 11345 18037 11379 18071
rect 11379 18037 11388 18071
rect 11336 18028 11388 18037
rect 23664 18028 23716 18080
rect 27896 18028 27948 18080
rect 28724 18028 28776 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1584 17824 1636 17876
rect 4712 17824 4764 17876
rect 9864 17824 9916 17876
rect 11336 17824 11388 17876
rect 19064 17867 19116 17876
rect 19064 17833 19073 17867
rect 19073 17833 19107 17867
rect 19107 17833 19116 17867
rect 19064 17824 19116 17833
rect 22376 17867 22428 17876
rect 22376 17833 22385 17867
rect 22385 17833 22419 17867
rect 22419 17833 22428 17867
rect 22376 17824 22428 17833
rect 22560 17824 22612 17876
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 26240 17824 26292 17876
rect 27620 17824 27672 17876
rect 31944 17824 31996 17876
rect 33324 17867 33376 17876
rect 33324 17833 33333 17867
rect 33333 17833 33367 17867
rect 33367 17833 33376 17867
rect 33324 17824 33376 17833
rect 1492 17620 1544 17672
rect 3884 17620 3936 17672
rect 4896 17688 4948 17740
rect 4528 17663 4580 17672
rect 4528 17629 4537 17663
rect 4537 17629 4571 17663
rect 4571 17629 4580 17663
rect 4528 17620 4580 17629
rect 4620 17663 4672 17672
rect 4620 17629 4629 17663
rect 4629 17629 4663 17663
rect 4663 17629 4672 17663
rect 4620 17620 4672 17629
rect 5080 17663 5132 17672
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 6920 17688 6972 17740
rect 9864 17620 9916 17672
rect 14280 17688 14332 17740
rect 16856 17688 16908 17740
rect 22284 17688 22336 17740
rect 23664 17688 23716 17740
rect 26240 17688 26292 17740
rect 4712 17552 4764 17604
rect 6552 17595 6604 17604
rect 6552 17561 6561 17595
rect 6561 17561 6595 17595
rect 6595 17561 6604 17595
rect 6552 17552 6604 17561
rect 6828 17552 6880 17604
rect 3424 17484 3476 17536
rect 4344 17484 4396 17536
rect 5264 17527 5316 17536
rect 5264 17493 5273 17527
rect 5273 17493 5307 17527
rect 5307 17493 5316 17527
rect 5264 17484 5316 17493
rect 7472 17484 7524 17536
rect 10508 17620 10560 17672
rect 11336 17620 11388 17672
rect 14556 17552 14608 17604
rect 11060 17527 11112 17536
rect 11060 17493 11069 17527
rect 11069 17493 11103 17527
rect 11103 17493 11112 17527
rect 11060 17484 11112 17493
rect 16028 17663 16080 17672
rect 16028 17629 16037 17663
rect 16037 17629 16071 17663
rect 16071 17629 16080 17663
rect 16028 17620 16080 17629
rect 23756 17663 23808 17672
rect 23756 17629 23765 17663
rect 23765 17629 23799 17663
rect 23799 17629 23808 17663
rect 23756 17620 23808 17629
rect 24124 17620 24176 17672
rect 29000 17688 29052 17740
rect 31852 17688 31904 17740
rect 26976 17620 27028 17672
rect 33784 17731 33836 17740
rect 33784 17697 33793 17731
rect 33793 17697 33827 17731
rect 33827 17697 33836 17731
rect 33784 17688 33836 17697
rect 33048 17620 33100 17672
rect 33416 17620 33468 17672
rect 34796 17688 34848 17740
rect 16488 17552 16540 17604
rect 17868 17552 17920 17604
rect 18052 17552 18104 17604
rect 20904 17595 20956 17604
rect 20904 17561 20913 17595
rect 20913 17561 20947 17595
rect 20947 17561 20956 17595
rect 20904 17552 20956 17561
rect 20996 17552 21048 17604
rect 25596 17552 25648 17604
rect 26332 17552 26384 17604
rect 28172 17595 28224 17604
rect 28172 17561 28181 17595
rect 28181 17561 28215 17595
rect 28215 17561 28224 17595
rect 28172 17552 28224 17561
rect 28724 17552 28776 17604
rect 30472 17552 30524 17604
rect 30840 17552 30892 17604
rect 18604 17484 18656 17536
rect 21640 17484 21692 17536
rect 26884 17484 26936 17536
rect 34060 17484 34112 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 1492 17144 1544 17196
rect 3056 17144 3108 17196
rect 3424 17212 3476 17264
rect 3792 17255 3844 17264
rect 3792 17221 3817 17255
rect 3817 17221 3844 17255
rect 3792 17212 3844 17221
rect 4620 17280 4672 17332
rect 4712 17280 4764 17332
rect 6552 17280 6604 17332
rect 17868 17280 17920 17332
rect 19064 17323 19116 17332
rect 19064 17289 19073 17323
rect 19073 17289 19107 17323
rect 19107 17289 19116 17323
rect 19064 17280 19116 17289
rect 22376 17280 22428 17332
rect 4344 17255 4396 17264
rect 4344 17221 4353 17255
rect 4353 17221 4387 17255
rect 4387 17221 4396 17255
rect 4344 17212 4396 17221
rect 5632 17212 5684 17264
rect 6920 17212 6972 17264
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 7932 17212 7984 17264
rect 9404 17212 9456 17264
rect 14556 17255 14608 17264
rect 14556 17221 14565 17255
rect 14565 17221 14599 17255
rect 14599 17221 14608 17255
rect 14556 17212 14608 17221
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 3424 16983 3476 16992
rect 3424 16949 3433 16983
rect 3433 16949 3467 16983
rect 3467 16949 3476 16983
rect 3424 16940 3476 16949
rect 4712 17076 4764 17128
rect 4528 16940 4580 16992
rect 8024 17119 8076 17128
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 9864 17144 9916 17196
rect 11060 17144 11112 17196
rect 14096 17144 14148 17196
rect 14280 17187 14332 17196
rect 14280 17153 14289 17187
rect 14289 17153 14323 17187
rect 14323 17153 14332 17187
rect 14280 17144 14332 17153
rect 15660 17144 15712 17196
rect 17592 17212 17644 17264
rect 20812 17212 20864 17264
rect 22284 17212 22336 17264
rect 20444 17144 20496 17196
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 16856 17119 16908 17128
rect 16856 17085 16865 17119
rect 16865 17085 16899 17119
rect 16899 17085 16908 17119
rect 16856 17076 16908 17085
rect 17776 17076 17828 17128
rect 18512 17076 18564 17128
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 26240 17280 26292 17332
rect 26884 17280 26936 17332
rect 34060 17280 34112 17332
rect 25596 17212 25648 17264
rect 28816 17212 28868 17264
rect 30656 17212 30708 17264
rect 31760 17212 31812 17264
rect 29000 17187 29052 17196
rect 29000 17153 29009 17187
rect 29009 17153 29043 17187
rect 29043 17153 29052 17187
rect 29000 17144 29052 17153
rect 29552 17187 29604 17196
rect 29552 17153 29561 17187
rect 29561 17153 29595 17187
rect 29595 17153 29604 17187
rect 29552 17144 29604 17153
rect 31944 17187 31996 17196
rect 31944 17153 31953 17187
rect 31953 17153 31987 17187
rect 31987 17153 31996 17187
rect 31944 17144 31996 17153
rect 33508 17144 33560 17196
rect 18236 17008 18288 17060
rect 21640 17008 21692 17060
rect 26792 17076 26844 17128
rect 29828 17119 29880 17128
rect 29828 17085 29837 17119
rect 29837 17085 29871 17119
rect 29871 17085 29880 17119
rect 29828 17076 29880 17085
rect 8576 16940 8628 16992
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 9588 16983 9640 16992
rect 9588 16949 9597 16983
rect 9597 16949 9631 16983
rect 9631 16949 9640 16983
rect 9588 16940 9640 16949
rect 10876 16940 10928 16992
rect 16028 16983 16080 16992
rect 16028 16949 16037 16983
rect 16037 16949 16071 16983
rect 16071 16949 16080 16983
rect 16028 16940 16080 16949
rect 16396 16940 16448 16992
rect 16488 16940 16540 16992
rect 19340 16940 19392 16992
rect 21916 16940 21968 16992
rect 27804 16940 27856 16992
rect 31208 16940 31260 16992
rect 31944 16940 31996 16992
rect 32128 17119 32180 17128
rect 32128 17085 32137 17119
rect 32137 17085 32171 17119
rect 32171 17085 32180 17119
rect 32128 17076 32180 17085
rect 32404 17119 32456 17128
rect 32404 17085 32413 17119
rect 32413 17085 32447 17119
rect 32447 17085 32456 17119
rect 32404 17076 32456 17085
rect 33048 17076 33100 17128
rect 34244 17119 34296 17128
rect 34244 17085 34253 17119
rect 34253 17085 34287 17119
rect 34287 17085 34296 17119
rect 34244 17076 34296 17085
rect 33416 16940 33468 16992
rect 33508 16940 33560 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1952 16736 2004 16788
rect 4436 16736 4488 16788
rect 5264 16736 5316 16788
rect 8024 16736 8076 16788
rect 2228 16643 2280 16652
rect 2228 16609 2237 16643
rect 2237 16609 2271 16643
rect 2271 16609 2280 16643
rect 2228 16600 2280 16609
rect 3424 16532 3476 16584
rect 3976 16532 4028 16584
rect 4068 16575 4120 16584
rect 4068 16541 4077 16575
rect 4077 16541 4111 16575
rect 4111 16541 4120 16575
rect 4068 16532 4120 16541
rect 4804 16668 4856 16720
rect 4620 16600 4672 16652
rect 4436 16575 4488 16584
rect 4436 16541 4445 16575
rect 4445 16541 4479 16575
rect 4479 16541 4488 16575
rect 4436 16532 4488 16541
rect 9588 16736 9640 16788
rect 11060 16736 11112 16788
rect 20444 16779 20496 16788
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 25688 16736 25740 16788
rect 26792 16779 26844 16788
rect 26792 16745 26801 16779
rect 26801 16745 26835 16779
rect 26835 16745 26844 16779
rect 26792 16736 26844 16745
rect 27068 16736 27120 16788
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 9496 16668 9548 16720
rect 29552 16736 29604 16788
rect 10048 16600 10100 16652
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 14096 16643 14148 16652
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14096 16600 14148 16609
rect 15936 16600 15988 16652
rect 18972 16600 19024 16652
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 21916 16600 21968 16609
rect 22284 16600 22336 16652
rect 26148 16600 26200 16652
rect 27528 16643 27580 16652
rect 27528 16609 27537 16643
rect 27537 16609 27571 16643
rect 27571 16609 27580 16643
rect 27528 16600 27580 16609
rect 27804 16643 27856 16652
rect 27804 16609 27813 16643
rect 27813 16609 27847 16643
rect 27847 16609 27856 16643
rect 27804 16600 27856 16609
rect 9864 16532 9916 16584
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 5540 16464 5592 16516
rect 7288 16464 7340 16516
rect 9404 16464 9456 16516
rect 11336 16464 11388 16516
rect 15660 16464 15712 16516
rect 17316 16507 17368 16516
rect 17316 16473 17325 16507
rect 17325 16473 17359 16507
rect 17359 16473 17368 16507
rect 17316 16464 17368 16473
rect 18420 16575 18472 16584
rect 18420 16541 18429 16575
rect 18429 16541 18463 16575
rect 18463 16541 18472 16575
rect 18420 16532 18472 16541
rect 18512 16575 18564 16584
rect 18512 16541 18521 16575
rect 18521 16541 18555 16575
rect 18555 16541 18564 16575
rect 18512 16532 18564 16541
rect 26884 16532 26936 16584
rect 30656 16532 30708 16584
rect 20628 16464 20680 16516
rect 20904 16464 20956 16516
rect 22652 16507 22704 16516
rect 22652 16473 22661 16507
rect 22661 16473 22695 16507
rect 22695 16473 22704 16507
rect 22652 16464 22704 16473
rect 23940 16464 23992 16516
rect 4712 16396 4764 16448
rect 15844 16439 15896 16448
rect 15844 16405 15853 16439
rect 15853 16405 15887 16439
rect 15887 16405 15896 16439
rect 15844 16396 15896 16405
rect 25044 16396 25096 16448
rect 25596 16464 25648 16516
rect 25964 16396 26016 16448
rect 29276 16464 29328 16516
rect 33508 16736 33560 16788
rect 31760 16668 31812 16720
rect 32128 16668 32180 16720
rect 32036 16600 32088 16652
rect 32404 16643 32456 16652
rect 32404 16609 32413 16643
rect 32413 16609 32447 16643
rect 32447 16609 32456 16643
rect 32404 16600 32456 16609
rect 33048 16600 33100 16652
rect 36452 16643 36504 16652
rect 36452 16609 36461 16643
rect 36461 16609 36495 16643
rect 36495 16609 36504 16643
rect 36452 16600 36504 16609
rect 31944 16575 31996 16584
rect 31944 16541 31953 16575
rect 31953 16541 31987 16575
rect 31987 16541 31996 16575
rect 31944 16532 31996 16541
rect 31668 16464 31720 16516
rect 29828 16396 29880 16448
rect 29920 16396 29972 16448
rect 36636 16507 36688 16516
rect 36636 16473 36645 16507
rect 36645 16473 36679 16507
rect 36679 16473 36688 16507
rect 36636 16464 36688 16473
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 3424 16192 3476 16244
rect 4068 16235 4120 16244
rect 4068 16201 4077 16235
rect 4077 16201 4111 16235
rect 4111 16201 4120 16235
rect 4068 16192 4120 16201
rect 2228 16099 2280 16108
rect 2228 16065 2243 16099
rect 2243 16065 2277 16099
rect 2277 16065 2280 16099
rect 10508 16167 10560 16176
rect 10508 16133 10517 16167
rect 10517 16133 10551 16167
rect 10551 16133 10560 16167
rect 10508 16124 10560 16133
rect 2228 16056 2280 16065
rect 3424 16056 3476 16108
rect 3700 16099 3752 16108
rect 3700 16065 3709 16099
rect 3709 16065 3743 16099
rect 3743 16065 3752 16099
rect 3700 16056 3752 16065
rect 3884 16056 3936 16108
rect 14280 16056 14332 16108
rect 17132 16192 17184 16244
rect 15660 16124 15712 16176
rect 15292 16056 15344 16108
rect 15844 16056 15896 16108
rect 18604 16056 18656 16108
rect 18972 16056 19024 16108
rect 19524 16192 19576 16244
rect 20812 16235 20864 16244
rect 20812 16201 20821 16235
rect 20821 16201 20855 16235
rect 20855 16201 20864 16235
rect 20812 16192 20864 16201
rect 21824 16192 21876 16244
rect 26608 16192 26660 16244
rect 19340 16167 19392 16176
rect 19340 16133 19349 16167
rect 19349 16133 19383 16167
rect 19383 16133 19392 16167
rect 19340 16124 19392 16133
rect 22652 16167 22704 16176
rect 22652 16133 22661 16167
rect 22661 16133 22695 16167
rect 22695 16133 22704 16167
rect 22652 16124 22704 16133
rect 23940 16124 23992 16176
rect 25964 16167 26016 16176
rect 25964 16133 25973 16167
rect 25973 16133 26007 16167
rect 26007 16133 26016 16167
rect 25964 16124 26016 16133
rect 28172 16192 28224 16244
rect 29092 16192 29144 16244
rect 33508 16235 33560 16244
rect 33508 16201 33517 16235
rect 33517 16201 33551 16235
rect 33551 16201 33560 16235
rect 33508 16192 33560 16201
rect 34244 16192 34296 16244
rect 4068 15988 4120 16040
rect 7656 15988 7708 16040
rect 14372 15988 14424 16040
rect 15476 16031 15528 16040
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 18788 15988 18840 16040
rect 19984 15988 20036 16040
rect 21824 16056 21876 16108
rect 23112 16099 23164 16108
rect 23112 16065 23121 16099
rect 23121 16065 23155 16099
rect 23155 16065 23164 16099
rect 23112 16056 23164 16065
rect 23296 16099 23348 16108
rect 23296 16065 23305 16099
rect 23305 16065 23339 16099
rect 23339 16065 23348 16099
rect 23296 16056 23348 16065
rect 20904 15988 20956 16040
rect 3148 15920 3200 15972
rect 7748 15920 7800 15972
rect 11060 15920 11112 15972
rect 1676 15852 1728 15904
rect 7196 15852 7248 15904
rect 10876 15852 10928 15904
rect 18420 15852 18472 15904
rect 23756 16031 23808 16040
rect 23756 15997 23765 16031
rect 23765 15997 23799 16031
rect 23799 15997 23808 16031
rect 23756 15988 23808 15997
rect 24400 15988 24452 16040
rect 25504 16031 25556 16040
rect 25504 15997 25513 16031
rect 25513 15997 25547 16031
rect 25547 15997 25556 16031
rect 27528 16124 27580 16176
rect 29000 16124 29052 16176
rect 30656 16124 30708 16176
rect 34060 16124 34112 16176
rect 25504 15988 25556 15997
rect 26332 15988 26384 16040
rect 28540 15988 28592 16040
rect 28908 16031 28960 16040
rect 28908 15997 28917 16031
rect 28917 15997 28951 16031
rect 28951 15997 28960 16031
rect 28908 15988 28960 15997
rect 29276 15988 29328 16040
rect 31760 16099 31812 16108
rect 31760 16065 31769 16099
rect 31769 16065 31803 16099
rect 31803 16065 31812 16099
rect 31760 16056 31812 16065
rect 30840 16031 30892 16040
rect 30840 15997 30849 16031
rect 30849 15997 30883 16031
rect 30883 15997 30892 16031
rect 30840 15988 30892 15997
rect 31944 15988 31996 16040
rect 32772 16031 32824 16040
rect 32772 15997 32781 16031
rect 32781 15997 32815 16031
rect 32815 15997 32824 16031
rect 32772 15988 32824 15997
rect 33140 15988 33192 16040
rect 25688 15963 25740 15972
rect 25688 15929 25697 15963
rect 25697 15929 25731 15963
rect 25731 15929 25740 15963
rect 25688 15920 25740 15929
rect 25044 15852 25096 15904
rect 28172 15852 28224 15904
rect 29920 15852 29972 15904
rect 32220 15895 32272 15904
rect 32220 15861 32229 15895
rect 32229 15861 32263 15895
rect 32263 15861 32272 15895
rect 32220 15852 32272 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 3884 15648 3936 15700
rect 10508 15691 10560 15700
rect 10508 15657 10517 15691
rect 10517 15657 10551 15691
rect 10551 15657 10560 15691
rect 10508 15648 10560 15657
rect 15476 15648 15528 15700
rect 15660 15648 15712 15700
rect 15936 15691 15988 15700
rect 15936 15657 15945 15691
rect 15945 15657 15979 15691
rect 15979 15657 15988 15691
rect 15936 15648 15988 15657
rect 23296 15648 23348 15700
rect 28908 15648 28960 15700
rect 1676 15555 1728 15564
rect 1676 15521 1685 15555
rect 1685 15521 1719 15555
rect 1719 15521 1728 15555
rect 1676 15512 1728 15521
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 7196 15555 7248 15564
rect 7196 15521 7205 15555
rect 7205 15521 7239 15555
rect 7239 15521 7248 15555
rect 7196 15512 7248 15521
rect 7656 15512 7708 15564
rect 3516 15444 3568 15496
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 6920 15487 6972 15496
rect 6920 15453 6929 15487
rect 6929 15453 6963 15487
rect 6963 15453 6972 15487
rect 6920 15444 6972 15453
rect 3056 15376 3108 15428
rect 3148 15376 3200 15428
rect 5540 15376 5592 15428
rect 10600 15555 10652 15564
rect 10600 15521 10609 15555
rect 10609 15521 10643 15555
rect 10643 15521 10652 15555
rect 10600 15512 10652 15521
rect 10876 15555 10928 15564
rect 10876 15521 10885 15555
rect 10885 15521 10919 15555
rect 10919 15521 10928 15555
rect 10876 15512 10928 15521
rect 14372 15555 14424 15564
rect 14372 15521 14381 15555
rect 14381 15521 14415 15555
rect 14415 15521 14424 15555
rect 14372 15512 14424 15521
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 15568 15512 15620 15564
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 16856 15555 16908 15564
rect 16856 15521 16865 15555
rect 16865 15521 16899 15555
rect 16899 15521 16908 15555
rect 16856 15512 16908 15521
rect 10048 15376 10100 15428
rect 11336 15376 11388 15428
rect 15844 15444 15896 15496
rect 14280 15376 14332 15428
rect 15936 15376 15988 15428
rect 16212 15376 16264 15428
rect 18420 15512 18472 15564
rect 31944 15580 31996 15632
rect 32036 15580 32088 15632
rect 18788 15555 18840 15564
rect 18788 15521 18797 15555
rect 18797 15521 18831 15555
rect 18831 15521 18840 15555
rect 18788 15512 18840 15521
rect 20720 15512 20772 15564
rect 20812 15512 20864 15564
rect 17316 15376 17368 15428
rect 3332 15308 3384 15360
rect 3700 15308 3752 15360
rect 4068 15308 4120 15360
rect 7288 15308 7340 15360
rect 8024 15308 8076 15360
rect 8484 15308 8536 15360
rect 9220 15308 9272 15360
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 10140 15351 10192 15360
rect 10140 15317 10149 15351
rect 10149 15317 10183 15351
rect 10183 15317 10192 15351
rect 10140 15308 10192 15317
rect 10600 15308 10652 15360
rect 17960 15376 18012 15428
rect 20628 15487 20680 15496
rect 20628 15453 20637 15487
rect 20637 15453 20671 15487
rect 20671 15453 20680 15487
rect 20628 15444 20680 15453
rect 23112 15512 23164 15564
rect 20720 15419 20772 15428
rect 20720 15385 20729 15419
rect 20729 15385 20763 15419
rect 20763 15385 20772 15419
rect 20720 15376 20772 15385
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 24400 15555 24452 15564
rect 24400 15521 24409 15555
rect 24409 15521 24443 15555
rect 24443 15521 24452 15555
rect 24400 15512 24452 15521
rect 25504 15512 25556 15564
rect 27896 15512 27948 15564
rect 28724 15512 28776 15564
rect 21916 15308 21968 15360
rect 22100 15419 22152 15428
rect 22100 15385 22109 15419
rect 22109 15385 22143 15419
rect 22143 15385 22152 15419
rect 22100 15376 22152 15385
rect 23848 15376 23900 15428
rect 25044 15487 25096 15496
rect 25044 15453 25053 15487
rect 25053 15453 25087 15487
rect 25087 15453 25096 15487
rect 25044 15444 25096 15453
rect 28816 15444 28868 15496
rect 29000 15512 29052 15564
rect 32220 15512 32272 15564
rect 33508 15512 33560 15564
rect 27068 15376 27120 15428
rect 29092 15376 29144 15428
rect 22284 15308 22336 15360
rect 27620 15351 27672 15360
rect 27620 15317 27629 15351
rect 27629 15317 27663 15351
rect 27663 15317 27672 15351
rect 27620 15308 27672 15317
rect 28080 15351 28132 15360
rect 28080 15317 28089 15351
rect 28089 15317 28123 15351
rect 28123 15317 28132 15351
rect 28080 15308 28132 15317
rect 29552 15308 29604 15360
rect 30564 15376 30616 15428
rect 31392 15419 31444 15428
rect 31392 15385 31401 15419
rect 31401 15385 31435 15419
rect 31435 15385 31444 15419
rect 31392 15376 31444 15385
rect 30472 15308 30524 15360
rect 30840 15308 30892 15360
rect 31576 15308 31628 15360
rect 31944 15444 31996 15496
rect 32128 15487 32180 15496
rect 32128 15453 32137 15487
rect 32137 15453 32171 15487
rect 32171 15453 32180 15487
rect 32128 15444 32180 15453
rect 33416 15444 33468 15496
rect 34520 15308 34572 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 3516 15147 3568 15156
rect 3516 15113 3525 15147
rect 3525 15113 3559 15147
rect 3559 15113 3568 15147
rect 3516 15104 3568 15113
rect 7288 15147 7340 15156
rect 7288 15113 7297 15147
rect 7297 15113 7331 15147
rect 7331 15113 7340 15147
rect 7288 15104 7340 15113
rect 7656 15147 7708 15156
rect 7656 15113 7665 15147
rect 7665 15113 7699 15147
rect 7699 15113 7708 15147
rect 7656 15104 7708 15113
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 10324 15104 10376 15156
rect 3148 15079 3200 15088
rect 3148 15045 3157 15079
rect 3157 15045 3191 15079
rect 3191 15045 3200 15079
rect 3148 15036 3200 15045
rect 3240 15036 3292 15088
rect 4068 15036 4120 15088
rect 5724 15079 5776 15088
rect 5724 15045 5733 15079
rect 5733 15045 5767 15079
rect 5767 15045 5776 15079
rect 5724 15036 5776 15045
rect 7932 15036 7984 15088
rect 10140 15036 10192 15088
rect 8484 14968 8536 15020
rect 5724 14832 5776 14884
rect 7932 14943 7984 14952
rect 7932 14909 7941 14943
rect 7941 14909 7975 14943
rect 7975 14909 7984 14943
rect 7932 14900 7984 14909
rect 8024 14943 8076 14952
rect 8024 14909 8033 14943
rect 8033 14909 8067 14943
rect 8067 14909 8076 14943
rect 8024 14900 8076 14909
rect 6736 14832 6788 14884
rect 3332 14807 3384 14816
rect 3332 14773 3341 14807
rect 3341 14773 3375 14807
rect 3375 14773 3384 14807
rect 3332 14764 3384 14773
rect 5264 14764 5316 14816
rect 5632 14764 5684 14816
rect 8852 14943 8904 14952
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 10600 14968 10652 14977
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 19064 15104 19116 15156
rect 19984 15036 20036 15088
rect 20720 15104 20772 15156
rect 22100 15104 22152 15156
rect 23296 15147 23348 15156
rect 23296 15113 23305 15147
rect 23305 15113 23339 15147
rect 23339 15113 23348 15147
rect 23296 15104 23348 15113
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 21824 15036 21876 15088
rect 23756 15036 23808 15088
rect 24400 15036 24452 15088
rect 26148 15036 26200 15088
rect 27620 15036 27672 15088
rect 27804 15036 27856 15088
rect 28816 15147 28868 15156
rect 28816 15113 28825 15147
rect 28825 15113 28859 15147
rect 28859 15113 28868 15147
rect 28816 15104 28868 15113
rect 30472 15104 30524 15156
rect 32772 15104 32824 15156
rect 34612 15104 34664 15156
rect 30656 15036 30708 15088
rect 33600 15036 33652 15088
rect 21916 15011 21968 15020
rect 21916 14977 21925 15011
rect 21925 14977 21959 15011
rect 21959 14977 21968 15011
rect 21916 14968 21968 14977
rect 26332 14968 26384 15020
rect 31300 14968 31352 15020
rect 10048 14900 10100 14952
rect 10784 14943 10836 14952
rect 10784 14909 10793 14943
rect 10793 14909 10827 14943
rect 10827 14909 10836 14943
rect 10784 14900 10836 14909
rect 15568 14900 15620 14952
rect 15752 14943 15804 14952
rect 15752 14909 15761 14943
rect 15761 14909 15795 14943
rect 15795 14909 15804 14943
rect 15752 14900 15804 14909
rect 16672 14943 16724 14952
rect 16672 14909 16681 14943
rect 16681 14909 16715 14943
rect 16715 14909 16724 14943
rect 16672 14900 16724 14909
rect 17592 14900 17644 14952
rect 21456 14900 21508 14952
rect 11336 14832 11388 14884
rect 23664 14900 23716 14952
rect 25964 14943 26016 14952
rect 25964 14909 25973 14943
rect 25973 14909 26007 14943
rect 26007 14909 26016 14943
rect 25964 14900 26016 14909
rect 26240 14900 26292 14952
rect 23940 14832 23992 14884
rect 24860 14832 24912 14884
rect 30840 14900 30892 14952
rect 9864 14764 9916 14816
rect 17960 14764 18012 14816
rect 25504 14807 25556 14816
rect 25504 14773 25513 14807
rect 25513 14773 25547 14807
rect 25547 14773 25556 14807
rect 25504 14764 25556 14773
rect 31760 14764 31812 14816
rect 32864 14943 32916 14952
rect 32864 14909 32873 14943
rect 32873 14909 32907 14943
rect 32907 14909 32916 14943
rect 32864 14900 32916 14909
rect 33600 14900 33652 14952
rect 34428 14943 34480 14952
rect 34428 14909 34437 14943
rect 34437 14909 34471 14943
rect 34471 14909 34480 14943
rect 34428 14900 34480 14909
rect 34704 14943 34756 14952
rect 34704 14909 34713 14943
rect 34713 14909 34747 14943
rect 34747 14909 34756 14943
rect 34704 14900 34756 14909
rect 34336 14807 34388 14816
rect 34336 14773 34345 14807
rect 34345 14773 34379 14807
rect 34379 14773 34388 14807
rect 34336 14764 34388 14773
rect 35440 14764 35492 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 6736 14603 6788 14612
rect 6736 14569 6745 14603
rect 6745 14569 6779 14603
rect 6779 14569 6788 14603
rect 6736 14560 6788 14569
rect 1676 14467 1728 14476
rect 1676 14433 1685 14467
rect 1685 14433 1719 14467
rect 1719 14433 1728 14467
rect 1676 14424 1728 14433
rect 1860 14424 1912 14476
rect 3240 14356 3292 14408
rect 3516 14356 3568 14408
rect 4620 14424 4672 14476
rect 5264 14467 5316 14476
rect 5264 14433 5273 14467
rect 5273 14433 5307 14467
rect 5307 14433 5316 14467
rect 5264 14424 5316 14433
rect 10784 14560 10836 14612
rect 15752 14560 15804 14612
rect 23940 14603 23992 14612
rect 23940 14569 23949 14603
rect 23949 14569 23983 14603
rect 23983 14569 23992 14603
rect 23940 14560 23992 14569
rect 28080 14560 28132 14612
rect 32128 14560 32180 14612
rect 33508 14603 33560 14612
rect 33508 14569 33517 14603
rect 33517 14569 33551 14603
rect 33551 14569 33560 14603
rect 33508 14560 33560 14569
rect 9680 14424 9732 14476
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 11336 14424 11388 14476
rect 14280 14424 14332 14476
rect 16672 14424 16724 14476
rect 18604 14467 18656 14476
rect 18604 14433 18613 14467
rect 18613 14433 18647 14467
rect 18647 14433 18656 14467
rect 18604 14424 18656 14433
rect 21824 14424 21876 14476
rect 24400 14467 24452 14476
rect 24400 14433 24409 14467
rect 24409 14433 24443 14467
rect 24443 14433 24452 14467
rect 24400 14424 24452 14433
rect 31392 14467 31444 14476
rect 31392 14433 31401 14467
rect 31401 14433 31435 14467
rect 31435 14433 31444 14467
rect 31392 14424 31444 14433
rect 31760 14467 31812 14476
rect 31760 14433 31769 14467
rect 31769 14433 31803 14467
rect 31803 14433 31812 14467
rect 31760 14424 31812 14433
rect 32036 14467 32088 14476
rect 32036 14433 32045 14467
rect 32045 14433 32079 14467
rect 32079 14433 32088 14467
rect 32036 14424 32088 14433
rect 34704 14467 34756 14476
rect 34704 14433 34713 14467
rect 34713 14433 34747 14467
rect 34747 14433 34756 14467
rect 34704 14424 34756 14433
rect 35440 14467 35492 14476
rect 35440 14433 35449 14467
rect 35449 14433 35483 14467
rect 35483 14433 35492 14467
rect 35440 14424 35492 14433
rect 2964 14288 3016 14340
rect 3332 14288 3384 14340
rect 5540 14288 5592 14340
rect 6920 14288 6972 14340
rect 26240 14399 26292 14408
rect 26240 14365 26249 14399
rect 26249 14365 26283 14399
rect 26283 14365 26292 14399
rect 26240 14356 26292 14365
rect 34520 14356 34572 14408
rect 3148 14220 3200 14272
rect 4436 14220 4488 14272
rect 15476 14288 15528 14340
rect 15568 14331 15620 14340
rect 15568 14297 15577 14331
rect 15577 14297 15611 14331
rect 15611 14297 15620 14331
rect 15568 14288 15620 14297
rect 16396 14220 16448 14272
rect 18420 14288 18472 14340
rect 20628 14288 20680 14340
rect 21272 14288 21324 14340
rect 22744 14288 22796 14340
rect 23848 14288 23900 14340
rect 18052 14220 18104 14272
rect 21640 14220 21692 14272
rect 22836 14220 22888 14272
rect 24676 14331 24728 14340
rect 24676 14297 24685 14331
rect 24685 14297 24719 14331
rect 24719 14297 24728 14331
rect 24676 14288 24728 14297
rect 26516 14331 26568 14340
rect 26516 14297 26525 14331
rect 26525 14297 26559 14331
rect 26559 14297 26568 14331
rect 26516 14288 26568 14297
rect 27804 14288 27856 14340
rect 30656 14288 30708 14340
rect 33324 14288 33376 14340
rect 33600 14288 33652 14340
rect 34336 14288 34388 14340
rect 26148 14263 26200 14272
rect 26148 14229 26157 14263
rect 26157 14229 26191 14263
rect 26191 14229 26200 14263
rect 26148 14220 26200 14229
rect 26332 14220 26384 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 1308 14016 1360 14068
rect 2964 14059 3016 14068
rect 2964 14025 2973 14059
rect 2973 14025 3007 14059
rect 3007 14025 3016 14059
rect 2964 14016 3016 14025
rect 5540 14016 5592 14068
rect 3056 13948 3108 14000
rect 4436 13991 4488 14000
rect 4436 13957 4445 13991
rect 4445 13957 4479 13991
rect 4479 13957 4488 13991
rect 4436 13948 4488 13957
rect 1676 13880 1728 13932
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 6920 13948 6972 14000
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 17960 14059 18012 14068
rect 17960 14025 17969 14059
rect 17969 14025 18003 14059
rect 18003 14025 18012 14059
rect 17960 14016 18012 14025
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 8852 13948 8904 14000
rect 15568 13948 15620 14000
rect 18420 13991 18472 14000
rect 18420 13957 18429 13991
rect 18429 13957 18463 13991
rect 18463 13957 18472 13991
rect 18420 13948 18472 13957
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9680 13880 9732 13932
rect 18972 13880 19024 13932
rect 21456 14016 21508 14068
rect 7932 13812 7984 13864
rect 14280 13855 14332 13864
rect 14280 13821 14289 13855
rect 14289 13821 14323 13855
rect 14323 13821 14332 13855
rect 14280 13812 14332 13821
rect 14556 13855 14608 13864
rect 14556 13821 14565 13855
rect 14565 13821 14599 13855
rect 14599 13821 14608 13855
rect 14556 13812 14608 13821
rect 18512 13812 18564 13864
rect 19984 13880 20036 13932
rect 21732 13880 21784 13932
rect 22008 13880 22060 13932
rect 22744 13948 22796 14000
rect 23020 13812 23072 13864
rect 23572 13923 23624 13932
rect 23572 13889 23581 13923
rect 23581 13889 23615 13923
rect 23615 13889 23624 13923
rect 23572 13880 23624 13889
rect 23940 13880 23992 13932
rect 26240 14016 26292 14068
rect 26516 14016 26568 14068
rect 28080 14016 28132 14068
rect 31668 14016 31720 14068
rect 32588 14016 32640 14068
rect 25504 13948 25556 14000
rect 26240 13880 26292 13932
rect 29644 13923 29696 13932
rect 29644 13889 29653 13923
rect 29653 13889 29687 13923
rect 29687 13889 29696 13923
rect 29644 13880 29696 13889
rect 32772 13948 32824 14000
rect 32864 13948 32916 14000
rect 32036 13880 32088 13932
rect 33416 13880 33468 13932
rect 33600 13880 33652 13932
rect 34336 13880 34388 13932
rect 24860 13812 24912 13864
rect 25964 13812 26016 13864
rect 18236 13744 18288 13796
rect 28908 13855 28960 13864
rect 28908 13821 28917 13855
rect 28917 13821 28951 13855
rect 28951 13821 28960 13855
rect 28908 13812 28960 13821
rect 29276 13812 29328 13864
rect 29552 13855 29604 13864
rect 29552 13821 29561 13855
rect 29561 13821 29595 13855
rect 29595 13821 29604 13855
rect 29552 13812 29604 13821
rect 30288 13855 30340 13864
rect 30288 13821 30297 13855
rect 30297 13821 30331 13855
rect 30331 13821 30340 13855
rect 30288 13812 30340 13821
rect 32404 13855 32456 13864
rect 32404 13821 32413 13855
rect 32413 13821 32447 13855
rect 32447 13821 32456 13855
rect 32404 13812 32456 13821
rect 27896 13744 27948 13796
rect 16028 13719 16080 13728
rect 16028 13685 16037 13719
rect 16037 13685 16071 13719
rect 16071 13685 16080 13719
rect 16028 13676 16080 13685
rect 33876 13676 33928 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 3148 13472 3200 13524
rect 22560 13515 22612 13524
rect 22560 13481 22569 13515
rect 22569 13481 22603 13515
rect 22603 13481 22612 13515
rect 22560 13472 22612 13481
rect 23572 13472 23624 13524
rect 32404 13515 32456 13524
rect 32404 13481 32413 13515
rect 32413 13481 32447 13515
rect 32447 13481 32456 13515
rect 32404 13472 32456 13481
rect 28080 13447 28132 13456
rect 28080 13413 28089 13447
rect 28089 13413 28123 13447
rect 28123 13413 28132 13447
rect 28080 13404 28132 13413
rect 1400 13336 1452 13388
rect 1860 13379 1912 13388
rect 1860 13345 1869 13379
rect 1869 13345 1903 13379
rect 1903 13345 1912 13379
rect 1860 13336 1912 13345
rect 3056 13336 3108 13388
rect 14556 13336 14608 13388
rect 16028 13336 16080 13388
rect 18604 13336 18656 13388
rect 21732 13336 21784 13388
rect 24676 13336 24728 13388
rect 26148 13336 26200 13388
rect 28908 13336 28960 13388
rect 34428 13336 34480 13388
rect 35348 13336 35400 13388
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 24860 13268 24912 13277
rect 24952 13268 25004 13320
rect 30104 13268 30156 13320
rect 30656 13268 30708 13320
rect 17040 13243 17092 13252
rect 17040 13209 17049 13243
rect 17049 13209 17083 13243
rect 17083 13209 17092 13243
rect 17040 13200 17092 13209
rect 16396 13132 16448 13184
rect 19984 13200 20036 13252
rect 21088 13243 21140 13252
rect 21088 13209 21097 13243
rect 21097 13209 21131 13243
rect 21131 13209 21140 13243
rect 21088 13200 21140 13209
rect 18512 13175 18564 13184
rect 18512 13141 18521 13175
rect 18521 13141 18555 13175
rect 18555 13141 18564 13175
rect 18512 13132 18564 13141
rect 21548 13200 21600 13252
rect 27712 13200 27764 13252
rect 29000 13200 29052 13252
rect 29552 13200 29604 13252
rect 30748 13132 30800 13184
rect 32128 13200 32180 13252
rect 33324 13200 33376 13252
rect 33876 13243 33928 13252
rect 33876 13209 33885 13243
rect 33885 13209 33919 13243
rect 33919 13209 33928 13243
rect 33876 13200 33928 13209
rect 34612 13200 34664 13252
rect 33600 13132 33652 13184
rect 33692 13132 33744 13184
rect 35440 13132 35492 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 16396 12860 16448 12912
rect 22008 12928 22060 12980
rect 14280 12792 14332 12844
rect 15200 12724 15252 12776
rect 15660 12724 15712 12776
rect 18052 12724 18104 12776
rect 19984 12860 20036 12912
rect 21732 12860 21784 12912
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 21088 12792 21140 12844
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 18604 12724 18656 12776
rect 19616 12724 19668 12776
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 24952 12971 25004 12980
rect 24952 12937 24961 12971
rect 24961 12937 24995 12971
rect 24995 12937 25004 12971
rect 24952 12928 25004 12937
rect 29000 12928 29052 12980
rect 29644 12928 29696 12980
rect 26240 12860 26292 12912
rect 29920 12860 29972 12912
rect 30288 12860 30340 12912
rect 24584 12792 24636 12844
rect 27344 12835 27396 12844
rect 27344 12801 27353 12835
rect 27353 12801 27387 12835
rect 27387 12801 27396 12835
rect 27344 12792 27396 12801
rect 30748 12835 30800 12844
rect 30748 12801 30757 12835
rect 30757 12801 30791 12835
rect 30791 12801 30800 12835
rect 30748 12792 30800 12801
rect 31116 12792 31168 12844
rect 34612 12928 34664 12980
rect 32128 12903 32180 12912
rect 32128 12869 32137 12903
rect 32137 12869 32171 12903
rect 32171 12869 32180 12903
rect 32128 12860 32180 12869
rect 32404 12860 32456 12912
rect 32588 12835 32640 12844
rect 32588 12801 32597 12835
rect 32597 12801 32631 12835
rect 32631 12801 32640 12835
rect 32588 12792 32640 12801
rect 33692 12903 33744 12912
rect 33692 12869 33701 12903
rect 33701 12869 33735 12903
rect 33735 12869 33744 12903
rect 33692 12860 33744 12869
rect 33784 12860 33836 12912
rect 20720 12724 20772 12733
rect 25504 12767 25556 12776
rect 25504 12733 25513 12767
rect 25513 12733 25547 12767
rect 25547 12733 25556 12767
rect 25504 12724 25556 12733
rect 26976 12724 27028 12776
rect 26056 12656 26108 12708
rect 30564 12724 30616 12776
rect 31024 12724 31076 12776
rect 33048 12724 33100 12776
rect 15844 12588 15896 12640
rect 28356 12588 28408 12640
rect 35348 12588 35400 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 29644 12384 29696 12436
rect 32772 12427 32824 12436
rect 32772 12393 32781 12427
rect 32781 12393 32815 12427
rect 32815 12393 32824 12427
rect 32772 12384 32824 12393
rect 10324 12248 10376 12300
rect 15200 12180 15252 12232
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 16212 12180 16264 12232
rect 18604 12180 18656 12232
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 19616 12180 19668 12189
rect 19800 12180 19852 12232
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20260 12180 20312 12189
rect 20628 12180 20680 12232
rect 20720 12223 20772 12232
rect 20720 12189 20729 12223
rect 20729 12189 20763 12223
rect 20763 12189 20772 12223
rect 20720 12180 20772 12189
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 23296 12248 23348 12300
rect 26056 12248 26108 12300
rect 28356 12291 28408 12300
rect 28356 12257 28365 12291
rect 28365 12257 28399 12291
rect 28399 12257 28408 12291
rect 28356 12248 28408 12257
rect 30564 12248 30616 12300
rect 31392 12248 31444 12300
rect 16028 12112 16080 12164
rect 16396 12112 16448 12164
rect 17960 12155 18012 12164
rect 17960 12121 17969 12155
rect 17969 12121 18003 12155
rect 18003 12121 18012 12155
rect 17960 12112 18012 12121
rect 21548 12112 21600 12164
rect 26608 12155 26660 12164
rect 26608 12121 26617 12155
rect 26617 12121 26651 12155
rect 26651 12121 26660 12155
rect 26608 12112 26660 12121
rect 17868 12044 17920 12096
rect 22928 12087 22980 12096
rect 22928 12053 22937 12087
rect 22937 12053 22971 12087
rect 22971 12053 22980 12087
rect 22928 12044 22980 12053
rect 23112 12044 23164 12096
rect 23848 12087 23900 12096
rect 23848 12053 23857 12087
rect 23857 12053 23891 12087
rect 23891 12053 23900 12087
rect 23848 12044 23900 12053
rect 25044 12044 25096 12096
rect 26332 12044 26384 12096
rect 27344 12044 27396 12096
rect 27436 12044 27488 12096
rect 28448 12112 28500 12164
rect 34520 12223 34572 12232
rect 34520 12189 34529 12223
rect 34529 12189 34563 12223
rect 34563 12189 34572 12223
rect 34520 12180 34572 12189
rect 34612 12180 34664 12232
rect 35348 12223 35400 12232
rect 35348 12189 35357 12223
rect 35357 12189 35391 12223
rect 35391 12189 35400 12223
rect 35348 12180 35400 12189
rect 30012 12112 30064 12164
rect 31024 12155 31076 12164
rect 31024 12121 31033 12155
rect 31033 12121 31067 12155
rect 31067 12121 31076 12155
rect 31024 12112 31076 12121
rect 33600 12112 33652 12164
rect 29000 12044 29052 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 16028 11840 16080 11892
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 23848 11840 23900 11892
rect 25504 11840 25556 11892
rect 27712 11840 27764 11892
rect 16396 11772 16448 11824
rect 17040 11772 17092 11824
rect 17868 11772 17920 11824
rect 18052 11704 18104 11756
rect 23112 11772 23164 11824
rect 24584 11772 24636 11824
rect 25964 11772 26016 11824
rect 26240 11772 26292 11824
rect 27436 11772 27488 11824
rect 29000 11840 29052 11892
rect 30012 11840 30064 11892
rect 28448 11772 28500 11824
rect 18512 11704 18564 11756
rect 19984 11704 20036 11756
rect 13728 11636 13780 11688
rect 16212 11636 16264 11688
rect 16488 11636 16540 11688
rect 18604 11679 18656 11688
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 19340 11636 19392 11688
rect 20720 11636 20772 11688
rect 21916 11636 21968 11688
rect 24400 11679 24452 11688
rect 24400 11645 24409 11679
rect 24409 11645 24443 11679
rect 24443 11645 24452 11679
rect 24400 11636 24452 11645
rect 24676 11679 24728 11688
rect 24676 11645 24685 11679
rect 24685 11645 24719 11679
rect 24719 11645 24728 11679
rect 24676 11636 24728 11645
rect 28080 11636 28132 11688
rect 32128 11704 32180 11756
rect 31208 11568 31260 11620
rect 31668 11679 31720 11688
rect 31668 11645 31677 11679
rect 31677 11645 31711 11679
rect 31711 11645 31720 11679
rect 31668 11636 31720 11645
rect 31760 11679 31812 11688
rect 31760 11645 31769 11679
rect 31769 11645 31803 11679
rect 31803 11645 31812 11679
rect 31760 11636 31812 11645
rect 20076 11500 20128 11552
rect 20260 11500 20312 11552
rect 25044 11500 25096 11552
rect 30840 11543 30892 11552
rect 30840 11509 30849 11543
rect 30849 11509 30883 11543
rect 30883 11509 30892 11543
rect 30840 11500 30892 11509
rect 31116 11543 31168 11552
rect 31116 11509 31125 11543
rect 31125 11509 31159 11543
rect 31159 11509 31168 11543
rect 31116 11500 31168 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 16212 11296 16264 11348
rect 16764 11228 16816 11280
rect 16120 11160 16172 11212
rect 21364 11296 21416 11348
rect 24676 11339 24728 11348
rect 24676 11305 24685 11339
rect 24685 11305 24719 11339
rect 24719 11305 24728 11339
rect 24676 11296 24728 11305
rect 31116 11296 31168 11348
rect 32128 11296 32180 11348
rect 23296 11228 23348 11280
rect 26976 11271 27028 11280
rect 20168 11160 20220 11212
rect 21272 11203 21324 11212
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 18604 11092 18656 11144
rect 22100 11092 22152 11144
rect 22284 11092 22336 11144
rect 22560 11135 22612 11144
rect 22560 11101 22569 11135
rect 22569 11101 22603 11135
rect 22603 11101 22612 11135
rect 22560 11092 22612 11101
rect 22928 11160 22980 11212
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 26976 11237 26985 11271
rect 26985 11237 27019 11271
rect 27019 11237 27028 11271
rect 26976 11228 27028 11237
rect 16396 11024 16448 11076
rect 17592 10956 17644 11008
rect 17868 10956 17920 11008
rect 19524 11067 19576 11076
rect 19524 11033 19533 11067
rect 19533 11033 19567 11067
rect 19567 11033 19576 11067
rect 19524 11024 19576 11033
rect 19984 11024 20036 11076
rect 25044 11135 25096 11144
rect 25044 11101 25053 11135
rect 25053 11101 25087 11135
rect 25087 11101 25096 11135
rect 25044 11092 25096 11101
rect 26240 11092 26292 11144
rect 22836 11024 22888 11076
rect 23204 11067 23256 11076
rect 23204 11033 23213 11067
rect 23213 11033 23247 11067
rect 23247 11033 23256 11067
rect 23204 11024 23256 11033
rect 23388 11024 23440 11076
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 18696 10956 18748 11008
rect 22192 10956 22244 11008
rect 25136 10999 25188 11008
rect 25136 10965 25145 10999
rect 25145 10965 25179 10999
rect 25179 10965 25188 10999
rect 25136 10956 25188 10965
rect 27712 11160 27764 11212
rect 28448 11160 28500 11212
rect 30380 11160 30432 11212
rect 31392 11203 31444 11212
rect 31392 11169 31401 11203
rect 31401 11169 31435 11203
rect 31435 11169 31444 11203
rect 31392 11160 31444 11169
rect 32680 11160 32732 11212
rect 33048 11160 33100 11212
rect 34704 11228 34756 11280
rect 35440 11160 35492 11212
rect 33968 11135 34020 11144
rect 33968 11101 33977 11135
rect 33977 11101 34011 11135
rect 34011 11101 34020 11135
rect 33968 11092 34020 11101
rect 29000 11024 29052 11076
rect 26608 10956 26660 11008
rect 31668 10956 31720 11008
rect 31852 10956 31904 11008
rect 33600 10956 33652 11008
rect 34244 10956 34296 11008
rect 34428 10999 34480 11008
rect 34428 10965 34437 10999
rect 34437 10965 34471 10999
rect 34471 10965 34480 10999
rect 34428 10956 34480 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 15384 10752 15436 10804
rect 16028 10795 16080 10804
rect 16028 10761 16037 10795
rect 16037 10761 16071 10795
rect 16071 10761 16080 10795
rect 16028 10752 16080 10761
rect 17592 10752 17644 10804
rect 18052 10752 18104 10804
rect 19064 10752 19116 10804
rect 23848 10752 23900 10804
rect 26332 10795 26384 10804
rect 26332 10761 26341 10795
rect 26341 10761 26375 10795
rect 26375 10761 26384 10795
rect 26332 10752 26384 10761
rect 30380 10795 30432 10804
rect 30380 10761 30395 10795
rect 30395 10761 30429 10795
rect 30429 10761 30432 10795
rect 30380 10752 30432 10761
rect 16396 10684 16448 10736
rect 17960 10684 18012 10736
rect 18420 10684 18472 10736
rect 22100 10684 22152 10736
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 16764 10616 16816 10668
rect 17408 10616 17460 10668
rect 16212 10591 16264 10600
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 17684 10548 17736 10600
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 21272 10616 21324 10668
rect 23664 10616 23716 10668
rect 18236 10548 18288 10600
rect 20812 10548 20864 10600
rect 21364 10591 21416 10600
rect 21364 10557 21373 10591
rect 21373 10557 21407 10591
rect 21407 10557 21416 10591
rect 21364 10548 21416 10557
rect 22284 10548 22336 10600
rect 23296 10480 23348 10532
rect 28632 10684 28684 10736
rect 30012 10684 30064 10736
rect 30840 10684 30892 10736
rect 31852 10727 31904 10736
rect 31852 10693 31861 10727
rect 31861 10693 31895 10727
rect 31895 10693 31904 10727
rect 31852 10684 31904 10693
rect 34428 10752 34480 10804
rect 33600 10684 33652 10736
rect 34244 10684 34296 10736
rect 25136 10659 25188 10668
rect 25136 10625 25145 10659
rect 25145 10625 25179 10659
rect 25179 10625 25188 10659
rect 25136 10616 25188 10625
rect 26148 10616 26200 10668
rect 26608 10616 26660 10668
rect 27988 10616 28040 10668
rect 25320 10548 25372 10600
rect 26056 10548 26108 10600
rect 26240 10591 26292 10600
rect 26240 10557 26249 10591
rect 26249 10557 26283 10591
rect 26283 10557 26292 10591
rect 26240 10548 26292 10557
rect 26976 10548 27028 10600
rect 28448 10591 28500 10600
rect 28448 10557 28457 10591
rect 28457 10557 28491 10591
rect 28491 10557 28500 10591
rect 28448 10548 28500 10557
rect 28724 10591 28776 10600
rect 28724 10557 28733 10591
rect 28733 10557 28767 10591
rect 28767 10557 28776 10591
rect 28724 10548 28776 10557
rect 17960 10412 18012 10464
rect 19064 10412 19116 10464
rect 20720 10455 20772 10464
rect 20720 10421 20729 10455
rect 20729 10421 20763 10455
rect 20763 10421 20772 10455
rect 20720 10412 20772 10421
rect 22928 10455 22980 10464
rect 22928 10421 22937 10455
rect 22937 10421 22971 10455
rect 22971 10421 22980 10455
rect 22928 10412 22980 10421
rect 26700 10480 26752 10532
rect 31484 10659 31536 10668
rect 31484 10625 31493 10659
rect 31493 10625 31527 10659
rect 31527 10625 31536 10659
rect 31484 10616 31536 10625
rect 31208 10591 31260 10600
rect 31208 10557 31217 10591
rect 31217 10557 31251 10591
rect 31251 10557 31260 10591
rect 31208 10548 31260 10557
rect 32496 10616 32548 10668
rect 32680 10659 32732 10668
rect 32680 10625 32689 10659
rect 32689 10625 32723 10659
rect 32723 10625 32732 10659
rect 32680 10616 32732 10625
rect 33416 10548 33468 10600
rect 34520 10591 34572 10600
rect 34520 10557 34529 10591
rect 34529 10557 34563 10591
rect 34563 10557 34572 10591
rect 34520 10548 34572 10557
rect 34796 10591 34848 10600
rect 34796 10557 34805 10591
rect 34805 10557 34839 10591
rect 34839 10557 34848 10591
rect 34796 10548 34848 10557
rect 32404 10480 32456 10532
rect 23940 10412 23992 10464
rect 24676 10412 24728 10464
rect 26792 10455 26844 10464
rect 26792 10421 26801 10455
rect 26801 10421 26835 10455
rect 26835 10421 26844 10455
rect 26792 10412 26844 10421
rect 30380 10412 30432 10464
rect 33968 10412 34020 10464
rect 34428 10455 34480 10464
rect 34428 10421 34437 10455
rect 34437 10421 34471 10455
rect 34471 10421 34480 10455
rect 34428 10412 34480 10421
rect 35348 10412 35400 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 17868 10251 17920 10260
rect 17868 10217 17877 10251
rect 17877 10217 17911 10251
rect 17911 10217 17920 10251
rect 17868 10208 17920 10217
rect 22192 10208 22244 10260
rect 22560 10208 22612 10260
rect 25136 10208 25188 10260
rect 28724 10208 28776 10260
rect 31760 10251 31812 10260
rect 31760 10217 31769 10251
rect 31769 10217 31803 10251
rect 31803 10217 31812 10251
rect 31760 10208 31812 10217
rect 31852 10208 31904 10260
rect 15936 10072 15988 10124
rect 18144 10072 18196 10124
rect 18236 10072 18288 10124
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 15476 10047 15528 10056
rect 15476 10013 15485 10047
rect 15485 10013 15519 10047
rect 15519 10013 15528 10047
rect 15476 10004 15528 10013
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 13912 9936 13964 9988
rect 16396 9936 16448 9988
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 19524 10072 19576 10124
rect 20076 10115 20128 10124
rect 20076 10081 20085 10115
rect 20085 10081 20119 10115
rect 20119 10081 20128 10115
rect 20076 10072 20128 10081
rect 21916 10072 21968 10124
rect 23572 10072 23624 10124
rect 24400 10115 24452 10124
rect 24400 10081 24409 10115
rect 24409 10081 24443 10115
rect 24443 10081 24452 10115
rect 24400 10072 24452 10081
rect 24676 10115 24728 10124
rect 24676 10081 24685 10115
rect 24685 10081 24719 10115
rect 24719 10081 24728 10115
rect 24676 10072 24728 10081
rect 19340 10047 19392 10056
rect 19340 10013 19349 10047
rect 19349 10013 19383 10047
rect 19383 10013 19392 10047
rect 19340 10004 19392 10013
rect 19800 10047 19852 10056
rect 19800 10013 19809 10047
rect 19809 10013 19843 10047
rect 19843 10013 19852 10047
rect 19800 10004 19852 10013
rect 20168 10004 20220 10056
rect 23020 10004 23072 10056
rect 23388 10004 23440 10056
rect 26976 10004 27028 10056
rect 29644 10047 29696 10056
rect 29644 10013 29653 10047
rect 29653 10013 29687 10047
rect 29687 10013 29696 10047
rect 29644 10004 29696 10013
rect 30196 10047 30248 10056
rect 30196 10013 30205 10047
rect 30205 10013 30239 10047
rect 30239 10013 30248 10047
rect 30196 10004 30248 10013
rect 31208 10072 31260 10124
rect 32496 10208 32548 10260
rect 33692 10208 33744 10260
rect 34612 10208 34664 10260
rect 34796 10208 34848 10260
rect 35440 10251 35492 10260
rect 35440 10217 35449 10251
rect 35449 10217 35483 10251
rect 35483 10217 35492 10251
rect 35440 10208 35492 10217
rect 32404 10140 32456 10192
rect 21548 9936 21600 9988
rect 25964 9936 26016 9988
rect 30380 9936 30432 9988
rect 31852 10047 31904 10056
rect 31852 10013 31861 10047
rect 31861 10013 31895 10047
rect 31895 10013 31904 10047
rect 31852 10004 31904 10013
rect 32128 10004 32180 10056
rect 32312 9936 32364 9988
rect 32496 10047 32548 10056
rect 32496 10013 32505 10047
rect 32505 10013 32539 10047
rect 32539 10013 32548 10047
rect 32496 10004 32548 10013
rect 32680 10047 32732 10056
rect 32680 10013 32689 10047
rect 32689 10013 32723 10047
rect 32723 10013 32732 10047
rect 32680 10004 32732 10013
rect 34428 10072 34480 10124
rect 34704 10047 34756 10056
rect 34704 10013 34713 10047
rect 34713 10013 34747 10047
rect 34747 10013 34756 10047
rect 34704 10004 34756 10013
rect 34796 10047 34848 10056
rect 34796 10013 34805 10047
rect 34805 10013 34839 10047
rect 34839 10013 34848 10047
rect 34796 10004 34848 10013
rect 34612 9936 34664 9988
rect 24952 9868 25004 9920
rect 29828 9911 29880 9920
rect 29828 9877 29837 9911
rect 29837 9877 29871 9911
rect 29871 9877 29880 9911
rect 29828 9868 29880 9877
rect 33784 9868 33836 9920
rect 34060 9911 34112 9920
rect 34060 9877 34069 9911
rect 34069 9877 34103 9911
rect 34103 9877 34112 9911
rect 34060 9868 34112 9877
rect 34244 9911 34296 9920
rect 34244 9877 34253 9911
rect 34253 9877 34287 9911
rect 34287 9877 34296 9911
rect 34244 9868 34296 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 15476 9664 15528 9716
rect 18420 9664 18472 9716
rect 13912 9639 13964 9648
rect 13912 9605 13921 9639
rect 13921 9605 13955 9639
rect 13955 9605 13964 9639
rect 13912 9596 13964 9605
rect 16396 9596 16448 9648
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 16488 9571 16540 9580
rect 16488 9537 16497 9571
rect 16497 9537 16531 9571
rect 16531 9537 16540 9571
rect 16488 9528 16540 9537
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 17868 9596 17920 9648
rect 18052 9596 18104 9648
rect 19984 9664 20036 9716
rect 20628 9664 20680 9716
rect 20720 9596 20772 9648
rect 26148 9707 26200 9716
rect 26148 9673 26157 9707
rect 26157 9673 26191 9707
rect 26191 9673 26200 9707
rect 26148 9664 26200 9673
rect 28632 9664 28684 9716
rect 23204 9596 23256 9648
rect 23388 9596 23440 9648
rect 24952 9596 25004 9648
rect 25136 9596 25188 9648
rect 26240 9596 26292 9648
rect 26700 9639 26752 9648
rect 26700 9605 26709 9639
rect 26709 9605 26743 9639
rect 26743 9605 26752 9639
rect 26700 9596 26752 9605
rect 26792 9596 26844 9648
rect 30196 9664 30248 9716
rect 32496 9664 32548 9716
rect 32680 9664 32732 9716
rect 32036 9596 32088 9648
rect 32312 9639 32364 9648
rect 32312 9605 32321 9639
rect 32321 9605 32355 9639
rect 32355 9605 32364 9639
rect 32312 9596 32364 9605
rect 33416 9639 33468 9648
rect 33416 9605 33425 9639
rect 33425 9605 33459 9639
rect 33459 9605 33468 9639
rect 33416 9596 33468 9605
rect 16120 9460 16172 9512
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 23572 9571 23624 9580
rect 23572 9537 23581 9571
rect 23581 9537 23615 9571
rect 23615 9537 23624 9571
rect 23572 9528 23624 9537
rect 28356 9528 28408 9580
rect 28724 9528 28776 9580
rect 29828 9571 29880 9580
rect 29828 9537 29837 9571
rect 29837 9537 29871 9571
rect 29871 9537 29880 9571
rect 29828 9528 29880 9537
rect 17868 9460 17920 9512
rect 17224 9392 17276 9444
rect 20076 9460 20128 9512
rect 22284 9460 22336 9512
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 26976 9503 27028 9512
rect 26976 9469 26985 9503
rect 26985 9469 27019 9503
rect 27019 9469 27028 9503
rect 26976 9460 27028 9469
rect 29276 9460 29328 9512
rect 29552 9460 29604 9512
rect 29736 9460 29788 9512
rect 30288 9571 30340 9580
rect 30288 9537 30297 9571
rect 30297 9537 30331 9571
rect 30331 9537 30340 9571
rect 30288 9528 30340 9537
rect 30748 9528 30800 9580
rect 31300 9528 31352 9580
rect 32680 9571 32732 9580
rect 32680 9537 32689 9571
rect 32689 9537 32723 9571
rect 32723 9537 32732 9571
rect 32680 9528 32732 9537
rect 32772 9528 32824 9580
rect 34612 9639 34664 9648
rect 34612 9605 34621 9639
rect 34621 9605 34655 9639
rect 34655 9605 34664 9639
rect 34612 9596 34664 9605
rect 33692 9571 33744 9580
rect 33692 9537 33701 9571
rect 33701 9537 33735 9571
rect 33735 9537 33744 9571
rect 33692 9528 33744 9537
rect 34244 9528 34296 9580
rect 35348 9528 35400 9580
rect 34796 9460 34848 9512
rect 33048 9392 33100 9444
rect 33784 9392 33836 9444
rect 28816 9367 28868 9376
rect 28816 9333 28825 9367
rect 28825 9333 28859 9367
rect 28859 9333 28868 9367
rect 28816 9324 28868 9333
rect 33140 9324 33192 9376
rect 34060 9324 34112 9376
rect 34244 9367 34296 9376
rect 34244 9333 34253 9367
rect 34253 9333 34287 9367
rect 34287 9333 34296 9367
rect 34244 9324 34296 9333
rect 34704 9324 34756 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 23664 9163 23716 9172
rect 23664 9129 23673 9163
rect 23673 9129 23707 9163
rect 23707 9129 23716 9163
rect 23664 9120 23716 9129
rect 24676 9120 24728 9172
rect 26700 9120 26752 9172
rect 28724 9163 28776 9172
rect 28724 9129 28733 9163
rect 28733 9129 28767 9163
rect 28767 9129 28776 9163
rect 28724 9120 28776 9129
rect 29644 9120 29696 9172
rect 31484 9120 31536 9172
rect 32772 9120 32824 9172
rect 34244 9120 34296 9172
rect 14280 8984 14332 9036
rect 16672 8984 16724 9036
rect 15292 8916 15344 8968
rect 15384 8959 15436 8968
rect 15384 8925 15393 8959
rect 15393 8925 15427 8959
rect 15427 8925 15436 8959
rect 15384 8916 15436 8925
rect 15476 8959 15528 8968
rect 15476 8925 15485 8959
rect 15485 8925 15519 8959
rect 15519 8925 15528 8959
rect 15476 8916 15528 8925
rect 18236 8916 18288 8968
rect 20444 8984 20496 9036
rect 21916 9027 21968 9036
rect 21916 8993 21925 9027
rect 21925 8993 21959 9027
rect 21959 8993 21968 9027
rect 21916 8984 21968 8993
rect 22928 8984 22980 9036
rect 23388 8984 23440 9036
rect 23572 8984 23624 9036
rect 14096 8848 14148 8900
rect 15936 8848 15988 8900
rect 16212 8848 16264 8900
rect 16396 8848 16448 8900
rect 18696 8916 18748 8968
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 23848 8916 23900 8968
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 26056 9027 26108 9036
rect 26056 8993 26065 9027
rect 26065 8993 26099 9027
rect 26099 8993 26108 9027
rect 26056 8984 26108 8993
rect 26976 9027 27028 9036
rect 26976 8993 26985 9027
rect 26985 8993 27019 9027
rect 27019 8993 27028 9027
rect 26976 8984 27028 8993
rect 28816 8984 28868 9036
rect 25596 8916 25648 8968
rect 26148 8916 26200 8968
rect 20628 8848 20680 8900
rect 21180 8891 21232 8900
rect 21180 8857 21189 8891
rect 21189 8857 21223 8891
rect 21223 8857 21232 8891
rect 21180 8848 21232 8857
rect 24584 8848 24636 8900
rect 25964 8823 26016 8832
rect 25964 8789 25973 8823
rect 25973 8789 26007 8823
rect 26007 8789 26016 8823
rect 25964 8780 26016 8789
rect 28356 8916 28408 8968
rect 30196 9052 30248 9104
rect 29552 8984 29604 9036
rect 31392 8984 31444 9036
rect 31668 9027 31720 9036
rect 31668 8993 31677 9027
rect 31677 8993 31711 9027
rect 31711 8993 31720 9027
rect 31668 8984 31720 8993
rect 33140 8984 33192 9036
rect 33416 8984 33468 9036
rect 34612 8984 34664 9036
rect 29460 8848 29512 8900
rect 30472 8916 30524 8968
rect 31208 8916 31260 8968
rect 32128 8916 32180 8968
rect 34060 8916 34112 8968
rect 34796 8916 34848 8968
rect 34980 8959 35032 8968
rect 34980 8925 34989 8959
rect 34989 8925 35023 8959
rect 35023 8925 35032 8959
rect 34980 8916 35032 8925
rect 30564 8848 30616 8900
rect 30656 8891 30708 8900
rect 30656 8857 30665 8891
rect 30665 8857 30699 8891
rect 30699 8857 30708 8891
rect 30656 8848 30708 8857
rect 27620 8780 27672 8832
rect 31300 8848 31352 8900
rect 30840 8823 30892 8832
rect 30840 8789 30849 8823
rect 30849 8789 30883 8823
rect 30883 8789 30892 8823
rect 30840 8780 30892 8789
rect 31576 8780 31628 8832
rect 33600 8848 33652 8900
rect 33416 8780 33468 8832
rect 35992 8848 36044 8900
rect 36452 8848 36504 8900
rect 34244 8780 34296 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 15476 8576 15528 8628
rect 16212 8576 16264 8628
rect 18696 8576 18748 8628
rect 19800 8576 19852 8628
rect 27988 8576 28040 8628
rect 14096 8551 14148 8560
rect 14096 8517 14105 8551
rect 14105 8517 14139 8551
rect 14139 8517 14148 8551
rect 14096 8508 14148 8517
rect 15660 8508 15712 8560
rect 16396 8508 16448 8560
rect 16488 8508 16540 8560
rect 23020 8551 23072 8560
rect 23020 8517 23029 8551
rect 23029 8517 23063 8551
rect 23063 8517 23072 8551
rect 23020 8508 23072 8517
rect 24032 8508 24084 8560
rect 26700 8508 26752 8560
rect 27620 8551 27672 8560
rect 27620 8517 27629 8551
rect 27629 8517 27663 8551
rect 27663 8517 27672 8551
rect 27620 8508 27672 8517
rect 33692 8576 33744 8628
rect 28724 8508 28776 8560
rect 29736 8508 29788 8560
rect 31208 8508 31260 8560
rect 31668 8508 31720 8560
rect 18604 8440 18656 8492
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 20444 8483 20496 8492
rect 20444 8449 20453 8483
rect 20453 8449 20487 8483
rect 20487 8449 20496 8483
rect 20444 8440 20496 8449
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 16672 8372 16724 8424
rect 18788 8372 18840 8424
rect 19800 8372 19852 8424
rect 21180 8483 21232 8492
rect 21180 8449 21189 8483
rect 21189 8449 21223 8483
rect 21223 8449 21232 8483
rect 21180 8440 21232 8449
rect 23756 8483 23808 8492
rect 23756 8449 23765 8483
rect 23765 8449 23799 8483
rect 23799 8449 23808 8483
rect 23756 8440 23808 8449
rect 23848 8440 23900 8492
rect 27896 8440 27948 8492
rect 32680 8508 32732 8560
rect 34244 8508 34296 8560
rect 34980 8576 35032 8628
rect 22100 8372 22152 8424
rect 23572 8372 23624 8424
rect 24032 8372 24084 8424
rect 27528 8372 27580 8424
rect 28356 8372 28408 8424
rect 18328 8304 18380 8356
rect 20812 8304 20864 8356
rect 26240 8304 26292 8356
rect 27712 8304 27764 8356
rect 14280 8236 14332 8288
rect 27988 8236 28040 8288
rect 29460 8372 29512 8424
rect 30196 8372 30248 8424
rect 30840 8372 30892 8424
rect 31300 8347 31352 8356
rect 31300 8313 31309 8347
rect 31309 8313 31343 8347
rect 31343 8313 31352 8347
rect 31300 8304 31352 8313
rect 31392 8347 31444 8356
rect 31392 8313 31401 8347
rect 31401 8313 31435 8347
rect 31435 8313 31444 8347
rect 31392 8304 31444 8313
rect 32128 8372 32180 8424
rect 32496 8440 32548 8492
rect 33416 8483 33468 8492
rect 33416 8449 33425 8483
rect 33425 8449 33459 8483
rect 33459 8449 33468 8483
rect 33416 8440 33468 8449
rect 33508 8440 33560 8492
rect 29920 8236 29972 8288
rect 32496 8236 32548 8288
rect 33048 8304 33100 8356
rect 33692 8236 33744 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 18328 8032 18380 8084
rect 25964 8032 26016 8084
rect 34612 8032 34664 8084
rect 14280 7939 14332 7948
rect 14280 7905 14289 7939
rect 14289 7905 14323 7939
rect 14323 7905 14332 7939
rect 14280 7896 14332 7905
rect 18788 7939 18840 7948
rect 18788 7905 18797 7939
rect 18797 7905 18831 7939
rect 18831 7905 18840 7939
rect 18788 7896 18840 7905
rect 21456 7939 21508 7948
rect 21456 7905 21465 7939
rect 21465 7905 21499 7939
rect 21499 7905 21508 7939
rect 21456 7896 21508 7905
rect 23664 7896 23716 7948
rect 23940 7939 23992 7948
rect 23940 7905 23949 7939
rect 23949 7905 23983 7939
rect 23983 7905 23992 7939
rect 23940 7896 23992 7905
rect 24124 7896 24176 7948
rect 25136 7896 25188 7948
rect 25688 7896 25740 7948
rect 27528 7896 27580 7948
rect 27620 7896 27672 7948
rect 30196 7939 30248 7948
rect 30196 7905 30205 7939
rect 30205 7905 30239 7939
rect 30239 7905 30248 7939
rect 30196 7896 30248 7905
rect 30656 7939 30708 7948
rect 30656 7905 30665 7939
rect 30665 7905 30699 7939
rect 30699 7905 30708 7939
rect 30656 7896 30708 7905
rect 15660 7828 15712 7880
rect 14556 7803 14608 7812
rect 14556 7769 14565 7803
rect 14565 7769 14599 7803
rect 14599 7769 14608 7803
rect 14556 7760 14608 7769
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 23296 7828 23348 7880
rect 23388 7828 23440 7880
rect 29920 7871 29972 7880
rect 29920 7837 29929 7871
rect 29929 7837 29963 7871
rect 29963 7837 29972 7871
rect 29920 7828 29972 7837
rect 31852 7828 31904 7880
rect 34060 7871 34112 7880
rect 34060 7837 34069 7871
rect 34069 7837 34103 7871
rect 34103 7837 34112 7871
rect 35992 7896 36044 7948
rect 34060 7828 34112 7837
rect 17408 7760 17460 7812
rect 20628 7760 20680 7812
rect 23756 7803 23808 7812
rect 16028 7735 16080 7744
rect 16028 7701 16037 7735
rect 16037 7701 16071 7735
rect 16071 7701 16080 7735
rect 16028 7692 16080 7701
rect 20536 7692 20588 7744
rect 22192 7692 22244 7744
rect 23756 7769 23765 7803
rect 23765 7769 23799 7803
rect 23799 7769 23808 7803
rect 23756 7760 23808 7769
rect 24952 7760 25004 7812
rect 25136 7760 25188 7812
rect 27528 7760 27580 7812
rect 27988 7803 28040 7812
rect 27988 7769 27997 7803
rect 27997 7769 28031 7803
rect 28031 7769 28040 7803
rect 27988 7760 28040 7769
rect 30564 7760 30616 7812
rect 32956 7803 33008 7812
rect 32956 7769 32965 7803
rect 32965 7769 32999 7803
rect 32999 7769 33008 7803
rect 32956 7760 33008 7769
rect 33324 7760 33376 7812
rect 35440 7828 35492 7880
rect 36176 7803 36228 7812
rect 36176 7769 36185 7803
rect 36185 7769 36219 7803
rect 36219 7769 36228 7803
rect 36176 7760 36228 7769
rect 27896 7692 27948 7744
rect 28448 7692 28500 7744
rect 30196 7692 30248 7744
rect 34336 7692 34388 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 14556 7420 14608 7472
rect 15200 7352 15252 7404
rect 18972 7488 19024 7540
rect 23572 7488 23624 7540
rect 25596 7488 25648 7540
rect 27896 7488 27948 7540
rect 30104 7488 30156 7540
rect 17408 7420 17460 7472
rect 20628 7420 20680 7472
rect 23296 7420 23348 7472
rect 24032 7420 24084 7472
rect 24584 7463 24636 7472
rect 24584 7429 24593 7463
rect 24593 7429 24627 7463
rect 24627 7429 24636 7463
rect 24584 7420 24636 7429
rect 25136 7420 25188 7472
rect 27804 7420 27856 7472
rect 28448 7463 28500 7472
rect 28448 7429 28457 7463
rect 28457 7429 28491 7463
rect 28491 7429 28500 7463
rect 28448 7420 28500 7429
rect 29736 7420 29788 7472
rect 31024 7420 31076 7472
rect 31852 7463 31904 7472
rect 31852 7429 31861 7463
rect 31861 7429 31895 7463
rect 31895 7429 31904 7463
rect 31852 7420 31904 7429
rect 33692 7420 33744 7472
rect 34060 7420 34112 7472
rect 35440 7420 35492 7472
rect 15568 7352 15620 7404
rect 16028 7352 16080 7404
rect 21456 7352 21508 7404
rect 27620 7352 27672 7404
rect 28172 7395 28224 7404
rect 28172 7361 28181 7395
rect 28181 7361 28215 7395
rect 28215 7361 28224 7395
rect 28172 7352 28224 7361
rect 30288 7395 30340 7404
rect 30288 7361 30297 7395
rect 30297 7361 30331 7395
rect 30331 7361 30340 7395
rect 30288 7352 30340 7361
rect 30564 7352 30616 7404
rect 32128 7395 32180 7404
rect 32128 7361 32137 7395
rect 32137 7361 32171 7395
rect 32171 7361 32180 7395
rect 32128 7352 32180 7361
rect 34336 7395 34388 7404
rect 34336 7361 34345 7395
rect 34345 7361 34379 7395
rect 34379 7361 34388 7395
rect 34336 7352 34388 7361
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 18512 7284 18564 7336
rect 20904 7327 20956 7336
rect 20904 7293 20913 7327
rect 20913 7293 20947 7327
rect 20947 7293 20956 7327
rect 20904 7284 20956 7293
rect 22100 7284 22152 7336
rect 18604 7148 18656 7200
rect 19248 7148 19300 7200
rect 20444 7148 20496 7200
rect 23388 7148 23440 7200
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 30012 7327 30064 7336
rect 30012 7293 30021 7327
rect 30021 7293 30055 7327
rect 30055 7293 30064 7327
rect 30012 7284 30064 7293
rect 31760 7284 31812 7336
rect 26976 7191 27028 7200
rect 26976 7157 26985 7191
rect 26985 7157 27019 7191
rect 27019 7157 27028 7191
rect 26976 7148 27028 7157
rect 34520 7216 34572 7268
rect 32496 7148 32548 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 22192 6987 22244 6996
rect 22192 6953 22201 6987
rect 22201 6953 22235 6987
rect 22235 6953 22244 6987
rect 22192 6944 22244 6953
rect 26976 6944 27028 6996
rect 27804 6987 27856 6996
rect 27804 6953 27813 6987
rect 27813 6953 27847 6987
rect 27847 6953 27856 6987
rect 27804 6944 27856 6953
rect 30288 6876 30340 6928
rect 16028 6808 16080 6860
rect 16672 6851 16724 6860
rect 16672 6817 16681 6851
rect 16681 6817 16715 6851
rect 16715 6817 16724 6851
rect 16672 6808 16724 6817
rect 19064 6808 19116 6860
rect 20444 6808 20496 6860
rect 14832 6672 14884 6724
rect 15752 6740 15804 6792
rect 18972 6740 19024 6792
rect 21272 6740 21324 6792
rect 21548 6783 21600 6792
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 21732 6783 21784 6792
rect 21732 6749 21741 6783
rect 21741 6749 21775 6783
rect 21775 6749 21784 6783
rect 21732 6740 21784 6749
rect 21824 6783 21876 6792
rect 21824 6749 21833 6783
rect 21833 6749 21867 6783
rect 21867 6749 21876 6783
rect 21824 6740 21876 6749
rect 22468 6808 22520 6860
rect 24124 6808 24176 6860
rect 24952 6851 25004 6860
rect 24952 6817 24961 6851
rect 24961 6817 24995 6851
rect 24995 6817 25004 6851
rect 24952 6808 25004 6817
rect 25964 6808 26016 6860
rect 28172 6808 28224 6860
rect 30012 6808 30064 6860
rect 22928 6740 22980 6792
rect 25320 6740 25372 6792
rect 25596 6783 25648 6792
rect 25596 6749 25605 6783
rect 25605 6749 25639 6783
rect 25639 6749 25648 6783
rect 25596 6740 25648 6749
rect 26056 6783 26108 6792
rect 26056 6749 26065 6783
rect 26065 6749 26099 6783
rect 26099 6749 26108 6783
rect 26056 6740 26108 6749
rect 27344 6740 27396 6792
rect 30656 6808 30708 6860
rect 34152 6919 34204 6928
rect 34152 6885 34161 6919
rect 34161 6885 34195 6919
rect 34195 6885 34204 6919
rect 34152 6876 34204 6885
rect 16948 6715 17000 6724
rect 16948 6681 16957 6715
rect 16957 6681 16991 6715
rect 16991 6681 17000 6715
rect 16948 6672 17000 6681
rect 17408 6672 17460 6724
rect 19524 6672 19576 6724
rect 17868 6604 17920 6656
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 20536 6604 20588 6656
rect 30380 6672 30432 6724
rect 30564 6672 30616 6724
rect 29736 6604 29788 6656
rect 31760 6808 31812 6860
rect 32128 6808 32180 6860
rect 33048 6808 33100 6860
rect 32220 6740 32272 6792
rect 33692 6740 33744 6792
rect 34336 6740 34388 6792
rect 32588 6715 32640 6724
rect 32588 6681 32597 6715
rect 32597 6681 32631 6715
rect 32631 6681 32640 6715
rect 32588 6672 32640 6681
rect 34060 6672 34112 6724
rect 33324 6604 33376 6656
rect 34612 6604 34664 6656
rect 34796 6647 34848 6656
rect 34796 6613 34805 6647
rect 34805 6613 34839 6647
rect 34839 6613 34848 6647
rect 34796 6604 34848 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 14280 6400 14332 6452
rect 14096 6332 14148 6384
rect 15660 6332 15712 6384
rect 16948 6332 17000 6384
rect 18144 6332 18196 6384
rect 18972 6400 19024 6452
rect 21548 6400 21600 6452
rect 14832 6196 14884 6248
rect 18420 6264 18472 6316
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 20904 6332 20956 6384
rect 18328 6196 18380 6248
rect 17868 6128 17920 6180
rect 19248 6307 19300 6316
rect 19248 6273 19257 6307
rect 19257 6273 19291 6307
rect 19291 6273 19300 6307
rect 19248 6264 19300 6273
rect 20444 6307 20496 6316
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 22928 6332 22980 6384
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 24676 6264 24728 6316
rect 25688 6400 25740 6452
rect 29736 6400 29788 6452
rect 28540 6332 28592 6384
rect 30380 6332 30432 6384
rect 32588 6332 32640 6384
rect 33600 6332 33652 6384
rect 33784 6332 33836 6384
rect 32220 6264 32272 6316
rect 21824 6196 21876 6248
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 22468 6239 22520 6248
rect 22468 6205 22477 6239
rect 22477 6205 22511 6239
rect 22511 6205 22520 6239
rect 22468 6196 22520 6205
rect 23112 6196 23164 6248
rect 23388 6239 23440 6248
rect 23388 6205 23397 6239
rect 23397 6205 23431 6239
rect 23431 6205 23440 6239
rect 23388 6196 23440 6205
rect 24400 6196 24452 6248
rect 27436 6196 27488 6248
rect 27712 6196 27764 6248
rect 28080 6196 28132 6248
rect 28172 6239 28224 6248
rect 28172 6205 28181 6239
rect 28181 6205 28215 6239
rect 28215 6205 28224 6239
rect 28172 6196 28224 6205
rect 30104 6196 30156 6248
rect 22100 6128 22152 6180
rect 29460 6128 29512 6180
rect 30472 6239 30524 6248
rect 30472 6205 30481 6239
rect 30481 6205 30515 6239
rect 30515 6205 30524 6239
rect 30472 6196 30524 6205
rect 32680 6239 32732 6248
rect 32680 6205 32689 6239
rect 32689 6205 32723 6239
rect 32723 6205 32732 6239
rect 32680 6196 32732 6205
rect 34152 6332 34204 6384
rect 34336 6332 34388 6384
rect 33048 6196 33100 6248
rect 34796 6196 34848 6248
rect 15384 6060 15436 6112
rect 15752 6060 15804 6112
rect 23296 6060 23348 6112
rect 25136 6103 25188 6112
rect 25136 6069 25145 6103
rect 25145 6069 25179 6103
rect 25179 6069 25188 6103
rect 25136 6060 25188 6069
rect 27160 6103 27212 6112
rect 27160 6069 27169 6103
rect 27169 6069 27203 6103
rect 27203 6069 27212 6103
rect 27160 6060 27212 6069
rect 29920 6103 29972 6112
rect 29920 6069 29929 6103
rect 29929 6069 29963 6103
rect 29963 6069 29972 6103
rect 29920 6060 29972 6069
rect 36728 6171 36780 6180
rect 36728 6137 36737 6171
rect 36737 6137 36771 6171
rect 36771 6137 36780 6171
rect 36728 6128 36780 6137
rect 32128 6060 32180 6112
rect 32312 6060 32364 6112
rect 33692 6103 33744 6112
rect 33692 6069 33701 6103
rect 33701 6069 33735 6103
rect 33735 6069 33744 6103
rect 33692 6060 33744 6069
rect 33784 6060 33836 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 21824 5856 21876 5908
rect 30472 5856 30524 5908
rect 33600 5899 33652 5908
rect 33600 5865 33609 5899
rect 33609 5865 33643 5899
rect 33643 5865 33652 5899
rect 33600 5856 33652 5865
rect 33692 5856 33744 5908
rect 34612 5856 34664 5908
rect 35348 5856 35400 5908
rect 27436 5831 27488 5840
rect 27436 5797 27445 5831
rect 27445 5797 27479 5831
rect 27479 5797 27488 5831
rect 27436 5788 27488 5797
rect 15844 5720 15896 5772
rect 14372 5627 14424 5636
rect 14372 5593 14381 5627
rect 14381 5593 14415 5627
rect 14415 5593 14424 5627
rect 14372 5584 14424 5593
rect 15384 5652 15436 5704
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16580 5763 16632 5772
rect 16580 5729 16589 5763
rect 16589 5729 16623 5763
rect 16623 5729 16632 5763
rect 16580 5720 16632 5729
rect 19064 5720 19116 5772
rect 19524 5763 19576 5772
rect 19524 5729 19533 5763
rect 19533 5729 19567 5763
rect 19567 5729 19576 5763
rect 19524 5720 19576 5729
rect 22284 5720 22336 5772
rect 24400 5763 24452 5772
rect 24400 5729 24409 5763
rect 24409 5729 24443 5763
rect 24443 5729 24452 5763
rect 24400 5720 24452 5729
rect 25136 5763 25188 5772
rect 25136 5729 25145 5763
rect 25145 5729 25179 5763
rect 25179 5729 25188 5763
rect 25136 5720 25188 5729
rect 15200 5584 15252 5636
rect 15568 5584 15620 5636
rect 23112 5695 23164 5704
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 16764 5584 16816 5636
rect 16856 5627 16908 5636
rect 16856 5593 16865 5627
rect 16865 5593 16899 5627
rect 16899 5593 16908 5627
rect 16856 5584 16908 5593
rect 17408 5584 17460 5636
rect 20536 5584 20588 5636
rect 22284 5584 22336 5636
rect 18328 5559 18380 5568
rect 18328 5525 18337 5559
rect 18337 5525 18371 5559
rect 18371 5525 18380 5559
rect 18328 5516 18380 5525
rect 21548 5516 21600 5568
rect 23848 5695 23900 5704
rect 23848 5661 23857 5695
rect 23857 5661 23891 5695
rect 23891 5661 23900 5695
rect 23848 5652 23900 5661
rect 24860 5695 24912 5704
rect 24860 5661 24869 5695
rect 24869 5661 24903 5695
rect 24903 5661 24912 5695
rect 24860 5652 24912 5661
rect 24952 5652 25004 5704
rect 25412 5652 25464 5704
rect 26056 5720 26108 5772
rect 27344 5652 27396 5704
rect 33784 5788 33836 5840
rect 27804 5720 27856 5772
rect 28080 5720 28132 5772
rect 30288 5720 30340 5772
rect 32312 5720 32364 5772
rect 33140 5763 33192 5772
rect 33140 5729 33149 5763
rect 33149 5729 33183 5763
rect 33183 5729 33192 5763
rect 33140 5720 33192 5729
rect 28540 5695 28592 5704
rect 28540 5661 28549 5695
rect 28549 5661 28583 5695
rect 28583 5661 28592 5695
rect 28540 5652 28592 5661
rect 31116 5652 31168 5704
rect 33232 5695 33284 5704
rect 33232 5661 33241 5695
rect 33241 5661 33275 5695
rect 33275 5661 33284 5695
rect 33232 5652 33284 5661
rect 33416 5695 33468 5704
rect 33416 5661 33425 5695
rect 33425 5661 33459 5695
rect 33459 5661 33468 5695
rect 33416 5652 33468 5661
rect 29828 5584 29880 5636
rect 29552 5516 29604 5568
rect 33324 5584 33376 5636
rect 33784 5652 33836 5704
rect 34520 5584 34572 5636
rect 35072 5584 35124 5636
rect 36176 5516 36228 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 14372 5287 14424 5296
rect 14372 5253 14381 5287
rect 14381 5253 14415 5287
rect 14415 5253 14424 5287
rect 14372 5244 14424 5253
rect 15660 5244 15712 5296
rect 16856 5244 16908 5296
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 18144 5244 18196 5296
rect 16764 5108 16816 5160
rect 18328 5176 18380 5228
rect 23112 5312 23164 5364
rect 23296 5287 23348 5296
rect 23296 5253 23305 5287
rect 23305 5253 23339 5287
rect 23339 5253 23348 5287
rect 23296 5244 23348 5253
rect 20536 5176 20588 5228
rect 20812 5108 20864 5160
rect 22100 5108 22152 5160
rect 22284 5176 22336 5228
rect 24676 5244 24728 5296
rect 28172 5312 28224 5364
rect 28540 5312 28592 5364
rect 25412 5219 25464 5228
rect 25412 5185 25421 5219
rect 25421 5185 25455 5219
rect 25455 5185 25464 5219
rect 25412 5176 25464 5185
rect 27160 5244 27212 5296
rect 29736 5244 29788 5296
rect 30012 5312 30064 5364
rect 30104 5312 30156 5364
rect 32312 5355 32364 5364
rect 32312 5321 32339 5355
rect 32339 5321 32364 5355
rect 32312 5312 32364 5321
rect 29920 5287 29972 5296
rect 29920 5253 29929 5287
rect 29929 5253 29963 5287
rect 29963 5253 29972 5287
rect 29920 5244 29972 5253
rect 29552 5219 29604 5228
rect 29552 5185 29561 5219
rect 29561 5185 29595 5219
rect 29595 5185 29604 5219
rect 29552 5176 29604 5185
rect 24400 5108 24452 5160
rect 30196 5176 30248 5228
rect 30380 5287 30432 5296
rect 30380 5253 30389 5287
rect 30389 5253 30423 5287
rect 30423 5253 30432 5287
rect 30380 5244 30432 5253
rect 21732 5040 21784 5092
rect 23848 4972 23900 5024
rect 24492 4972 24544 5024
rect 24952 4972 25004 5024
rect 30840 5219 30892 5228
rect 30840 5185 30849 5219
rect 30849 5185 30883 5219
rect 30883 5185 30892 5219
rect 30840 5176 30892 5185
rect 31024 5219 31076 5228
rect 31024 5185 31033 5219
rect 31033 5185 31067 5219
rect 31067 5185 31076 5219
rect 31024 5176 31076 5185
rect 31116 5219 31168 5228
rect 31116 5185 31125 5219
rect 31125 5185 31159 5219
rect 31159 5185 31168 5219
rect 31116 5176 31168 5185
rect 32496 5287 32548 5296
rect 32496 5253 32505 5287
rect 32505 5253 32539 5287
rect 32539 5253 32548 5287
rect 32496 5244 32548 5253
rect 33324 5244 33376 5296
rect 33140 5219 33192 5228
rect 33140 5185 33149 5219
rect 33149 5185 33183 5219
rect 33183 5185 33192 5219
rect 33140 5176 33192 5185
rect 33416 5219 33468 5228
rect 33416 5185 33425 5219
rect 33425 5185 33459 5219
rect 33459 5185 33468 5219
rect 33416 5176 33468 5185
rect 35072 5287 35124 5296
rect 35072 5253 35081 5287
rect 35081 5253 35115 5287
rect 35115 5253 35124 5287
rect 35072 5244 35124 5253
rect 34704 5219 34756 5228
rect 34704 5185 34713 5219
rect 34713 5185 34747 5219
rect 34747 5185 34756 5219
rect 34704 5176 34756 5185
rect 34888 5219 34940 5228
rect 34888 5185 34897 5219
rect 34897 5185 34931 5219
rect 34931 5185 34940 5219
rect 34888 5176 34940 5185
rect 34060 5151 34112 5160
rect 34060 5117 34069 5151
rect 34069 5117 34103 5151
rect 34103 5117 34112 5151
rect 34060 5108 34112 5117
rect 34428 5108 34480 5160
rect 30472 5040 30524 5092
rect 34336 5040 34388 5092
rect 30656 4972 30708 5024
rect 32312 5015 32364 5024
rect 32312 4981 32321 5015
rect 32321 4981 32355 5015
rect 32355 4981 32364 5015
rect 32312 4972 32364 4981
rect 33232 4972 33284 5024
rect 34796 4972 34848 5024
rect 35532 4972 35584 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 16764 4768 16816 4820
rect 14096 4632 14148 4684
rect 15568 4675 15620 4684
rect 15568 4641 15577 4675
rect 15577 4641 15611 4675
rect 15611 4641 15620 4675
rect 15568 4632 15620 4641
rect 20812 4675 20864 4684
rect 20812 4641 20821 4675
rect 20821 4641 20855 4675
rect 20855 4641 20864 4675
rect 20812 4632 20864 4641
rect 21548 4700 21600 4752
rect 30380 4700 30432 4752
rect 22100 4632 22152 4684
rect 24400 4675 24452 4684
rect 24400 4641 24409 4675
rect 24409 4641 24443 4675
rect 24443 4641 24452 4675
rect 24400 4632 24452 4641
rect 24492 4632 24544 4684
rect 21732 4564 21784 4616
rect 15660 4496 15712 4548
rect 25044 4607 25096 4616
rect 25044 4573 25053 4607
rect 25053 4573 25087 4607
rect 25087 4573 25096 4607
rect 25044 4564 25096 4573
rect 30840 4632 30892 4684
rect 32312 4700 32364 4752
rect 34704 4700 34756 4752
rect 31944 4632 31996 4684
rect 25320 4496 25372 4548
rect 29460 4496 29512 4548
rect 30472 4564 30524 4616
rect 32036 4564 32088 4616
rect 31024 4496 31076 4548
rect 33140 4564 33192 4616
rect 33232 4607 33284 4616
rect 33232 4573 33241 4607
rect 33241 4573 33275 4607
rect 33275 4573 33284 4607
rect 33232 4564 33284 4573
rect 33324 4564 33376 4616
rect 34428 4632 34480 4684
rect 33692 4564 33744 4616
rect 33416 4496 33468 4548
rect 34336 4496 34388 4548
rect 34888 4607 34940 4616
rect 34888 4573 34897 4607
rect 34897 4573 34931 4607
rect 34931 4573 34940 4607
rect 34888 4564 34940 4573
rect 35348 4564 35400 4616
rect 35532 4539 35584 4548
rect 35532 4505 35559 4539
rect 35559 4505 35584 4539
rect 35532 4496 35584 4505
rect 30380 4428 30432 4480
rect 31300 4428 31352 4480
rect 32312 4471 32364 4480
rect 32312 4437 32321 4471
rect 32321 4437 32355 4471
rect 32355 4437 32364 4471
rect 32312 4428 32364 4437
rect 32496 4471 32548 4480
rect 32496 4437 32505 4471
rect 32505 4437 32539 4471
rect 32539 4437 32548 4471
rect 32496 4428 32548 4437
rect 35348 4471 35400 4480
rect 35348 4437 35357 4471
rect 35357 4437 35391 4471
rect 35391 4437 35400 4471
rect 35348 4428 35400 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 30380 4267 30432 4276
rect 30380 4233 30389 4267
rect 30389 4233 30423 4267
rect 30423 4233 30432 4267
rect 30380 4224 30432 4233
rect 31760 4224 31812 4276
rect 31944 4224 31996 4276
rect 32312 4224 32364 4276
rect 32404 4224 32456 4276
rect 30288 4156 30340 4208
rect 28172 4088 28224 4140
rect 31300 4199 31352 4208
rect 31300 4165 31309 4199
rect 31309 4165 31343 4199
rect 31343 4165 31352 4199
rect 31300 4156 31352 4165
rect 32036 4156 32088 4208
rect 33324 4267 33376 4276
rect 33324 4233 33333 4267
rect 33333 4233 33367 4267
rect 33367 4233 33376 4267
rect 33324 4224 33376 4233
rect 33416 4224 33468 4276
rect 33692 4156 33744 4208
rect 35348 4156 35400 4208
rect 30748 4088 30800 4140
rect 29460 4020 29512 4072
rect 32496 4088 32548 4140
rect 31852 4020 31904 4072
rect 32404 4020 32456 4072
rect 32680 4063 32732 4072
rect 32680 4029 32689 4063
rect 32689 4029 32723 4063
rect 32723 4029 32732 4063
rect 33968 4088 34020 4140
rect 32680 4020 32732 4029
rect 33048 4020 33100 4072
rect 30472 3884 30524 3936
rect 33600 3884 33652 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 31760 3680 31812 3732
rect 32956 3680 33008 3732
rect 33600 3612 33652 3664
rect 30656 3544 30708 3596
rect 31852 3544 31904 3596
rect 30012 3519 30064 3528
rect 30012 3485 30021 3519
rect 30021 3485 30055 3519
rect 30055 3485 30064 3519
rect 30012 3476 30064 3485
rect 33232 3544 33284 3596
rect 30932 3408 30984 3460
rect 32956 3476 33008 3528
rect 33692 3408 33744 3460
rect 34704 3408 34756 3460
rect 32404 3340 32456 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 34704 3136 34756 3188
rect 30472 3111 30524 3120
rect 30472 3077 30481 3111
rect 30481 3077 30515 3111
rect 30515 3077 30524 3111
rect 30472 3068 30524 3077
rect 30932 3068 30984 3120
rect 32404 3111 32456 3120
rect 32404 3077 32413 3111
rect 32413 3077 32447 3111
rect 32447 3077 32456 3111
rect 32404 3068 32456 3077
rect 33968 3068 34020 3120
rect 30012 2932 30064 2984
rect 32036 2932 32088 2984
rect 33048 2932 33100 2984
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 24952 2592 25004 2644
rect 23204 2388 23256 2440
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 25134 39658 25190 40352
rect 29642 39658 29698 40352
rect 30930 39658 30986 40352
rect 25134 39630 25268 39658
rect 25134 39552 25190 39630
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 25240 37874 25268 39630
rect 29642 39630 29776 39658
rect 29642 39552 29698 39630
rect 29748 37874 29776 39630
rect 30852 39630 30986 39658
rect 12532 37868 12584 37874
rect 12532 37810 12584 37816
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 16396 37868 16448 37874
rect 16396 37810 16448 37816
rect 18604 37868 18656 37874
rect 18604 37810 18656 37816
rect 23848 37868 23900 37874
rect 23848 37810 23900 37816
rect 25228 37868 25280 37874
rect 25228 37810 25280 37816
rect 28080 37868 28132 37874
rect 28080 37810 28132 37816
rect 29736 37868 29788 37874
rect 29736 37810 29788 37816
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 848 37256 900 37262
rect 848 37198 900 37204
rect 860 36961 888 37198
rect 3332 37188 3384 37194
rect 3332 37130 3384 37136
rect 846 36952 902 36961
rect 846 36887 902 36896
rect 3344 30258 3372 37130
rect 12544 37126 12572 37810
rect 13084 37800 13136 37806
rect 13084 37742 13136 37748
rect 13728 37800 13780 37806
rect 13728 37742 13780 37748
rect 12992 37188 13044 37194
rect 12992 37130 13044 37136
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 12544 36922 12572 37062
rect 12532 36916 12584 36922
rect 12532 36858 12584 36864
rect 13004 36854 13032 37130
rect 12348 36848 12400 36854
rect 12348 36790 12400 36796
rect 12992 36848 13044 36854
rect 12992 36790 13044 36796
rect 11704 36576 11756 36582
rect 11704 36518 11756 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 11716 36242 11744 36518
rect 11704 36236 11756 36242
rect 11704 36178 11756 36184
rect 12360 36106 12388 36790
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 12452 36378 12480 36722
rect 13096 36582 13124 37742
rect 13452 37664 13504 37670
rect 13452 37606 13504 37612
rect 13464 37330 13492 37606
rect 13452 37324 13504 37330
rect 13452 37266 13504 37272
rect 13740 36718 13768 37742
rect 16040 37466 16068 37810
rect 16212 37664 16264 37670
rect 16212 37606 16264 37612
rect 15476 37460 15528 37466
rect 15476 37402 15528 37408
rect 16028 37460 16080 37466
rect 16028 37402 16080 37408
rect 14648 37256 14700 37262
rect 14648 37198 14700 37204
rect 14660 36786 14688 37198
rect 15200 37120 15252 37126
rect 15200 37062 15252 37068
rect 14648 36780 14700 36786
rect 14648 36722 14700 36728
rect 13728 36712 13780 36718
rect 13728 36654 13780 36660
rect 14372 36712 14424 36718
rect 14372 36654 14424 36660
rect 13084 36576 13136 36582
rect 13084 36518 13136 36524
rect 12440 36372 12492 36378
rect 12440 36314 12492 36320
rect 12992 36372 13044 36378
rect 12992 36314 13044 36320
rect 12348 36100 12400 36106
rect 12348 36042 12400 36048
rect 11520 36032 11572 36038
rect 11520 35974 11572 35980
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 11532 35154 11560 35974
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 11900 35290 11928 35634
rect 11888 35284 11940 35290
rect 11888 35226 11940 35232
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 11532 34066 11560 35090
rect 11900 34746 11928 35226
rect 12360 35018 12388 36042
rect 13004 35834 13032 36314
rect 13096 36174 13124 36518
rect 13740 36242 13768 36654
rect 14384 36378 14412 36654
rect 15212 36582 15240 37062
rect 15200 36576 15252 36582
rect 15200 36518 15252 36524
rect 14372 36372 14424 36378
rect 14372 36314 14424 36320
rect 13728 36236 13780 36242
rect 13728 36178 13780 36184
rect 13084 36168 13136 36174
rect 13084 36110 13136 36116
rect 12992 35828 13044 35834
rect 12992 35770 13044 35776
rect 13740 35630 13768 36178
rect 13728 35624 13780 35630
rect 13728 35566 13780 35572
rect 13360 35488 13412 35494
rect 13360 35430 13412 35436
rect 13372 35018 13400 35430
rect 15212 35154 15240 36518
rect 15488 36174 15516 37402
rect 16224 37330 16252 37606
rect 16212 37324 16264 37330
rect 16212 37266 16264 37272
rect 15568 37188 15620 37194
rect 15568 37130 15620 37136
rect 15580 36854 15608 37130
rect 16408 36922 16436 37810
rect 17500 37664 17552 37670
rect 17500 37606 17552 37612
rect 17512 37330 17540 37606
rect 18616 37466 18644 37810
rect 18696 37800 18748 37806
rect 18696 37742 18748 37748
rect 18880 37800 18932 37806
rect 18880 37742 18932 37748
rect 23664 37800 23716 37806
rect 23664 37742 23716 37748
rect 18604 37460 18656 37466
rect 18604 37402 18656 37408
rect 17500 37324 17552 37330
rect 17500 37266 17552 37272
rect 16488 37120 16540 37126
rect 16488 37062 16540 37068
rect 16396 36916 16448 36922
rect 16396 36858 16448 36864
rect 15568 36848 15620 36854
rect 15568 36790 15620 36796
rect 15476 36168 15528 36174
rect 15476 36110 15528 36116
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 14188 35148 14240 35154
rect 14188 35090 14240 35096
rect 15200 35148 15252 35154
rect 15200 35090 15252 35096
rect 12348 35012 12400 35018
rect 12348 34954 12400 34960
rect 13360 35012 13412 35018
rect 13360 34954 13412 34960
rect 11888 34740 11940 34746
rect 11888 34682 11940 34688
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 12084 34066 12112 34342
rect 11520 34060 11572 34066
rect 11520 34002 11572 34008
rect 12072 34060 12124 34066
rect 12072 34002 12124 34008
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 11532 33522 11560 34002
rect 12360 33862 12388 34954
rect 13544 34672 13596 34678
rect 13544 34614 13596 34620
rect 13084 34604 13136 34610
rect 13084 34546 13136 34552
rect 12716 34400 12768 34406
rect 12716 34342 12768 34348
rect 12348 33856 12400 33862
rect 12348 33798 12400 33804
rect 12360 33590 12388 33798
rect 12728 33658 12756 34342
rect 13096 33658 13124 34546
rect 13360 34536 13412 34542
rect 13360 34478 13412 34484
rect 12716 33652 12768 33658
rect 12716 33594 12768 33600
rect 13084 33652 13136 33658
rect 13084 33594 13136 33600
rect 12348 33584 12400 33590
rect 12348 33526 12400 33532
rect 11520 33516 11572 33522
rect 11520 33458 11572 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 13096 32978 13124 33594
rect 13372 32978 13400 34478
rect 13556 34202 13584 34614
rect 14200 34610 14228 35090
rect 15488 35018 15516 35430
rect 15580 35018 15608 36790
rect 16396 36780 16448 36786
rect 16396 36722 16448 36728
rect 16408 36242 16436 36722
rect 16500 36242 16528 37062
rect 18616 36922 18644 37402
rect 18708 37108 18736 37742
rect 18788 37120 18840 37126
rect 18708 37080 18788 37108
rect 18708 36922 18736 37080
rect 18788 37062 18840 37068
rect 18604 36916 18656 36922
rect 18604 36858 18656 36864
rect 18696 36916 18748 36922
rect 18696 36858 18748 36864
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 17132 36712 17184 36718
rect 17132 36654 17184 36660
rect 17684 36712 17736 36718
rect 17684 36654 17736 36660
rect 16396 36236 16448 36242
rect 16396 36178 16448 36184
rect 16488 36236 16540 36242
rect 16488 36178 16540 36184
rect 16408 35630 16436 36178
rect 17144 35894 17172 36654
rect 17500 36576 17552 36582
rect 17500 36518 17552 36524
rect 17512 36242 17540 36518
rect 17500 36236 17552 36242
rect 17500 36178 17552 36184
rect 16960 35866 17172 35894
rect 16960 35766 16988 35866
rect 16948 35760 17000 35766
rect 16948 35702 17000 35708
rect 16212 35624 16264 35630
rect 16212 35566 16264 35572
rect 16396 35624 16448 35630
rect 16396 35566 16448 35572
rect 15476 35012 15528 35018
rect 15476 34954 15528 34960
rect 15568 35012 15620 35018
rect 15568 34954 15620 34960
rect 15580 34610 15608 34954
rect 16224 34746 16252 35566
rect 16960 35290 16988 35702
rect 17592 35488 17644 35494
rect 17592 35430 17644 35436
rect 16948 35284 17000 35290
rect 16948 35226 17000 35232
rect 17604 35154 17632 35430
rect 17592 35148 17644 35154
rect 17592 35090 17644 35096
rect 16396 34944 16448 34950
rect 16396 34886 16448 34892
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 13820 34468 13872 34474
rect 13820 34410 13872 34416
rect 13544 34196 13596 34202
rect 13544 34138 13596 34144
rect 13084 32972 13136 32978
rect 13084 32914 13136 32920
rect 13360 32972 13412 32978
rect 13360 32914 13412 32920
rect 12072 32768 12124 32774
rect 12072 32710 12124 32716
rect 13084 32768 13136 32774
rect 13084 32710 13136 32716
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 11612 32360 11664 32366
rect 11612 32302 11664 32308
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 11624 31822 11652 32302
rect 12084 31890 12112 32710
rect 13096 32026 13124 32710
rect 13176 32360 13228 32366
rect 13176 32302 13228 32308
rect 13084 32020 13136 32026
rect 13084 31962 13136 31968
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 11612 31816 11664 31822
rect 11612 31758 11664 31764
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 9404 31408 9456 31414
rect 9324 31356 9404 31362
rect 9324 31350 9456 31356
rect 9324 31334 9444 31350
rect 8116 31272 8168 31278
rect 8116 31214 8168 31220
rect 8944 31272 8996 31278
rect 8944 31214 8996 31220
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 8128 30818 8156 31214
rect 8956 30938 8984 31214
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 8128 30802 8248 30818
rect 5632 30796 5684 30802
rect 8128 30796 8260 30802
rect 8128 30790 8208 30796
rect 5632 30738 5684 30744
rect 8208 30738 8260 30744
rect 8576 30796 8628 30802
rect 8576 30738 8628 30744
rect 3516 30728 3568 30734
rect 3516 30670 3568 30676
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 2596 30252 2648 30258
rect 2596 30194 2648 30200
rect 2964 30252 3016 30258
rect 2964 30194 3016 30200
rect 3332 30252 3384 30258
rect 3332 30194 3384 30200
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1122 29336 1178 29345
rect 1122 29271 1178 29280
rect 848 25424 900 25430
rect 846 25392 848 25401
rect 900 25392 902 25401
rect 846 25327 902 25336
rect 846 23760 902 23769
rect 846 23695 848 23704
rect 900 23695 902 23704
rect 848 23666 900 23672
rect 1136 22778 1164 29271
rect 1412 29102 1440 29582
rect 2608 29578 2636 30194
rect 2596 29572 2648 29578
rect 2596 29514 2648 29520
rect 2976 29238 3004 30194
rect 2964 29232 3016 29238
rect 2964 29174 3016 29180
rect 1400 29096 1452 29102
rect 1400 29038 1452 29044
rect 1676 29096 1728 29102
rect 1676 29038 1728 29044
rect 1412 27470 1440 29038
rect 1688 28762 1716 29038
rect 2872 29028 2924 29034
rect 2872 28970 2924 28976
rect 1676 28756 1728 28762
rect 1676 28698 1728 28704
rect 2884 28558 2912 28970
rect 2872 28552 2924 28558
rect 2872 28494 2924 28500
rect 2228 28416 2280 28422
rect 2228 28358 2280 28364
rect 2240 28082 2268 28358
rect 2884 28218 2912 28494
rect 2872 28212 2924 28218
rect 2872 28154 2924 28160
rect 2228 28076 2280 28082
rect 2228 28018 2280 28024
rect 2136 27872 2188 27878
rect 2136 27814 2188 27820
rect 2148 27674 2176 27814
rect 2136 27668 2188 27674
rect 2136 27610 2188 27616
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1860 27464 1912 27470
rect 1860 27406 1912 27412
rect 1676 26920 1728 26926
rect 1676 26862 1728 26868
rect 1688 26586 1716 26862
rect 1872 26790 1900 27406
rect 2872 27396 2924 27402
rect 2976 27384 3004 29174
rect 3528 28490 3556 30670
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 3792 30184 3844 30190
rect 4172 30138 4200 30534
rect 3792 30126 3844 30132
rect 3804 29850 3832 30126
rect 4080 30110 4200 30138
rect 3792 29844 3844 29850
rect 3792 29786 3844 29792
rect 4080 29730 4108 30110
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4528 29844 4580 29850
rect 4528 29786 4580 29792
rect 4080 29702 4200 29730
rect 4540 29714 4568 29786
rect 4172 29510 4200 29702
rect 4528 29708 4580 29714
rect 4528 29650 4580 29656
rect 4252 29640 4304 29646
rect 4252 29582 4304 29588
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 4160 29504 4212 29510
rect 4160 29446 4212 29452
rect 3620 28966 3648 29446
rect 4264 29306 4292 29582
rect 4540 29458 4568 29650
rect 4632 29646 4660 30670
rect 4712 30660 4764 30666
rect 4712 30602 4764 30608
rect 4724 30394 4752 30602
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4712 30388 4764 30394
rect 4712 30330 4764 30336
rect 5644 30258 5672 30738
rect 6368 30660 6420 30666
rect 6368 30602 6420 30608
rect 7472 30660 7524 30666
rect 7472 30602 7524 30608
rect 6380 30394 6408 30602
rect 6736 30592 6788 30598
rect 6736 30534 6788 30540
rect 6368 30388 6420 30394
rect 6368 30330 6420 30336
rect 5908 30320 5960 30326
rect 5908 30262 5960 30268
rect 5632 30252 5684 30258
rect 5632 30194 5684 30200
rect 5816 30252 5868 30258
rect 5816 30194 5868 30200
rect 5644 30161 5672 30194
rect 5724 30184 5776 30190
rect 5630 30152 5686 30161
rect 5724 30126 5776 30132
rect 5630 30087 5686 30096
rect 4712 30048 4764 30054
rect 4712 29990 4764 29996
rect 5172 30048 5224 30054
rect 5172 29990 5224 29996
rect 4724 29714 4752 29990
rect 5184 29850 5212 29990
rect 5172 29844 5224 29850
rect 5172 29786 5224 29792
rect 4712 29708 4764 29714
rect 4712 29650 4764 29656
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 4540 29430 4660 29458
rect 4252 29300 4304 29306
rect 4252 29242 4304 29248
rect 3976 29232 4028 29238
rect 3976 29174 4028 29180
rect 3608 28960 3660 28966
rect 3608 28902 3660 28908
rect 3620 28626 3648 28902
rect 3988 28626 4016 29174
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 3608 28620 3660 28626
rect 3608 28562 3660 28568
rect 3976 28620 4028 28626
rect 3976 28562 4028 28568
rect 3516 28484 3568 28490
rect 3516 28426 3568 28432
rect 3700 28484 3752 28490
rect 3700 28426 3752 28432
rect 3424 28144 3476 28150
rect 3424 28086 3476 28092
rect 3056 28008 3108 28014
rect 3436 27996 3464 28086
rect 3108 27968 3464 27996
rect 3056 27950 3108 27956
rect 3148 27872 3200 27878
rect 3148 27814 3200 27820
rect 3160 27538 3188 27814
rect 3436 27606 3464 27968
rect 3424 27600 3476 27606
rect 3424 27542 3476 27548
rect 3148 27532 3200 27538
rect 3148 27474 3200 27480
rect 2924 27356 3004 27384
rect 2872 27338 2924 27344
rect 2976 27062 3004 27356
rect 2964 27056 3016 27062
rect 2964 26998 3016 27004
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 1676 26580 1728 26586
rect 1676 26522 1728 26528
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 2228 26240 2280 26246
rect 2228 26182 2280 26188
rect 2240 25362 2268 26182
rect 2688 25968 2740 25974
rect 2688 25910 2740 25916
rect 2700 25430 2728 25910
rect 2792 25838 2820 26250
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2792 25498 2820 25774
rect 2780 25492 2832 25498
rect 2780 25434 2832 25440
rect 2688 25424 2740 25430
rect 2688 25366 2740 25372
rect 2228 25356 2280 25362
rect 2228 25298 2280 25304
rect 1584 25288 1636 25294
rect 1584 25230 1636 25236
rect 2136 25288 2188 25294
rect 2136 25230 2188 25236
rect 1596 24954 1624 25230
rect 1860 25152 1912 25158
rect 1860 25094 1912 25100
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1872 24138 1900 25094
rect 2148 24954 2176 25230
rect 2700 24954 2728 25366
rect 2792 25362 2820 25434
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2136 24948 2188 24954
rect 2136 24890 2188 24896
rect 2688 24948 2740 24954
rect 2688 24890 2740 24896
rect 1860 24132 1912 24138
rect 1860 24074 1912 24080
rect 2148 23730 2176 24890
rect 2976 24886 3004 26998
rect 3160 26790 3188 27474
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 3160 26450 3188 26726
rect 3148 26444 3200 26450
rect 3148 26386 3200 26392
rect 3528 25498 3556 28426
rect 3712 28150 3740 28426
rect 3700 28144 3752 28150
rect 3700 28086 3752 28092
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3620 27674 3648 28018
rect 3608 27668 3660 27674
rect 3608 27610 3660 27616
rect 3620 27470 3648 27610
rect 3608 27464 3660 27470
rect 3608 27406 3660 27412
rect 3712 26042 3740 28086
rect 3988 28082 4016 28562
rect 4080 28082 4108 28698
rect 4632 28642 4660 29430
rect 4540 28614 4660 28642
rect 4540 28422 4568 28614
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 4528 28416 4580 28422
rect 4528 28358 4580 28364
rect 4540 28082 4568 28358
rect 3976 28076 4028 28082
rect 3976 28018 4028 28024
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 4528 28076 4580 28082
rect 4528 28018 4580 28024
rect 4632 27878 4660 28494
rect 4620 27872 4672 27878
rect 4620 27814 4672 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27674 4660 27814
rect 4620 27668 4672 27674
rect 4620 27610 4672 27616
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 3700 26036 3752 26042
rect 3700 25978 3752 25984
rect 3792 25900 3844 25906
rect 3792 25842 3844 25848
rect 3516 25492 3568 25498
rect 3516 25434 3568 25440
rect 3804 25362 3832 25842
rect 4080 25838 4108 27542
rect 4724 26926 4752 29650
rect 4896 29640 4948 29646
rect 4816 29588 4896 29594
rect 4816 29582 4948 29588
rect 4816 29566 4936 29582
rect 5540 29572 5592 29578
rect 4816 28694 4844 29566
rect 5540 29514 5592 29520
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5552 29306 5580 29514
rect 5540 29300 5592 29306
rect 5540 29242 5592 29248
rect 5356 29232 5408 29238
rect 5356 29174 5408 29180
rect 4804 28688 4856 28694
rect 4804 28630 4856 28636
rect 5368 28422 5396 29174
rect 5736 29170 5764 30126
rect 5828 29238 5856 30194
rect 5920 29578 5948 30262
rect 6748 30122 6776 30534
rect 7484 30326 7512 30602
rect 7472 30320 7524 30326
rect 7472 30262 7524 30268
rect 7840 30252 7892 30258
rect 7840 30194 7892 30200
rect 8116 30252 8168 30258
rect 8116 30194 8168 30200
rect 6736 30116 6788 30122
rect 6736 30058 6788 30064
rect 5908 29572 5960 29578
rect 5908 29514 5960 29520
rect 5920 29306 5948 29514
rect 6092 29504 6144 29510
rect 6092 29446 6144 29452
rect 5908 29300 5960 29306
rect 5908 29242 5960 29248
rect 5816 29232 5868 29238
rect 5816 29174 5868 29180
rect 6104 29170 6132 29446
rect 6460 29300 6512 29306
rect 6460 29242 6512 29248
rect 5724 29164 5776 29170
rect 5724 29106 5776 29112
rect 6092 29164 6144 29170
rect 6092 29106 6144 29112
rect 5908 28960 5960 28966
rect 5908 28902 5960 28908
rect 5724 28484 5776 28490
rect 5724 28426 5776 28432
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5368 28150 5396 28358
rect 5736 28150 5764 28426
rect 5816 28416 5868 28422
rect 5816 28358 5868 28364
rect 5264 28144 5316 28150
rect 5264 28086 5316 28092
rect 5356 28144 5408 28150
rect 5356 28086 5408 28092
rect 5724 28144 5776 28150
rect 5724 28086 5776 28092
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5276 26994 5304 28086
rect 5368 27334 5396 28086
rect 5632 27940 5684 27946
rect 5632 27882 5684 27888
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 5460 27470 5488 27814
rect 5644 27554 5672 27882
rect 5736 27674 5764 28086
rect 5724 27668 5776 27674
rect 5724 27610 5776 27616
rect 5644 27526 5764 27554
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 5264 26988 5316 26994
rect 5264 26930 5316 26936
rect 4712 26920 4764 26926
rect 4712 26862 4764 26868
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26586 4660 26726
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4724 26466 4752 26862
rect 4540 26450 4752 26466
rect 4528 26444 4752 26450
rect 4580 26438 4752 26444
rect 4528 26386 4580 26392
rect 4620 26240 4672 26246
rect 4620 26182 4672 26188
rect 4068 25832 4120 25838
rect 4068 25774 4120 25780
rect 3148 25356 3200 25362
rect 3148 25298 3200 25304
rect 3792 25356 3844 25362
rect 3792 25298 3844 25304
rect 2964 24880 3016 24886
rect 2964 24822 3016 24828
rect 2976 24562 3004 24822
rect 3160 24818 3188 25298
rect 3332 25152 3384 25158
rect 3332 25094 3384 25100
rect 3148 24812 3200 24818
rect 3148 24754 3200 24760
rect 3056 24608 3108 24614
rect 2976 24556 3056 24562
rect 2976 24550 3108 24556
rect 2976 24534 3096 24550
rect 2976 24206 3004 24534
rect 3160 24274 3188 24754
rect 3344 24750 3372 25094
rect 4080 24834 4108 25774
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25412 4660 26182
rect 4724 26042 4752 26438
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4540 25384 4660 25412
rect 4540 25226 4568 25384
rect 4344 25220 4396 25226
rect 4344 25162 4396 25168
rect 4528 25220 4580 25226
rect 4528 25162 4580 25168
rect 4356 24954 4384 25162
rect 4344 24948 4396 24954
rect 4344 24890 4396 24896
rect 4540 24886 4568 25162
rect 4528 24880 4580 24886
rect 4080 24818 4200 24834
rect 4528 24822 4580 24828
rect 4816 24818 4844 26930
rect 5368 26790 5396 27270
rect 5460 27062 5488 27406
rect 5552 27130 5580 27406
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 5356 26784 5408 26790
rect 5632 26784 5684 26790
rect 5356 26726 5408 26732
rect 5630 26752 5632 26761
rect 5684 26752 5686 26761
rect 5630 26687 5686 26696
rect 5736 26382 5764 27526
rect 5828 27470 5856 28358
rect 5920 28218 5948 28902
rect 6000 28756 6052 28762
rect 6000 28698 6052 28704
rect 5908 28212 5960 28218
rect 5908 28154 5960 28160
rect 6012 28098 6040 28698
rect 6104 28490 6132 29106
rect 6092 28484 6144 28490
rect 6092 28426 6144 28432
rect 6104 28218 6132 28426
rect 6092 28212 6144 28218
rect 6092 28154 6144 28160
rect 5920 28070 6040 28098
rect 5920 28014 5948 28070
rect 5908 28008 5960 28014
rect 5908 27950 5960 27956
rect 6000 27940 6052 27946
rect 6000 27882 6052 27888
rect 5816 27464 5868 27470
rect 5816 27406 5868 27412
rect 5816 27056 5868 27062
rect 5816 26998 5868 27004
rect 5828 26518 5856 26998
rect 5908 26920 5960 26926
rect 5908 26862 5960 26868
rect 5920 26586 5948 26862
rect 6012 26790 6040 27882
rect 6104 27878 6132 28154
rect 6092 27872 6144 27878
rect 6092 27814 6144 27820
rect 6276 27872 6328 27878
rect 6276 27814 6328 27820
rect 6092 27532 6144 27538
rect 6092 27474 6144 27480
rect 6104 26790 6132 27474
rect 6184 27328 6236 27334
rect 6184 27270 6236 27276
rect 6196 27130 6224 27270
rect 6184 27124 6236 27130
rect 6184 27066 6236 27072
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 6092 26784 6144 26790
rect 6092 26726 6144 26732
rect 5908 26580 5960 26586
rect 5908 26522 5960 26528
rect 5816 26512 5868 26518
rect 5816 26454 5868 26460
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5828 25922 5856 26454
rect 5644 25894 5856 25922
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5368 24818 5396 25434
rect 5448 25220 5500 25226
rect 5448 25162 5500 25168
rect 5460 24886 5488 25162
rect 5448 24880 5500 24886
rect 5448 24822 5500 24828
rect 4080 24812 4212 24818
rect 4080 24806 4160 24812
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 1124 22772 1176 22778
rect 1124 22714 1176 22720
rect 2700 22710 2728 22918
rect 2688 22704 2740 22710
rect 2688 22646 2740 22652
rect 2792 22574 2820 23054
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 1676 22432 1728 22438
rect 1676 22374 1728 22380
rect 1688 22234 1716 22374
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 2792 22166 2820 22510
rect 2780 22160 2832 22166
rect 2780 22102 2832 22108
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21486 1440 21966
rect 2976 21962 3004 24142
rect 3160 23186 3188 24210
rect 3712 23798 3740 24550
rect 4080 24274 4108 24806
rect 4160 24754 4212 24760
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24268 4120 24274
rect 4068 24210 4120 24216
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5368 23798 5396 24754
rect 5644 23866 5672 25894
rect 5724 25832 5776 25838
rect 5724 25774 5776 25780
rect 5736 25294 5764 25774
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5736 24954 5764 25230
rect 5724 24948 5776 24954
rect 5724 24890 5776 24896
rect 5736 24682 5764 24890
rect 5724 24676 5776 24682
rect 5724 24618 5776 24624
rect 5632 23860 5684 23866
rect 5632 23802 5684 23808
rect 3700 23792 3752 23798
rect 3700 23734 3752 23740
rect 5080 23792 5132 23798
rect 5080 23734 5132 23740
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 3148 23180 3200 23186
rect 3148 23122 3200 23128
rect 3160 22642 3188 23122
rect 3712 23118 3740 23734
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5092 23322 5120 23734
rect 5828 23594 5856 25638
rect 5920 25498 5948 26522
rect 6288 26450 6316 27814
rect 6472 27402 6500 29242
rect 6748 28762 6776 30058
rect 7852 29850 7880 30194
rect 8128 29850 8156 30194
rect 8220 29850 8248 30738
rect 8300 30592 8352 30598
rect 8300 30534 8352 30540
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 8312 30122 8340 30534
rect 8300 30116 8352 30122
rect 8300 30058 8352 30064
rect 8496 30054 8524 30534
rect 8588 30394 8616 30738
rect 8576 30388 8628 30394
rect 8576 30330 8628 30336
rect 8760 30320 8812 30326
rect 8760 30262 8812 30268
rect 8484 30048 8536 30054
rect 8484 29990 8536 29996
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 8116 29844 8168 29850
rect 8116 29786 8168 29792
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7760 28762 7788 29038
rect 6736 28756 6788 28762
rect 6736 28698 6788 28704
rect 7748 28756 7800 28762
rect 7748 28698 7800 28704
rect 8128 28558 8156 29786
rect 8220 28966 8248 29786
rect 8496 29782 8524 29990
rect 8484 29776 8536 29782
rect 8484 29718 8536 29724
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 8220 28014 8248 28902
rect 8312 28762 8340 29582
rect 8496 29510 8524 29582
rect 8772 29578 8800 30262
rect 9128 30184 9180 30190
rect 9126 30152 9128 30161
rect 9180 30152 9182 30161
rect 9126 30087 9182 30096
rect 9220 30116 9272 30122
rect 9220 30058 9272 30064
rect 9232 29646 9260 30058
rect 9220 29640 9272 29646
rect 9220 29582 9272 29588
rect 8760 29572 8812 29578
rect 8760 29514 8812 29520
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8300 28756 8352 28762
rect 8300 28698 8352 28704
rect 8772 28558 8800 29514
rect 9128 29504 9180 29510
rect 9128 29446 9180 29452
rect 8760 28552 8812 28558
rect 8760 28494 8812 28500
rect 6828 28008 6880 28014
rect 6828 27950 6880 27956
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 6840 27674 6868 27950
rect 6828 27668 6880 27674
rect 6828 27610 6880 27616
rect 6552 27600 6604 27606
rect 6552 27542 6604 27548
rect 6460 27396 6512 27402
rect 6460 27338 6512 27344
rect 6460 26852 6512 26858
rect 6460 26794 6512 26800
rect 6368 26580 6420 26586
rect 6368 26522 6420 26528
rect 6276 26444 6328 26450
rect 6276 26386 6328 26392
rect 6000 26308 6052 26314
rect 6000 26250 6052 26256
rect 5908 25492 5960 25498
rect 5908 25434 5960 25440
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5920 24818 5948 25230
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5816 23588 5868 23594
rect 5816 23530 5868 23536
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5080 23316 5132 23322
rect 5080 23258 5132 23264
rect 5276 23186 5304 23462
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 3700 23112 3752 23118
rect 3976 23112 4028 23118
rect 3752 23060 3832 23066
rect 3700 23054 3832 23060
rect 3976 23054 4028 23060
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 3712 23038 3832 23054
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3436 22710 3464 22918
rect 3424 22704 3476 22710
rect 3424 22646 3476 22652
rect 3700 22704 3752 22710
rect 3700 22646 3752 22652
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2976 21622 3004 21898
rect 3712 21622 3740 22646
rect 3804 22094 3832 23038
rect 3988 22234 4016 23054
rect 4080 22574 4108 23054
rect 5552 23050 5580 23462
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 5540 23044 5592 23050
rect 5540 22986 5592 22992
rect 4816 22710 4844 22986
rect 5264 22976 5316 22982
rect 5264 22918 5316 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4804 22704 4856 22710
rect 4632 22664 4804 22692
rect 4068 22568 4120 22574
rect 4068 22510 4120 22516
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 4080 22094 4108 22510
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3804 22066 3924 22094
rect 4080 22066 4200 22094
rect 3896 21962 3924 22066
rect 3976 22024 4028 22030
rect 4172 22012 4200 22066
rect 4028 21984 4200 22012
rect 3976 21966 4028 21972
rect 3884 21956 3936 21962
rect 3884 21898 3936 21904
rect 4344 21956 4396 21962
rect 4344 21898 4396 21904
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4356 21842 4384 21898
rect 4632 21842 4660 22664
rect 4804 22646 4856 22652
rect 5276 22574 5304 22918
rect 5540 22704 5592 22710
rect 5460 22664 5540 22692
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 2964 21616 3016 21622
rect 2964 21558 3016 21564
rect 3700 21616 3752 21622
rect 3700 21558 3752 21564
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 21010 1440 21422
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 19310 1440 20946
rect 2976 20874 3004 21558
rect 3424 21480 3476 21486
rect 4172 21434 4200 21830
rect 4356 21814 4660 21842
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 3424 21422 3476 21428
rect 3436 21146 3464 21422
rect 4080 21406 4200 21434
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3896 20942 3924 21286
rect 4080 20942 4108 21406
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21010 4660 21814
rect 4724 21350 4752 21830
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4816 20874 4844 22510
rect 5460 22438 5488 22664
rect 5540 22646 5592 22652
rect 5632 22704 5684 22710
rect 5632 22646 5684 22652
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 5448 22432 5500 22438
rect 5448 22374 5500 22380
rect 4908 22098 4936 22374
rect 5460 22234 5488 22374
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 4896 22092 4948 22098
rect 5644 22094 5672 22646
rect 5724 22500 5776 22506
rect 5724 22442 5776 22448
rect 4896 22034 4948 22040
rect 5552 22066 5672 22094
rect 5736 22094 5764 22442
rect 5816 22094 5868 22098
rect 5736 22092 5868 22094
rect 5736 22066 5816 22092
rect 5552 21894 5580 22066
rect 5816 22034 5868 22040
rect 6012 21894 6040 26250
rect 6380 25498 6408 26522
rect 6472 25906 6500 26794
rect 6564 26450 6592 27542
rect 8220 27538 8248 27950
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 6736 27056 6788 27062
rect 6736 26998 6788 27004
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6460 25900 6512 25906
rect 6460 25842 6512 25848
rect 6460 25764 6512 25770
rect 6460 25706 6512 25712
rect 6368 25492 6420 25498
rect 6368 25434 6420 25440
rect 6472 25378 6500 25706
rect 6092 25356 6144 25362
rect 6092 25298 6144 25304
rect 6380 25350 6500 25378
rect 6104 24954 6132 25298
rect 6380 25294 6408 25350
rect 6564 25294 6592 26386
rect 6748 25922 6776 26998
rect 6840 26926 6868 26998
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6656 25894 6776 25922
rect 6656 25378 6684 25894
rect 6736 25832 6788 25838
rect 6736 25774 6788 25780
rect 6748 25498 6776 25774
rect 6736 25492 6788 25498
rect 6736 25434 6788 25440
rect 6840 25430 6868 26182
rect 6828 25424 6880 25430
rect 6656 25350 6776 25378
rect 6828 25366 6880 25372
rect 6748 25294 6776 25350
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 6552 25288 6604 25294
rect 6552 25230 6604 25236
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6092 24948 6144 24954
rect 6092 24890 6144 24896
rect 6380 24886 6408 25230
rect 6368 24880 6420 24886
rect 6368 24822 6420 24828
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 6196 21894 6224 23462
rect 6380 23322 6408 24822
rect 6748 24818 6776 25230
rect 6932 25226 6960 27270
rect 8128 26858 8156 27270
rect 7380 26852 7432 26858
rect 7380 26794 7432 26800
rect 8116 26852 8168 26858
rect 8116 26794 8168 26800
rect 7104 26784 7156 26790
rect 7102 26752 7104 26761
rect 7156 26752 7158 26761
rect 7102 26687 7158 26696
rect 7392 26450 7420 26794
rect 8220 26586 8248 27474
rect 8772 27062 8800 28494
rect 9140 28014 9168 29446
rect 9232 29034 9260 29582
rect 9324 29510 9352 31334
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9956 31136 10008 31142
rect 9956 31078 10008 31084
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9404 30252 9456 30258
rect 9404 30194 9456 30200
rect 9416 29578 9444 30194
rect 9496 30048 9548 30054
rect 9600 30002 9628 30330
rect 9692 30326 9720 31078
rect 9968 30734 9996 31078
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 9680 30320 9732 30326
rect 9680 30262 9732 30268
rect 9548 29996 9628 30002
rect 9496 29990 9628 29996
rect 9508 29974 9628 29990
rect 9404 29572 9456 29578
rect 9404 29514 9456 29520
rect 9312 29504 9364 29510
rect 9312 29446 9364 29452
rect 9324 29306 9352 29446
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9220 29028 9272 29034
rect 9220 28970 9272 28976
rect 9600 28966 9628 29974
rect 9692 29102 9720 30262
rect 9784 30190 9812 30670
rect 11624 30258 11652 31758
rect 13188 31482 13216 32302
rect 13176 31476 13228 31482
rect 13176 31418 13228 31424
rect 13372 30938 13400 32914
rect 13544 32020 13596 32026
rect 13544 31962 13596 31968
rect 13556 31482 13584 31962
rect 13832 31958 13860 34410
rect 14200 34066 14228 34546
rect 14280 34196 14332 34202
rect 14280 34138 14332 34144
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 14292 33590 14320 34138
rect 15568 34060 15620 34066
rect 15568 34002 15620 34008
rect 15580 33930 15608 34002
rect 16408 33930 16436 34886
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 15568 33924 15620 33930
rect 15568 33866 15620 33872
rect 15936 33924 15988 33930
rect 15936 33866 15988 33872
rect 16396 33924 16448 33930
rect 16396 33866 16448 33872
rect 14280 33584 14332 33590
rect 14280 33526 14332 33532
rect 15396 33522 15424 33866
rect 15384 33516 15436 33522
rect 15384 33458 15436 33464
rect 13912 33448 13964 33454
rect 13912 33390 13964 33396
rect 13924 32910 13952 33390
rect 13912 32904 13964 32910
rect 13912 32846 13964 32852
rect 13924 32230 13952 32846
rect 15580 32502 15608 33866
rect 15948 33658 15976 33866
rect 15936 33652 15988 33658
rect 15936 33594 15988 33600
rect 16408 33522 16436 33866
rect 17408 33856 17460 33862
rect 17408 33798 17460 33804
rect 17420 33658 17448 33798
rect 17696 33658 17724 36654
rect 18800 36378 18828 36722
rect 18512 36372 18564 36378
rect 18512 36314 18564 36320
rect 18788 36372 18840 36378
rect 18788 36314 18840 36320
rect 18144 36032 18196 36038
rect 18144 35974 18196 35980
rect 18156 35154 18184 35974
rect 18524 35834 18552 36314
rect 18512 35828 18564 35834
rect 18512 35770 18564 35776
rect 18892 35630 18920 37742
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 22388 37330 22416 37606
rect 23676 37466 23704 37742
rect 23664 37460 23716 37466
rect 23664 37402 23716 37408
rect 23860 37398 23888 37810
rect 24860 37800 24912 37806
rect 24860 37742 24912 37748
rect 27252 37800 27304 37806
rect 27252 37742 27304 37748
rect 24400 37460 24452 37466
rect 24400 37402 24452 37408
rect 23848 37392 23900 37398
rect 23848 37334 23900 37340
rect 21548 37324 21600 37330
rect 21548 37266 21600 37272
rect 22376 37324 22428 37330
rect 22376 37266 22428 37272
rect 19432 37188 19484 37194
rect 21272 37188 21324 37194
rect 19484 37148 19564 37176
rect 19432 37130 19484 37136
rect 19536 36854 19564 37148
rect 21272 37130 21324 37136
rect 21456 37188 21508 37194
rect 21456 37130 21508 37136
rect 19892 37120 19944 37126
rect 19892 37062 19944 37068
rect 20076 37120 20128 37126
rect 20076 37062 20128 37068
rect 20536 37120 20588 37126
rect 20536 37062 20588 37068
rect 19524 36848 19576 36854
rect 19524 36790 19576 36796
rect 19536 36106 19564 36790
rect 19904 36718 19932 37062
rect 19892 36712 19944 36718
rect 19892 36654 19944 36660
rect 20088 36582 20116 37062
rect 20548 36718 20576 37062
rect 21284 36786 21312 37130
rect 21272 36780 21324 36786
rect 21272 36722 21324 36728
rect 20536 36712 20588 36718
rect 20536 36654 20588 36660
rect 20812 36712 20864 36718
rect 20812 36654 20864 36660
rect 20996 36712 21048 36718
rect 20996 36654 21048 36660
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19524 36100 19576 36106
rect 19524 36042 19576 36048
rect 19064 35692 19116 35698
rect 19064 35634 19116 35640
rect 18880 35624 18932 35630
rect 18880 35566 18932 35572
rect 19076 35290 19104 35634
rect 19064 35284 19116 35290
rect 19064 35226 19116 35232
rect 18144 35148 18196 35154
rect 18144 35090 18196 35096
rect 19800 35148 19852 35154
rect 19800 35090 19852 35096
rect 18880 35080 18932 35086
rect 18880 35022 18932 35028
rect 18892 34746 18920 35022
rect 19524 35012 19576 35018
rect 19524 34954 19576 34960
rect 19156 34944 19208 34950
rect 19156 34886 19208 34892
rect 18880 34740 18932 34746
rect 18880 34682 18932 34688
rect 17776 34536 17828 34542
rect 17776 34478 17828 34484
rect 17788 33930 17816 34478
rect 18892 33998 18920 34682
rect 19168 34542 19196 34886
rect 19536 34678 19564 34954
rect 19812 34746 19840 35090
rect 19800 34740 19852 34746
rect 19800 34682 19852 34688
rect 19340 34672 19392 34678
rect 19340 34614 19392 34620
rect 19524 34672 19576 34678
rect 19524 34614 19576 34620
rect 19156 34536 19208 34542
rect 19156 34478 19208 34484
rect 19352 34066 19380 34614
rect 19616 34400 19668 34406
rect 19616 34342 19668 34348
rect 19340 34060 19392 34066
rect 19340 34002 19392 34008
rect 18880 33992 18932 33998
rect 18880 33934 18932 33940
rect 17776 33924 17828 33930
rect 17776 33866 17828 33872
rect 19524 33924 19576 33930
rect 19524 33866 19576 33872
rect 17408 33652 17460 33658
rect 17408 33594 17460 33600
rect 17684 33652 17736 33658
rect 17684 33594 17736 33600
rect 16396 33516 16448 33522
rect 16396 33458 16448 33464
rect 17040 33516 17092 33522
rect 17040 33458 17092 33464
rect 16408 32842 16436 33458
rect 17052 33114 17080 33458
rect 17696 33454 17724 33594
rect 17788 33590 17816 33866
rect 19536 33590 19564 33866
rect 19628 33658 19656 34342
rect 19708 33924 19760 33930
rect 19708 33866 19760 33872
rect 19720 33658 19748 33866
rect 19616 33652 19668 33658
rect 19616 33594 19668 33600
rect 19708 33652 19760 33658
rect 19708 33594 19760 33600
rect 17776 33584 17828 33590
rect 17776 33526 17828 33532
rect 19524 33584 19576 33590
rect 19524 33526 19576 33532
rect 17684 33448 17736 33454
rect 17684 33390 17736 33396
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 17040 33108 17092 33114
rect 17040 33050 17092 33056
rect 18064 32858 18092 33390
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 18524 32978 18552 33254
rect 19628 33046 19656 33594
rect 19708 33516 19760 33522
rect 19708 33458 19760 33464
rect 19616 33040 19668 33046
rect 19616 32982 19668 32988
rect 19720 32978 19748 33458
rect 19812 33386 19840 34682
rect 19996 34066 20024 36110
rect 20548 36106 20576 36654
rect 20536 36100 20588 36106
rect 20536 36042 20588 36048
rect 20824 35766 20852 36654
rect 21008 36378 21036 36654
rect 20996 36372 21048 36378
rect 20996 36314 21048 36320
rect 20904 36236 20956 36242
rect 20904 36178 20956 36184
rect 20916 35834 20944 36178
rect 21008 35834 21036 36314
rect 21284 36106 21312 36722
rect 21468 36650 21496 37130
rect 21456 36644 21508 36650
rect 21456 36586 21508 36592
rect 21364 36576 21416 36582
rect 21364 36518 21416 36524
rect 21272 36100 21324 36106
rect 21272 36042 21324 36048
rect 20904 35828 20956 35834
rect 20904 35770 20956 35776
rect 20996 35828 21048 35834
rect 20996 35770 21048 35776
rect 20812 35760 20864 35766
rect 20812 35702 20864 35708
rect 20260 35624 20312 35630
rect 20260 35566 20312 35572
rect 19984 34060 20036 34066
rect 19984 34002 20036 34008
rect 20272 33454 20300 35566
rect 20536 34944 20588 34950
rect 20536 34886 20588 34892
rect 20548 34746 20576 34886
rect 20536 34740 20588 34746
rect 20456 34700 20536 34728
rect 20456 33658 20484 34700
rect 20536 34682 20588 34688
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20640 34066 20668 34546
rect 20628 34060 20680 34066
rect 20628 34002 20680 34008
rect 21284 33930 21312 36042
rect 21376 35834 21404 36518
rect 21560 35894 21588 37266
rect 22284 37188 22336 37194
rect 22284 37130 22336 37136
rect 22008 37120 22060 37126
rect 22008 37062 22060 37068
rect 22020 36922 22048 37062
rect 22008 36916 22060 36922
rect 22008 36858 22060 36864
rect 21824 36848 21876 36854
rect 21824 36790 21876 36796
rect 21836 36378 21864 36790
rect 22296 36786 22324 37130
rect 23860 36922 23888 37334
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 24412 36854 24440 37402
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 21824 36372 21876 36378
rect 21824 36314 21876 36320
rect 21468 35866 21588 35894
rect 21364 35828 21416 35834
rect 21364 35770 21416 35776
rect 21468 35630 21496 35866
rect 22296 35766 22324 36722
rect 24124 36712 24176 36718
rect 24124 36654 24176 36660
rect 24136 35834 24164 36654
rect 24872 36650 24900 37742
rect 25412 37664 25464 37670
rect 25412 37606 25464 37612
rect 25424 36922 25452 37606
rect 26148 37256 26200 37262
rect 26148 37198 26200 37204
rect 25872 37188 25924 37194
rect 25872 37130 25924 37136
rect 25884 36922 25912 37130
rect 25412 36916 25464 36922
rect 25412 36858 25464 36864
rect 25872 36916 25924 36922
rect 25872 36858 25924 36864
rect 25964 36780 26016 36786
rect 25964 36722 26016 36728
rect 25504 36712 25556 36718
rect 25502 36680 25504 36689
rect 25556 36680 25558 36689
rect 24676 36644 24728 36650
rect 24676 36586 24728 36592
rect 24860 36644 24912 36650
rect 25502 36615 25558 36624
rect 24860 36586 24912 36592
rect 24688 36038 24716 36586
rect 24768 36100 24820 36106
rect 24768 36042 24820 36048
rect 24676 36032 24728 36038
rect 24676 35974 24728 35980
rect 24124 35828 24176 35834
rect 24124 35770 24176 35776
rect 22284 35760 22336 35766
rect 22284 35702 22336 35708
rect 23570 35728 23626 35737
rect 23570 35663 23572 35672
rect 23624 35663 23626 35672
rect 23572 35634 23624 35640
rect 21456 35624 21508 35630
rect 21456 35566 21508 35572
rect 21468 34406 21496 35566
rect 24400 35080 24452 35086
rect 24400 35022 24452 35028
rect 23480 34604 23532 34610
rect 23480 34546 23532 34552
rect 22560 34536 22612 34542
rect 22560 34478 22612 34484
rect 21456 34400 21508 34406
rect 21456 34342 21508 34348
rect 22100 34400 22152 34406
rect 22100 34342 22152 34348
rect 21272 33924 21324 33930
rect 21272 33866 21324 33872
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20444 33652 20496 33658
rect 20444 33594 20496 33600
rect 20352 33584 20404 33590
rect 20352 33526 20404 33532
rect 20260 33448 20312 33454
rect 20260 33390 20312 33396
rect 19800 33380 19852 33386
rect 19800 33322 19852 33328
rect 18512 32972 18564 32978
rect 18512 32914 18564 32920
rect 19708 32972 19760 32978
rect 19708 32914 19760 32920
rect 19064 32904 19116 32910
rect 18064 32842 18276 32858
rect 19064 32846 19116 32852
rect 16396 32836 16448 32842
rect 16396 32778 16448 32784
rect 18064 32836 18288 32842
rect 18064 32830 18236 32836
rect 16408 32502 16436 32778
rect 18064 32570 18092 32830
rect 18236 32778 18288 32784
rect 18052 32564 18104 32570
rect 18052 32506 18104 32512
rect 15568 32496 15620 32502
rect 15568 32438 15620 32444
rect 16396 32496 16448 32502
rect 16396 32438 16448 32444
rect 14280 32428 14332 32434
rect 14280 32370 14332 32376
rect 13912 32224 13964 32230
rect 13912 32166 13964 32172
rect 14188 32224 14240 32230
rect 14188 32166 14240 32172
rect 13820 31952 13872 31958
rect 13820 31894 13872 31900
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13832 31278 13860 31894
rect 14200 31822 14228 32166
rect 14292 31890 14320 32370
rect 15292 32360 15344 32366
rect 15292 32302 15344 32308
rect 15936 32360 15988 32366
rect 15936 32302 15988 32308
rect 14832 32224 14884 32230
rect 14832 32166 14884 32172
rect 14844 31890 14872 32166
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14832 31884 14884 31890
rect 14832 31826 14884 31832
rect 14188 31816 14240 31822
rect 14188 31758 14240 31764
rect 14200 31346 14228 31758
rect 14464 31680 14516 31686
rect 14464 31622 14516 31628
rect 14476 31414 14504 31622
rect 14844 31482 14872 31826
rect 15304 31822 15332 32302
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 15580 31890 15608 32166
rect 15568 31884 15620 31890
rect 15568 31826 15620 31832
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 14832 31476 14884 31482
rect 14832 31418 14884 31424
rect 14464 31408 14516 31414
rect 14464 31350 14516 31356
rect 14188 31340 14240 31346
rect 14188 31282 14240 31288
rect 13820 31272 13872 31278
rect 13820 31214 13872 31220
rect 13360 30932 13412 30938
rect 13360 30874 13412 30880
rect 12624 30592 12676 30598
rect 12624 30534 12676 30540
rect 13176 30592 13228 30598
rect 13176 30534 13228 30540
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 10784 30252 10836 30258
rect 10784 30194 10836 30200
rect 11612 30252 11664 30258
rect 11612 30194 11664 30200
rect 9772 30184 9824 30190
rect 9772 30126 9824 30132
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 9784 29102 9812 30126
rect 9956 30048 10008 30054
rect 9956 29990 10008 29996
rect 9968 29714 9996 29990
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 10416 29708 10468 29714
rect 10416 29650 10468 29656
rect 10428 29578 10456 29650
rect 10416 29572 10468 29578
rect 10416 29514 10468 29520
rect 10520 29306 10548 30126
rect 10600 29504 10652 29510
rect 10600 29446 10652 29452
rect 10508 29300 10560 29306
rect 10508 29242 10560 29248
rect 10612 29170 10640 29446
rect 10796 29238 10824 30194
rect 12636 30190 12664 30534
rect 12624 30184 12676 30190
rect 12624 30126 12676 30132
rect 13188 30054 13216 30534
rect 13268 30320 13320 30326
rect 13268 30262 13320 30268
rect 12992 30048 13044 30054
rect 12992 29990 13044 29996
rect 13176 30048 13228 30054
rect 13176 29990 13228 29996
rect 11520 29640 11572 29646
rect 11520 29582 11572 29588
rect 10784 29232 10836 29238
rect 10784 29174 10836 29180
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9036 28008 9088 28014
rect 9036 27950 9088 27956
rect 9128 28008 9180 28014
rect 9128 27950 9180 27956
rect 9048 27674 9076 27950
rect 9036 27668 9088 27674
rect 9036 27610 9088 27616
rect 9140 27470 9168 27950
rect 10048 27940 10100 27946
rect 10048 27882 10100 27888
rect 10060 27470 10088 27882
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 10048 27464 10100 27470
rect 10048 27406 10100 27412
rect 10140 27464 10192 27470
rect 10140 27406 10192 27412
rect 8760 27056 8812 27062
rect 8760 26998 8812 27004
rect 8392 26988 8444 26994
rect 8392 26930 8444 26936
rect 8208 26580 8260 26586
rect 8208 26522 8260 26528
rect 7380 26444 7432 26450
rect 7380 26386 7432 26392
rect 7656 26308 7708 26314
rect 7656 26250 7708 26256
rect 7668 25974 7696 26250
rect 8220 25974 8248 26522
rect 7656 25968 7708 25974
rect 7656 25910 7708 25916
rect 8208 25968 8260 25974
rect 8208 25910 8260 25916
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 6920 25220 6972 25226
rect 6920 25162 6972 25168
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6748 24614 6776 24754
rect 6552 24608 6604 24614
rect 6552 24550 6604 24556
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 6564 23730 6592 24550
rect 6748 24138 6776 24550
rect 6932 24206 6960 25162
rect 7024 24886 7052 25842
rect 7012 24880 7064 24886
rect 7012 24822 7064 24828
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 7116 24410 7144 24686
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6932 23730 6960 24142
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6368 23316 6420 23322
rect 6368 23258 6420 23264
rect 6276 22704 6328 22710
rect 6276 22646 6328 22652
rect 6288 22234 6316 22646
rect 6564 22574 6592 23666
rect 6932 22642 6960 23666
rect 7288 23044 7340 23050
rect 7288 22986 7340 22992
rect 7300 22778 7328 22986
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6276 22228 6328 22234
rect 6276 22170 6328 22176
rect 6828 22092 6880 22098
rect 6932 22094 6960 22578
rect 7668 22438 7696 25910
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 7748 24200 7800 24206
rect 7748 24142 7800 24148
rect 7760 23866 7788 24142
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7656 22432 7708 22438
rect 7656 22374 7708 22380
rect 7104 22094 7156 22098
rect 6932 22092 7156 22094
rect 6932 22066 7104 22092
rect 6828 22034 6880 22040
rect 7104 22034 7156 22040
rect 6840 21962 6868 22034
rect 7300 22030 7328 22374
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 6828 21956 6880 21962
rect 6828 21898 6880 21904
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5552 21690 5580 21830
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5552 21146 5580 21626
rect 6472 21554 6500 21830
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 6104 21010 6132 21286
rect 6932 21010 6960 21490
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7024 21010 7052 21082
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 7116 20942 7144 21830
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 7484 20942 7512 21286
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 4804 20868 4856 20874
rect 4804 20810 4856 20816
rect 1688 20398 1716 20810
rect 2976 20618 3004 20810
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 2976 20590 3096 20618
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1768 19780 1820 19786
rect 1768 19722 1820 19728
rect 1780 19446 1808 19722
rect 1964 19446 1992 19994
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 1768 19440 1820 19446
rect 1768 19382 1820 19388
rect 1952 19440 2004 19446
rect 1952 19382 2004 19388
rect 2332 19310 2360 19654
rect 2424 19514 2452 19790
rect 2608 19718 2636 19790
rect 2976 19718 3004 20334
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 1412 18834 1440 19246
rect 1400 18828 1452 18834
rect 1452 18788 1532 18816
rect 1400 18770 1452 18776
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 17785 1440 18022
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1504 17678 1532 18788
rect 1676 18692 1728 18698
rect 1676 18634 1728 18640
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17882 1624 18226
rect 1688 18222 1716 18634
rect 2608 18222 2636 19654
rect 2976 19514 3004 19654
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 3068 19446 3096 20590
rect 3160 20466 3188 20742
rect 4816 20602 4844 20810
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4804 20596 4856 20602
rect 4804 20538 4856 20544
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3160 19786 3188 20402
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 3148 19780 3200 19786
rect 3148 19722 3200 19728
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3056 19440 3108 19446
rect 3056 19382 3108 19388
rect 3068 18698 3096 19382
rect 3896 18766 3924 19722
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3988 19378 4016 19654
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3056 18692 3108 18698
rect 3056 18634 3108 18640
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1504 17202 1532 17614
rect 3068 17202 3096 18634
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3160 18290 3188 18566
rect 3988 18426 4016 19314
rect 4080 19174 4108 19994
rect 4816 19378 4844 20538
rect 6380 20398 6408 20878
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6656 20534 6684 20742
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 6380 19378 6408 20334
rect 6840 19446 6868 20538
rect 6828 19440 6880 19446
rect 6828 19382 6880 19388
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 4632 19258 4660 19314
rect 4632 19230 4752 19258
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4080 18834 4108 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4252 18692 4304 18698
rect 4252 18634 4304 18640
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 4264 18154 4292 18634
rect 4540 18426 4568 18770
rect 4632 18698 4660 19110
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17678 4660 18022
rect 4724 17882 4752 19230
rect 6840 18714 6868 19382
rect 6748 18698 6868 18714
rect 6736 18692 6868 18698
rect 6788 18686 6868 18692
rect 6736 18634 6788 18640
rect 6932 18630 6960 19382
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3436 17270 3464 17478
rect 3424 17264 3476 17270
rect 3424 17206 3476 17212
rect 3792 17264 3844 17270
rect 3896 17252 3924 17614
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4356 17270 4384 17478
rect 3844 17224 3924 17252
rect 3792 17206 3844 17212
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 1504 16574 1532 17138
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1964 16794 1992 17070
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 1412 16546 1532 16574
rect 1412 15502 1440 16546
rect 2240 16114 2268 16594
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15570 1716 15846
rect 1676 15564 1728 15570
rect 1676 15506 1728 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1306 14376 1362 14385
rect 1306 14311 1362 14320
rect 1320 14074 1348 14311
rect 1308 14068 1360 14074
rect 1308 14010 1360 14016
rect 1412 13394 1440 15438
rect 3068 15434 3096 17138
rect 3436 16998 3464 17206
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3436 16590 3464 16934
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3436 16250 3464 16526
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3896 16114 3924 17224
rect 4344 17264 4396 17270
rect 4344 17206 4396 17212
rect 4540 16998 4568 17614
rect 4632 17338 4660 17614
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4724 17338 4752 17546
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4448 16590 4476 16730
rect 4632 16658 4660 17274
rect 4724 17134 4752 17274
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3160 15434 3188 15914
rect 3436 15706 3464 16050
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1688 13938 1716 14418
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1872 13394 1900 14418
rect 2964 14340 3016 14346
rect 2964 14282 3016 14288
rect 2976 14074 3004 14282
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3068 14006 3096 15370
rect 3160 15094 3188 15370
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3160 14278 3188 15030
rect 3252 14414 3280 15030
rect 3344 14822 3372 15302
rect 3528 15162 3556 15438
rect 3712 15366 3740 16050
rect 3896 15706 3924 16050
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3988 15314 4016 16526
rect 4080 16250 4108 16526
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4080 15502 4108 15982
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4068 15360 4120 15366
rect 3988 15308 4068 15314
rect 3988 15302 4120 15308
rect 3988 15286 4108 15302
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3344 14346 3372 14758
rect 3528 14414 3556 15098
rect 4080 15094 4108 15286
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14482 4660 16594
rect 4724 16454 4752 17070
rect 4816 16726 4844 18566
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4908 17746 4936 18362
rect 5276 18358 5304 18566
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 5092 17678 5120 18090
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5276 17542 5304 18294
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 16794 5304 17478
rect 5644 17270 5672 18566
rect 6840 17610 6868 18566
rect 7668 18358 7696 22374
rect 8036 21690 8064 23666
rect 8312 23118 8340 24686
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 8404 22438 8432 26930
rect 8944 26784 8996 26790
rect 8944 26726 8996 26732
rect 8956 26586 8984 26726
rect 8944 26580 8996 26586
rect 8944 26522 8996 26528
rect 8956 26382 8984 26522
rect 9140 26518 9168 27406
rect 9600 27062 9628 27406
rect 9588 27056 9640 27062
rect 9588 26998 9640 27004
rect 10048 27056 10100 27062
rect 10048 26998 10100 27004
rect 9496 26988 9548 26994
rect 9496 26930 9548 26936
rect 9128 26512 9180 26518
rect 9128 26454 9180 26460
rect 9220 26512 9272 26518
rect 9220 26454 9272 26460
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 8668 25968 8720 25974
rect 8668 25910 8720 25916
rect 8680 24886 8708 25910
rect 9232 25838 9260 26454
rect 9508 25838 9536 26930
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9692 26042 9720 26318
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 9876 25922 9904 26862
rect 10060 26738 10088 26998
rect 10152 26926 10180 27406
rect 10140 26920 10192 26926
rect 10140 26862 10192 26868
rect 10060 26710 10180 26738
rect 10152 26382 10180 26710
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 10152 26042 10180 26318
rect 10140 26036 10192 26042
rect 10140 25978 10192 25984
rect 9876 25894 10088 25922
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 8668 24880 8720 24886
rect 8668 24822 8720 24828
rect 9508 23866 9536 25774
rect 9496 23860 9548 23866
rect 9496 23802 9548 23808
rect 9220 23792 9272 23798
rect 9220 23734 9272 23740
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8588 22778 8616 23666
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 8680 22778 8708 23462
rect 8772 23322 8800 23666
rect 9128 23520 9180 23526
rect 9128 23462 9180 23468
rect 8760 23316 8812 23322
rect 8760 23258 8812 23264
rect 9140 23118 9168 23462
rect 9232 23322 9260 23734
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9692 23322 9720 23462
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 9140 22710 9168 23054
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 9232 22658 9260 23258
rect 9496 23248 9548 23254
rect 9496 23190 9548 23196
rect 9508 23050 9536 23190
rect 9692 23118 9720 23258
rect 9784 23254 9812 23666
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9784 23118 9812 23190
rect 9876 23118 9904 25894
rect 10060 25838 10088 25894
rect 10048 25832 10100 25838
rect 10048 25774 10100 25780
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 10060 25294 10088 25638
rect 10140 25492 10192 25498
rect 10140 25434 10192 25440
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9956 25220 10008 25226
rect 9956 25162 10008 25168
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 8392 22432 8444 22438
rect 8392 22374 8444 22380
rect 8220 22030 8248 22374
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8024 21684 8076 21690
rect 8024 21626 8076 21632
rect 8036 21350 8064 21626
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8208 21412 8260 21418
rect 8208 21354 8260 21360
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 7932 21072 7984 21078
rect 7852 21020 7932 21026
rect 7852 21014 7984 21020
rect 7852 20998 7972 21014
rect 7852 20806 7880 20998
rect 8036 20942 8064 21286
rect 8220 21010 8248 21354
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 8024 20936 8076 20942
rect 8024 20878 8076 20884
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7760 18834 7788 20266
rect 7852 20058 7880 20742
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7944 19786 7972 20878
rect 8220 20602 8248 20946
rect 8312 20942 8340 21082
rect 8772 21010 8800 21558
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9048 21350 9076 21490
rect 9140 21486 9168 22646
rect 9232 22642 9444 22658
rect 9232 22636 9456 22642
rect 9232 22630 9404 22636
rect 9404 22578 9456 22584
rect 9692 22166 9720 23054
rect 9784 22438 9812 23054
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 9048 21162 9076 21286
rect 9048 21134 9168 21162
rect 9140 21078 9168 21134
rect 9128 21072 9180 21078
rect 9128 21014 9180 21020
rect 8760 21004 8812 21010
rect 8760 20946 8812 20952
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8312 20602 8340 20742
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 8128 20058 8156 20402
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 7932 19780 7984 19786
rect 7932 19722 7984 19728
rect 8036 19514 8064 19994
rect 8220 19854 8248 20538
rect 8772 20398 8800 20946
rect 9140 20806 9168 21014
rect 9324 21010 9352 21354
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 9600 20942 9628 21558
rect 9692 20942 9720 21626
rect 9876 21078 9904 23054
rect 9968 21690 9996 25162
rect 10152 23866 10180 25434
rect 10244 25362 10272 28970
rect 11532 28082 11560 29582
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11808 29306 11836 29514
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 13004 29238 13032 29990
rect 13280 29646 13308 30262
rect 13740 30054 13768 30534
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13740 29646 13768 29990
rect 13832 29714 13860 31214
rect 15304 30802 15332 31758
rect 15948 31686 15976 32302
rect 16408 31770 16436 32438
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 17052 32026 17080 32370
rect 17408 32360 17460 32366
rect 17408 32302 17460 32308
rect 17040 32020 17092 32026
rect 17040 31962 17092 31968
rect 16316 31742 16436 31770
rect 16316 31686 16344 31742
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 16304 31680 16356 31686
rect 16304 31622 16356 31628
rect 15948 31482 15976 31622
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 16316 31414 16344 31622
rect 17052 31482 17080 31962
rect 17040 31476 17092 31482
rect 17040 31418 17092 31424
rect 16304 31408 16356 31414
rect 16304 31350 16356 31356
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 15292 30796 15344 30802
rect 15292 30738 15344 30744
rect 15304 30326 15332 30738
rect 16040 30666 16068 31078
rect 16316 30666 16344 31350
rect 17420 31278 17448 32302
rect 19076 32230 19104 32846
rect 19524 32768 19576 32774
rect 19524 32710 19576 32716
rect 19536 32502 19564 32710
rect 20364 32502 20392 33526
rect 20640 33522 20668 33798
rect 21468 33522 21496 34342
rect 21548 33992 21600 33998
rect 21548 33934 21600 33940
rect 21560 33590 21588 33934
rect 22112 33930 22140 34342
rect 22100 33924 22152 33930
rect 22100 33866 22152 33872
rect 22192 33856 22244 33862
rect 22192 33798 22244 33804
rect 21548 33584 21600 33590
rect 21548 33526 21600 33532
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 21456 33516 21508 33522
rect 21456 33458 21508 33464
rect 21088 33312 21140 33318
rect 21088 33254 21140 33260
rect 21100 32978 21128 33254
rect 21088 32972 21140 32978
rect 21088 32914 21140 32920
rect 22204 32910 22232 33798
rect 22572 33658 22600 34478
rect 23492 34202 23520 34546
rect 23480 34196 23532 34202
rect 23480 34138 23532 34144
rect 22560 33652 22612 33658
rect 22560 33594 22612 33600
rect 22284 33448 22336 33454
rect 22284 33390 22336 33396
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 19524 32496 19576 32502
rect 19524 32438 19576 32444
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 22100 32360 22152 32366
rect 22100 32302 22152 32308
rect 19064 32224 19116 32230
rect 19064 32166 19116 32172
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 19076 31890 19104 32166
rect 21008 31890 21036 32166
rect 19064 31884 19116 31890
rect 19064 31826 19116 31832
rect 20996 31884 21048 31890
rect 20996 31826 21048 31832
rect 18880 31748 18932 31754
rect 18880 31690 18932 31696
rect 18892 31414 18920 31690
rect 19076 31482 19104 31826
rect 22112 31482 22140 32302
rect 22204 31890 22232 32846
rect 22296 32570 22324 33390
rect 22572 33114 22600 33594
rect 22928 33448 22980 33454
rect 22928 33390 22980 33396
rect 22940 33114 22968 33390
rect 22560 33108 22612 33114
rect 22560 33050 22612 33056
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 23492 32774 23520 34138
rect 24412 33998 24440 35022
rect 24688 34678 24716 35974
rect 24780 35601 24808 36042
rect 24766 35592 24822 35601
rect 24766 35527 24822 35536
rect 24676 34672 24728 34678
rect 24676 34614 24728 34620
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24412 33522 24440 33934
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24412 32910 24440 33254
rect 24688 33046 24716 34614
rect 24872 34474 24900 36586
rect 25228 36576 25280 36582
rect 25228 36518 25280 36524
rect 24952 36304 25004 36310
rect 24952 36246 25004 36252
rect 24964 35018 24992 36246
rect 25240 35766 25268 36518
rect 25516 36378 25544 36615
rect 25976 36378 26004 36722
rect 26160 36650 26188 37198
rect 26516 37188 26568 37194
rect 26516 37130 26568 37136
rect 26528 36922 26556 37130
rect 26608 37120 26660 37126
rect 26608 37062 26660 37068
rect 26516 36916 26568 36922
rect 26516 36858 26568 36864
rect 26620 36786 26648 37062
rect 26516 36780 26568 36786
rect 26516 36722 26568 36728
rect 26608 36780 26660 36786
rect 26608 36722 26660 36728
rect 27068 36780 27120 36786
rect 27068 36722 27120 36728
rect 26148 36644 26200 36650
rect 26148 36586 26200 36592
rect 25504 36372 25556 36378
rect 25504 36314 25556 36320
rect 25964 36372 26016 36378
rect 25964 36314 26016 36320
rect 26160 36242 26188 36586
rect 26528 36378 26556 36722
rect 26516 36372 26568 36378
rect 26516 36314 26568 36320
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 26148 36236 26200 36242
rect 26148 36178 26200 36184
rect 25228 35760 25280 35766
rect 25228 35702 25280 35708
rect 25424 35630 25452 36178
rect 25780 36168 25832 36174
rect 25964 36168 26016 36174
rect 25832 36116 25964 36122
rect 25780 36110 26016 36116
rect 25792 36094 26004 36110
rect 25504 36032 25556 36038
rect 25504 35974 25556 35980
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 25148 35018 25176 35566
rect 25424 35154 25452 35566
rect 25412 35148 25464 35154
rect 25412 35090 25464 35096
rect 24952 35012 25004 35018
rect 24952 34954 25004 34960
rect 25136 35012 25188 35018
rect 25188 34972 25268 35000
rect 25136 34954 25188 34960
rect 25240 34678 25268 34972
rect 25516 34746 25544 35974
rect 25976 35290 26004 36094
rect 26240 35624 26292 35630
rect 26240 35566 26292 35572
rect 26252 35290 26280 35566
rect 27080 35562 27108 36722
rect 27264 36650 27292 37742
rect 27712 37664 27764 37670
rect 27712 37606 27764 37612
rect 27988 37664 28040 37670
rect 27988 37606 28040 37612
rect 27528 37256 27580 37262
rect 27448 37204 27528 37210
rect 27448 37198 27580 37204
rect 27448 37182 27568 37198
rect 27344 36780 27396 36786
rect 27344 36722 27396 36728
rect 27356 36650 27384 36722
rect 27252 36644 27304 36650
rect 27252 36586 27304 36592
rect 27344 36644 27396 36650
rect 27344 36586 27396 36592
rect 27264 35630 27292 36586
rect 27448 36582 27476 37182
rect 27724 36854 27752 37606
rect 27712 36848 27764 36854
rect 27712 36790 27764 36796
rect 27436 36576 27488 36582
rect 27436 36518 27488 36524
rect 27252 35624 27304 35630
rect 27252 35566 27304 35572
rect 27068 35556 27120 35562
rect 27068 35498 27120 35504
rect 27448 35494 27476 36518
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 27632 35766 27660 36178
rect 27620 35760 27672 35766
rect 27620 35702 27672 35708
rect 28000 35698 28028 37606
rect 28092 37466 28120 37810
rect 29184 37800 29236 37806
rect 29184 37742 29236 37748
rect 30380 37800 30432 37806
rect 30380 37742 30432 37748
rect 28080 37460 28132 37466
rect 28080 37402 28132 37408
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28724 37256 28776 37262
rect 28724 37198 28776 37204
rect 28264 37120 28316 37126
rect 28264 37062 28316 37068
rect 27712 35692 27764 35698
rect 27712 35634 27764 35640
rect 27988 35692 28040 35698
rect 27988 35634 28040 35640
rect 27724 35494 27752 35634
rect 27436 35488 27488 35494
rect 27436 35430 27488 35436
rect 27712 35488 27764 35494
rect 27712 35430 27764 35436
rect 25964 35284 26016 35290
rect 25964 35226 26016 35232
rect 26240 35284 26292 35290
rect 26240 35226 26292 35232
rect 28276 35170 28304 37062
rect 28552 35698 28580 37198
rect 28736 36310 28764 37198
rect 28908 37188 28960 37194
rect 28908 37130 28960 37136
rect 28920 36836 28948 37130
rect 29000 36848 29052 36854
rect 28920 36808 29000 36836
rect 28814 36680 28870 36689
rect 28814 36615 28870 36624
rect 28724 36304 28776 36310
rect 28724 36246 28776 36252
rect 28724 36168 28776 36174
rect 28724 36110 28776 36116
rect 28540 35692 28592 35698
rect 28540 35634 28592 35640
rect 28632 35216 28684 35222
rect 28276 35164 28632 35170
rect 28276 35158 28684 35164
rect 28276 35142 28672 35158
rect 25964 35012 26016 35018
rect 25964 34954 26016 34960
rect 25504 34740 25556 34746
rect 25504 34682 25556 34688
rect 25228 34672 25280 34678
rect 25228 34614 25280 34620
rect 24860 34468 24912 34474
rect 24860 34410 24912 34416
rect 25044 34400 25096 34406
rect 25044 34342 25096 34348
rect 25056 34066 25084 34342
rect 25044 34060 25096 34066
rect 25044 34002 25096 34008
rect 25136 34060 25188 34066
rect 25136 34002 25188 34008
rect 25148 33590 25176 34002
rect 25240 33930 25268 34614
rect 25228 33924 25280 33930
rect 25228 33866 25280 33872
rect 25240 33658 25268 33866
rect 25516 33862 25544 34682
rect 25976 34678 26004 34954
rect 28172 34944 28224 34950
rect 28172 34886 28224 34892
rect 25964 34672 26016 34678
rect 25964 34614 26016 34620
rect 27620 34672 27672 34678
rect 27620 34614 27672 34620
rect 27804 34672 27856 34678
rect 27804 34614 27856 34620
rect 25780 34468 25832 34474
rect 25780 34410 25832 34416
rect 25504 33856 25556 33862
rect 25504 33798 25556 33804
rect 25228 33652 25280 33658
rect 25228 33594 25280 33600
rect 25136 33584 25188 33590
rect 25136 33526 25188 33532
rect 24860 33448 24912 33454
rect 24860 33390 24912 33396
rect 24872 33114 24900 33390
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24676 33040 24728 33046
rect 24676 32982 24728 32988
rect 25148 32910 25176 33526
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 24400 32904 24452 32910
rect 24400 32846 24452 32852
rect 25136 32904 25188 32910
rect 25136 32846 25188 32852
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22296 32026 22324 32506
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 22284 32020 22336 32026
rect 22284 31962 22336 31968
rect 22192 31884 22244 31890
rect 22192 31826 22244 31832
rect 19064 31476 19116 31482
rect 19064 31418 19116 31424
rect 22100 31476 22152 31482
rect 22100 31418 22152 31424
rect 18880 31408 18932 31414
rect 18880 31350 18932 31356
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17408 31272 17460 31278
rect 17408 31214 17460 31220
rect 16396 31204 16448 31210
rect 16396 31146 16448 31152
rect 16408 30938 16436 31146
rect 16396 30932 16448 30938
rect 16396 30874 16448 30880
rect 16028 30660 16080 30666
rect 16304 30660 16356 30666
rect 16028 30602 16080 30608
rect 16224 30620 16304 30648
rect 16224 30394 16252 30620
rect 16304 30602 16356 30608
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 15292 30320 15344 30326
rect 15292 30262 15344 30268
rect 15200 30184 15252 30190
rect 15200 30126 15252 30132
rect 15212 29850 15240 30126
rect 15200 29844 15252 29850
rect 15200 29786 15252 29792
rect 13820 29708 13872 29714
rect 13820 29650 13872 29656
rect 14648 29708 14700 29714
rect 14648 29650 14700 29656
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13280 29306 13308 29446
rect 13268 29300 13320 29306
rect 13268 29242 13320 29248
rect 12992 29232 13044 29238
rect 12992 29174 13044 29180
rect 13176 29096 13228 29102
rect 13176 29038 13228 29044
rect 13188 28626 13216 29038
rect 13176 28620 13228 28626
rect 13176 28562 13228 28568
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11992 28150 12020 28358
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 11520 28076 11572 28082
rect 11520 28018 11572 28024
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 10784 27872 10836 27878
rect 10784 27814 10836 27820
rect 10600 27532 10652 27538
rect 10428 27492 10600 27520
rect 10324 27464 10376 27470
rect 10324 27406 10376 27412
rect 10336 26382 10364 27406
rect 10428 26994 10456 27492
rect 10520 27402 10548 27492
rect 10600 27474 10652 27480
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 10324 26376 10376 26382
rect 10324 26318 10376 26324
rect 10232 25356 10284 25362
rect 10232 25298 10284 25304
rect 10232 25152 10284 25158
rect 10232 25094 10284 25100
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10244 23798 10272 25094
rect 10232 23792 10284 23798
rect 10232 23734 10284 23740
rect 10336 23186 10364 26318
rect 10428 26246 10456 26930
rect 10704 26586 10732 27066
rect 10796 26790 10824 27814
rect 11716 27520 11744 28018
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 11796 27532 11848 27538
rect 11716 27492 11796 27520
rect 12452 27520 12480 27950
rect 11796 27474 11848 27480
rect 12360 27492 12480 27520
rect 12808 27532 12860 27538
rect 10876 27396 10928 27402
rect 10876 27338 10928 27344
rect 11060 27396 11112 27402
rect 11060 27338 11112 27344
rect 10888 26858 10916 27338
rect 10968 27328 11020 27334
rect 10968 27270 11020 27276
rect 10980 27062 11008 27270
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 10876 26852 10928 26858
rect 10876 26794 10928 26800
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10692 26580 10744 26586
rect 10612 26540 10692 26568
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10508 25764 10560 25770
rect 10508 25706 10560 25712
rect 10520 25498 10548 25706
rect 10508 25492 10560 25498
rect 10508 25434 10560 25440
rect 10612 25226 10640 26540
rect 10692 26522 10744 26528
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10704 25498 10732 26250
rect 10796 25974 10824 26726
rect 11072 26314 11100 27338
rect 12360 26314 12388 27492
rect 12808 27474 12860 27480
rect 12440 27396 12492 27402
rect 12440 27338 12492 27344
rect 12452 26586 12480 27338
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 11060 26308 11112 26314
rect 11060 26250 11112 26256
rect 12348 26308 12400 26314
rect 12348 26250 12400 26256
rect 10876 26240 10928 26246
rect 10876 26182 10928 26188
rect 10784 25968 10836 25974
rect 10784 25910 10836 25916
rect 10888 25838 10916 26182
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10600 25220 10652 25226
rect 10600 25162 10652 25168
rect 11072 24818 11100 26250
rect 12072 26240 12124 26246
rect 12072 26182 12124 26188
rect 12084 25906 12112 26182
rect 12820 25906 12848 27474
rect 13188 26908 13216 28562
rect 13280 28558 13308 29242
rect 14660 29102 14688 29650
rect 16224 29578 16252 30330
rect 16212 29572 16264 29578
rect 16212 29514 16264 29520
rect 15660 29504 15712 29510
rect 15660 29446 15712 29452
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 15672 29306 15700 29446
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 14188 29096 14240 29102
rect 14188 29038 14240 29044
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14200 28762 14228 29038
rect 14740 28960 14792 28966
rect 14740 28902 14792 28908
rect 14188 28756 14240 28762
rect 14188 28698 14240 28704
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 13452 28416 13504 28422
rect 13452 28358 13504 28364
rect 13464 27878 13492 28358
rect 13728 28144 13780 28150
rect 13728 28086 13780 28092
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 13360 27328 13412 27334
rect 13360 27270 13412 27276
rect 13372 27130 13400 27270
rect 13360 27124 13412 27130
rect 13360 27066 13412 27072
rect 13268 26920 13320 26926
rect 13188 26880 13268 26908
rect 13268 26862 13320 26868
rect 13280 26518 13308 26862
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 13372 26382 13400 27066
rect 13464 26450 13492 27814
rect 13740 27402 13768 28086
rect 14752 28014 14780 28902
rect 15672 28558 15700 29242
rect 15764 29170 15792 29446
rect 16224 29238 16252 29514
rect 16212 29232 16264 29238
rect 16212 29174 16264 29180
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15660 28552 15712 28558
rect 15660 28494 15712 28500
rect 15764 28490 15792 29106
rect 16224 28506 16252 29174
rect 16408 28626 16436 30874
rect 16488 30796 16540 30802
rect 16488 30738 16540 30744
rect 16500 29714 16528 30738
rect 17592 30660 17644 30666
rect 17592 30602 17644 30608
rect 17604 30394 17632 30602
rect 17972 30598 18000 31282
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 18340 30938 18368 31214
rect 18328 30932 18380 30938
rect 18328 30874 18380 30880
rect 18236 30796 18288 30802
rect 18236 30738 18288 30744
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 18248 30394 18276 30738
rect 18892 30666 18920 31350
rect 19076 31278 19104 31418
rect 19064 31272 19116 31278
rect 19064 31214 19116 31220
rect 20168 31272 20220 31278
rect 20168 31214 20220 31220
rect 19340 31136 19392 31142
rect 19340 31078 19392 31084
rect 19616 31136 19668 31142
rect 19616 31078 19668 31084
rect 19352 30870 19380 31078
rect 19340 30864 19392 30870
rect 19340 30806 19392 30812
rect 19628 30734 19656 31078
rect 20180 30938 20208 31214
rect 20168 30932 20220 30938
rect 20168 30874 20220 30880
rect 20260 30864 20312 30870
rect 20260 30806 20312 30812
rect 19616 30728 19668 30734
rect 19616 30670 19668 30676
rect 18880 30660 18932 30666
rect 18880 30602 18932 30608
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 18340 30394 18368 30534
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 18236 30388 18288 30394
rect 18236 30330 18288 30336
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18420 30184 18472 30190
rect 18420 30126 18472 30132
rect 16488 29708 16540 29714
rect 16488 29650 16540 29656
rect 17224 29572 17276 29578
rect 17224 29514 17276 29520
rect 17236 29306 17264 29514
rect 17224 29300 17276 29306
rect 17224 29242 17276 29248
rect 17316 29164 17368 29170
rect 17316 29106 17368 29112
rect 16856 29096 16908 29102
rect 16856 29038 16908 29044
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 16132 28478 16252 28506
rect 16132 28082 16160 28478
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 14740 28008 14792 28014
rect 14740 27950 14792 27956
rect 14752 27520 14780 27950
rect 16132 27878 16160 28018
rect 16304 28008 16356 28014
rect 16304 27950 16356 27956
rect 15200 27872 15252 27878
rect 15200 27814 15252 27820
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 15212 27690 15240 27814
rect 15120 27662 15240 27690
rect 14832 27532 14884 27538
rect 14752 27492 14832 27520
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 14108 26926 14136 27270
rect 14752 27062 14780 27492
rect 14832 27474 14884 27480
rect 15120 27402 15148 27662
rect 16316 27606 16344 27950
rect 16408 27606 16436 28562
rect 16868 28218 16896 29038
rect 17328 28762 17356 29106
rect 18432 29034 18460 30126
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 17960 29028 18012 29034
rect 17960 28970 18012 28976
rect 18420 29028 18472 29034
rect 18420 28970 18472 28976
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16672 27872 16724 27878
rect 16672 27814 16724 27820
rect 16304 27600 16356 27606
rect 16304 27542 16356 27548
rect 16396 27600 16448 27606
rect 16448 27548 16528 27554
rect 16396 27542 16528 27548
rect 16408 27526 16528 27542
rect 16684 27538 16712 27814
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 15108 27396 15160 27402
rect 15108 27338 15160 27344
rect 15568 27396 15620 27402
rect 15568 27338 15620 27344
rect 15580 27130 15608 27338
rect 15568 27124 15620 27130
rect 15568 27066 15620 27072
rect 14740 27056 14792 27062
rect 14740 26998 14792 27004
rect 16408 26994 16436 27406
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 14096 26920 14148 26926
rect 14096 26862 14148 26868
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 14108 26450 14136 26862
rect 13452 26444 13504 26450
rect 13452 26386 13504 26392
rect 14096 26444 14148 26450
rect 14096 26386 14148 26392
rect 14740 26444 14792 26450
rect 14740 26386 14792 26392
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 13544 26308 13596 26314
rect 13544 26250 13596 26256
rect 13556 25974 13584 26250
rect 14096 26240 14148 26246
rect 14096 26182 14148 26188
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 13544 25968 13596 25974
rect 13544 25910 13596 25916
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 14108 25838 14136 26182
rect 14476 26042 14504 26182
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 14476 25430 14504 25978
rect 14464 25424 14516 25430
rect 14464 25366 14516 25372
rect 14752 25362 14780 26386
rect 14936 26382 14964 26862
rect 16408 26450 16436 26930
rect 16500 26858 16528 27526
rect 16672 27532 16724 27538
rect 16672 27474 16724 27480
rect 16868 27402 16896 28154
rect 17328 27402 17356 28698
rect 17972 27538 18000 28970
rect 18788 28960 18840 28966
rect 18788 28902 18840 28908
rect 18800 28626 18828 28902
rect 19260 28626 19288 29582
rect 19524 29572 19576 29578
rect 19524 29514 19576 29520
rect 19536 29306 19564 29514
rect 20168 29504 20220 29510
rect 20168 29446 20220 29452
rect 20180 29306 20208 29446
rect 19524 29300 19576 29306
rect 19524 29242 19576 29248
rect 20168 29300 20220 29306
rect 20168 29242 20220 29248
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 18788 28620 18840 28626
rect 18788 28562 18840 28568
rect 19248 28620 19300 28626
rect 19248 28562 19300 28568
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 18328 28484 18380 28490
rect 18328 28426 18380 28432
rect 18236 28144 18288 28150
rect 18340 28132 18368 28426
rect 18288 28104 18368 28132
rect 18236 28086 18288 28092
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18156 27674 18184 27950
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 17960 27532 18012 27538
rect 17960 27474 18012 27480
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 17316 27396 17368 27402
rect 17316 27338 17368 27344
rect 17040 26920 17092 26926
rect 17040 26862 17092 26868
rect 17776 26920 17828 26926
rect 17776 26862 17828 26868
rect 16488 26852 16540 26858
rect 16488 26794 16540 26800
rect 16500 26518 16528 26794
rect 16488 26512 16540 26518
rect 16488 26454 16540 26460
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10428 23322 10456 23462
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 10060 22778 10088 22986
rect 10520 22778 10548 23666
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9968 21146 9996 21422
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 9128 20800 9180 20806
rect 9128 20742 9180 20748
rect 8956 20466 8984 20742
rect 9600 20602 9628 20878
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 8772 18970 8800 20334
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 9416 18698 9444 19382
rect 9692 19310 9720 20266
rect 9784 19922 9812 20742
rect 9968 20618 9996 21082
rect 10060 21010 10088 21966
rect 10428 21690 10456 22578
rect 10520 22166 10548 22578
rect 10612 22234 10640 23462
rect 10704 22642 10732 23802
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10888 22982 10916 23598
rect 11072 23050 11100 24754
rect 11808 24274 11836 25230
rect 13820 25220 13872 25226
rect 13820 25162 13872 25168
rect 13832 24750 13860 25162
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 14016 24954 14044 25094
rect 14004 24948 14056 24954
rect 14004 24890 14056 24896
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13820 24744 13872 24750
rect 13820 24686 13872 24692
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 13096 24274 13124 24550
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 12164 24268 12216 24274
rect 12164 24210 12216 24216
rect 13084 24268 13136 24274
rect 13084 24210 13136 24216
rect 12176 23186 12204 24210
rect 13832 24138 13860 24686
rect 13924 24410 13952 24754
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12452 23186 12480 23462
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 11060 23044 11112 23050
rect 11060 22986 11112 22992
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10784 22704 10836 22710
rect 10784 22646 10836 22652
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10796 22438 10824 22646
rect 10888 22642 10916 22918
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10508 22160 10560 22166
rect 10508 22102 10560 22108
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10336 21010 10364 21286
rect 10428 21146 10456 21626
rect 10796 21486 10824 22374
rect 11072 21962 11100 22986
rect 12176 22642 12204 23122
rect 13832 23050 13860 24074
rect 13924 23866 13952 24346
rect 14476 24206 14504 25230
rect 14752 24750 14780 25298
rect 14936 25294 14964 26318
rect 17052 26042 17080 26862
rect 17224 26784 17276 26790
rect 17224 26726 17276 26732
rect 17040 26036 17092 26042
rect 17040 25978 17092 25984
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16948 25832 17000 25838
rect 16948 25774 17000 25780
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 15200 25220 15252 25226
rect 15200 25162 15252 25168
rect 15844 25220 15896 25226
rect 15844 25162 15896 25168
rect 15212 24954 15240 25162
rect 15200 24948 15252 24954
rect 15200 24890 15252 24896
rect 14740 24744 14792 24750
rect 14660 24692 14740 24698
rect 14660 24686 14792 24692
rect 14660 24670 14780 24686
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13924 23322 13952 23666
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13832 22710 13860 22986
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 14016 22574 14044 22918
rect 14476 22778 14504 24142
rect 14660 23186 14688 24670
rect 15856 24206 15884 25162
rect 16868 24750 16896 25774
rect 16960 25498 16988 25774
rect 16948 25492 17000 25498
rect 16948 25434 17000 25440
rect 16960 24954 16988 25434
rect 17236 25362 17264 26726
rect 17788 26586 17816 26862
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17408 26308 17460 26314
rect 17408 26250 17460 26256
rect 17420 26042 17448 26250
rect 17408 26036 17460 26042
rect 17408 25978 17460 25984
rect 17972 25974 18000 26726
rect 18340 26246 18368 28104
rect 19260 28014 19288 28562
rect 19352 28014 19380 28562
rect 19904 28490 19932 29106
rect 20180 28490 20208 29242
rect 20272 29102 20300 30806
rect 20904 30796 20956 30802
rect 20904 30738 20956 30744
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20824 29646 20852 30534
rect 20916 30190 20944 30738
rect 22112 30666 22140 31418
rect 22204 31414 22232 31826
rect 22192 31408 22244 31414
rect 22192 31350 22244 31356
rect 22100 30660 22152 30666
rect 22100 30602 22152 30608
rect 22204 30326 22232 31350
rect 22480 30938 22508 32302
rect 23584 31890 23612 32846
rect 24860 32496 24912 32502
rect 24860 32438 24912 32444
rect 23572 31884 23624 31890
rect 23572 31826 23624 31832
rect 24768 31884 24820 31890
rect 24768 31826 24820 31832
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24492 31680 24544 31686
rect 24492 31622 24544 31628
rect 22572 31414 22600 31622
rect 24412 31414 24440 31622
rect 24504 31482 24532 31622
rect 24492 31476 24544 31482
rect 24492 31418 24544 31424
rect 22560 31408 22612 31414
rect 22560 31350 22612 31356
rect 24400 31408 24452 31414
rect 24400 31350 24452 31356
rect 24400 31272 24452 31278
rect 24400 31214 24452 31220
rect 22468 30932 22520 30938
rect 22468 30874 22520 30880
rect 24412 30734 24440 31214
rect 24400 30728 24452 30734
rect 24400 30670 24452 30676
rect 22192 30320 22244 30326
rect 22192 30262 22244 30268
rect 20904 30184 20956 30190
rect 20904 30126 20956 30132
rect 20916 29714 20944 30126
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20720 28960 20772 28966
rect 20720 28902 20772 28908
rect 20732 28626 20760 28902
rect 20720 28620 20772 28626
rect 20720 28562 20772 28568
rect 20824 28490 20852 29582
rect 20916 29102 20944 29650
rect 22204 29646 22232 30262
rect 24412 30258 24440 30670
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 22560 30048 22612 30054
rect 22560 29990 22612 29996
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22204 29306 22232 29582
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 21272 29164 21324 29170
rect 21272 29106 21324 29112
rect 20904 29096 20956 29102
rect 20904 29038 20956 29044
rect 21284 28762 21312 29106
rect 21456 29096 21508 29102
rect 21456 29038 21508 29044
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 21468 28626 21496 29038
rect 22572 28626 22600 29990
rect 23296 29572 23348 29578
rect 23296 29514 23348 29520
rect 22652 29504 22704 29510
rect 22652 29446 22704 29452
rect 22664 29170 22692 29446
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 21456 28620 21508 28626
rect 21456 28562 21508 28568
rect 22560 28620 22612 28626
rect 22560 28562 22612 28568
rect 19892 28484 19944 28490
rect 19892 28426 19944 28432
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 19524 28416 19576 28422
rect 19524 28358 19576 28364
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19260 27538 19288 27950
rect 19352 27674 19380 27950
rect 19536 27674 19564 28358
rect 19904 27674 19932 28426
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19524 27668 19576 27674
rect 19524 27610 19576 27616
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 18880 27532 18932 27538
rect 18880 27474 18932 27480
rect 19248 27532 19300 27538
rect 19248 27474 19300 27480
rect 18892 26926 18920 27474
rect 19260 26994 19288 27474
rect 20824 27402 20852 28426
rect 22572 28422 22600 28562
rect 22664 28558 22692 29106
rect 23308 28762 23336 29514
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23296 28756 23348 28762
rect 23296 28698 23348 28704
rect 23492 28558 23520 29242
rect 23676 28762 23704 30126
rect 24780 29782 24808 31826
rect 24872 30122 24900 32438
rect 25240 31822 25268 33594
rect 25792 32978 25820 34410
rect 25976 33930 26004 34614
rect 26148 34604 26200 34610
rect 26148 34546 26200 34552
rect 25964 33924 26016 33930
rect 25964 33866 26016 33872
rect 26160 33658 26188 34546
rect 26148 33652 26200 33658
rect 26148 33594 26200 33600
rect 26056 33448 26108 33454
rect 26056 33390 26108 33396
rect 25780 32972 25832 32978
rect 25780 32914 25832 32920
rect 25688 32768 25740 32774
rect 25688 32710 25740 32716
rect 25700 31890 25728 32710
rect 25792 32570 25820 32914
rect 26068 32910 26096 33390
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26160 32842 26188 33594
rect 26148 32836 26200 32842
rect 26148 32778 26200 32784
rect 25780 32564 25832 32570
rect 25780 32506 25832 32512
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26068 32026 26096 32370
rect 27632 32026 27660 34614
rect 27712 33516 27764 33522
rect 27712 33458 27764 33464
rect 27724 32502 27752 33458
rect 27816 33046 27844 34614
rect 28184 34542 28212 34886
rect 28276 34542 28304 35142
rect 28736 35086 28764 36110
rect 28828 36106 28856 36615
rect 28816 36100 28868 36106
rect 28816 36042 28868 36048
rect 28828 35086 28856 36042
rect 28920 36038 28948 36808
rect 29000 36790 29052 36796
rect 29196 36378 29224 37742
rect 29828 37256 29880 37262
rect 29828 37198 29880 37204
rect 29736 37188 29788 37194
rect 29736 37130 29788 37136
rect 29748 36786 29776 37130
rect 29840 37126 29868 37198
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 29736 36780 29788 36786
rect 29736 36722 29788 36728
rect 29552 36712 29604 36718
rect 29552 36654 29604 36660
rect 29564 36378 29592 36654
rect 29184 36372 29236 36378
rect 29184 36314 29236 36320
rect 29552 36372 29604 36378
rect 29552 36314 29604 36320
rect 28908 36032 28960 36038
rect 28908 35974 28960 35980
rect 29000 36032 29052 36038
rect 29000 35974 29052 35980
rect 28448 35080 28500 35086
rect 28448 35022 28500 35028
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 28816 35080 28868 35086
rect 28816 35022 28868 35028
rect 28460 34746 28488 35022
rect 28448 34740 28500 34746
rect 28448 34682 28500 34688
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 28172 34536 28224 34542
rect 28172 34478 28224 34484
rect 28264 34536 28316 34542
rect 28264 34478 28316 34484
rect 28184 34202 28212 34478
rect 28172 34196 28224 34202
rect 28172 34138 28224 34144
rect 28540 34060 28592 34066
rect 28540 34002 28592 34008
rect 28080 33312 28132 33318
rect 28080 33254 28132 33260
rect 27804 33040 27856 33046
rect 27804 32982 27856 32988
rect 27712 32496 27764 32502
rect 27896 32496 27948 32502
rect 27712 32438 27764 32444
rect 27816 32456 27896 32484
rect 26056 32020 26108 32026
rect 26056 31962 26108 31968
rect 27620 32020 27672 32026
rect 27620 31962 27672 31968
rect 25688 31884 25740 31890
rect 25688 31826 25740 31832
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25240 31396 25268 31758
rect 25780 31748 25832 31754
rect 25780 31690 25832 31696
rect 25792 31482 25820 31690
rect 25780 31476 25832 31482
rect 25780 31418 25832 31424
rect 25320 31408 25372 31414
rect 25240 31368 25320 31396
rect 25240 30666 25268 31368
rect 25320 31350 25372 31356
rect 26068 31278 26096 31962
rect 26976 31884 27028 31890
rect 26976 31826 27028 31832
rect 26988 31754 27016 31826
rect 26976 31748 27028 31754
rect 26976 31690 27028 31696
rect 27528 31408 27580 31414
rect 27528 31350 27580 31356
rect 27712 31408 27764 31414
rect 27816 31396 27844 32456
rect 27896 32438 27948 32444
rect 28092 32366 28120 33254
rect 28552 33114 28580 34002
rect 28540 33108 28592 33114
rect 28540 33050 28592 33056
rect 28816 33108 28868 33114
rect 28816 33050 28868 33056
rect 28828 32774 28856 33050
rect 28920 32842 28948 34546
rect 29012 34542 29040 35974
rect 29196 35086 29224 36314
rect 29564 36242 29592 36314
rect 29552 36236 29604 36242
rect 29552 36178 29604 36184
rect 29368 36168 29420 36174
rect 29368 36110 29420 36116
rect 29380 35494 29408 36110
rect 29840 35698 29868 37062
rect 30392 36786 30420 37742
rect 30472 37324 30524 37330
rect 30472 37266 30524 37272
rect 30564 37324 30616 37330
rect 30564 37266 30616 37272
rect 30380 36780 30432 36786
rect 30380 36722 30432 36728
rect 30104 36576 30156 36582
rect 30104 36518 30156 36524
rect 29920 36372 29972 36378
rect 29920 36314 29972 36320
rect 29736 35692 29788 35698
rect 29736 35634 29788 35640
rect 29828 35692 29880 35698
rect 29828 35634 29880 35640
rect 29368 35488 29420 35494
rect 29368 35430 29420 35436
rect 29184 35080 29236 35086
rect 29184 35022 29236 35028
rect 29092 35012 29144 35018
rect 29092 34954 29144 34960
rect 29104 34542 29132 34954
rect 29380 34610 29408 35430
rect 29748 35290 29776 35634
rect 29736 35284 29788 35290
rect 29736 35226 29788 35232
rect 29460 34672 29512 34678
rect 29460 34614 29512 34620
rect 29368 34604 29420 34610
rect 29368 34546 29420 34552
rect 29000 34536 29052 34542
rect 29000 34478 29052 34484
rect 29092 34536 29144 34542
rect 29092 34478 29144 34484
rect 29276 34536 29328 34542
rect 29276 34478 29328 34484
rect 29184 34060 29236 34066
rect 29184 34002 29236 34008
rect 29092 33448 29144 33454
rect 29092 33390 29144 33396
rect 29000 33312 29052 33318
rect 29000 33254 29052 33260
rect 29012 32978 29040 33254
rect 29000 32972 29052 32978
rect 29000 32914 29052 32920
rect 29104 32858 29132 33390
rect 29196 32910 29224 34002
rect 29288 33998 29316 34478
rect 29380 34134 29408 34546
rect 29368 34128 29420 34134
rect 29368 34070 29420 34076
rect 29276 33992 29328 33998
rect 29276 33934 29328 33940
rect 29368 33992 29420 33998
rect 29368 33934 29420 33940
rect 29380 33522 29408 33934
rect 29472 33522 29500 34614
rect 29736 34536 29788 34542
rect 29736 34478 29788 34484
rect 29644 33924 29696 33930
rect 29644 33866 29696 33872
rect 29656 33522 29684 33866
rect 29368 33516 29420 33522
rect 29368 33458 29420 33464
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 29644 33516 29696 33522
rect 29644 33458 29696 33464
rect 29644 33040 29696 33046
rect 29644 32982 29696 32988
rect 28908 32836 28960 32842
rect 28908 32778 28960 32784
rect 29012 32830 29132 32858
rect 29184 32904 29236 32910
rect 29184 32846 29236 32852
rect 28816 32768 28868 32774
rect 28816 32710 28868 32716
rect 29012 32570 29040 32830
rect 29000 32564 29052 32570
rect 29000 32506 29052 32512
rect 29184 32496 29236 32502
rect 29184 32438 29236 32444
rect 28080 32360 28132 32366
rect 28080 32302 28132 32308
rect 27988 31884 28040 31890
rect 27988 31826 28040 31832
rect 27896 31680 27948 31686
rect 27896 31622 27948 31628
rect 27764 31368 27844 31396
rect 27712 31350 27764 31356
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 26056 31272 26108 31278
rect 26056 31214 26108 31220
rect 25228 30660 25280 30666
rect 25228 30602 25280 30608
rect 25044 30184 25096 30190
rect 25044 30126 25096 30132
rect 24860 30116 24912 30122
rect 24860 30058 24912 30064
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24780 29306 24808 29446
rect 24768 29300 24820 29306
rect 24768 29242 24820 29248
rect 23848 29232 23900 29238
rect 23848 29174 23900 29180
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 23480 28552 23532 28558
rect 23480 28494 23532 28500
rect 23860 28490 23888 29174
rect 23848 28484 23900 28490
rect 23848 28426 23900 28432
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22664 27538 22692 28018
rect 22652 27532 22704 27538
rect 22652 27474 22704 27480
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 22192 27396 22244 27402
rect 22192 27338 22244 27344
rect 20444 27328 20496 27334
rect 20444 27270 20496 27276
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18880 26920 18932 26926
rect 18880 26862 18932 26868
rect 18328 26240 18380 26246
rect 18328 26182 18380 26188
rect 17960 25968 18012 25974
rect 17960 25910 18012 25916
rect 18512 25832 18564 25838
rect 18512 25774 18564 25780
rect 17224 25356 17276 25362
rect 17224 25298 17276 25304
rect 18524 25226 18552 25774
rect 18800 25498 18828 26862
rect 18892 26042 18920 26862
rect 19260 26450 19288 26930
rect 19248 26444 19300 26450
rect 19248 26386 19300 26392
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 18880 26036 18932 26042
rect 18880 25978 18932 25984
rect 19260 25974 19288 26250
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 18788 25492 18840 25498
rect 18788 25434 18840 25440
rect 19260 25294 19288 25910
rect 19444 25702 19472 27066
rect 20456 27062 20484 27270
rect 20824 27130 20852 27338
rect 22100 27328 22152 27334
rect 22100 27270 22152 27276
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 20444 27056 20496 27062
rect 20444 26998 20496 27004
rect 20720 27056 20772 27062
rect 20824 27010 20852 27066
rect 20772 27004 20852 27010
rect 20720 26998 20852 27004
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 18512 25220 18564 25226
rect 18512 25162 18564 25168
rect 16948 24948 17000 24954
rect 16948 24890 17000 24896
rect 18524 24818 18552 25162
rect 19260 24886 19288 25230
rect 20364 25226 20392 25842
rect 20456 25294 20484 26998
rect 20732 26982 20852 26998
rect 20732 26314 20760 26982
rect 21836 26790 21864 27066
rect 22112 26926 22140 27270
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 21824 26784 21876 26790
rect 21824 26726 21876 26732
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20352 25220 20404 25226
rect 20352 25162 20404 25168
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 19248 24880 19300 24886
rect 19248 24822 19300 24828
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 16120 24744 16172 24750
rect 16120 24686 16172 24692
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16132 24410 16160 24686
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 14740 24132 14792 24138
rect 14740 24074 14792 24080
rect 14752 23866 14780 24074
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 14648 23180 14700 23186
rect 14648 23122 14700 23128
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14108 22642 14136 22714
rect 14096 22636 14148 22642
rect 14096 22578 14148 22584
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 14384 22234 14412 22510
rect 14568 22438 14596 22918
rect 15304 22778 15332 23054
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 14372 22228 14424 22234
rect 14372 22170 14424 22176
rect 15028 22098 15056 22374
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 15304 22030 15332 22714
rect 15396 22166 15424 23598
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15580 22234 15608 22986
rect 15856 22982 15884 24142
rect 16132 23866 16160 24346
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 16316 23662 16344 24686
rect 18524 24274 18552 24754
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 16408 23798 16436 24006
rect 17788 23866 17816 24074
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 16396 23792 16448 23798
rect 16396 23734 16448 23740
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15856 22710 15884 22918
rect 16868 22710 16896 22986
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 17052 22642 17080 22918
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15384 22160 15436 22166
rect 15384 22102 15436 22108
rect 15856 22098 15884 22374
rect 16868 22234 16896 22374
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 15844 22092 15896 22098
rect 17052 22094 17080 22578
rect 17144 22574 17172 23598
rect 17328 22778 17356 23598
rect 18708 23118 18736 23802
rect 19260 23798 19288 24822
rect 19892 24676 19944 24682
rect 19892 24618 19944 24624
rect 19904 24206 19932 24618
rect 20364 24614 20392 25162
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20352 24608 20404 24614
rect 20352 24550 20404 24556
rect 20364 24274 20392 24550
rect 20456 24342 20484 24754
rect 20444 24336 20496 24342
rect 20444 24278 20496 24284
rect 20824 24274 20852 25162
rect 21008 24818 21036 25638
rect 21836 25294 21864 26726
rect 22204 26382 22232 27338
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 22480 27130 22508 27270
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 22296 26450 22324 26726
rect 22664 26450 22692 27474
rect 23296 27396 23348 27402
rect 23296 27338 23348 27344
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 22848 26586 22876 26862
rect 23308 26790 23336 27338
rect 23860 27062 23888 28426
rect 24872 27690 24900 30058
rect 25056 29714 25084 30126
rect 25240 29782 25268 30602
rect 25228 29776 25280 29782
rect 25228 29718 25280 29724
rect 25792 29714 25820 31214
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25884 30802 25912 31078
rect 26344 30938 26372 31282
rect 26516 31272 26568 31278
rect 26516 31214 26568 31220
rect 27252 31272 27304 31278
rect 27252 31214 27304 31220
rect 26332 30932 26384 30938
rect 26332 30874 26384 30880
rect 25872 30796 25924 30802
rect 25872 30738 25924 30744
rect 26344 30394 26372 30874
rect 26528 30870 26556 31214
rect 27264 30938 27292 31214
rect 27252 30932 27304 30938
rect 27252 30874 27304 30880
rect 26516 30864 26568 30870
rect 26516 30806 26568 30812
rect 26332 30388 26384 30394
rect 26332 30330 26384 30336
rect 26528 30190 26556 30806
rect 26516 30184 26568 30190
rect 26516 30126 26568 30132
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 25780 29708 25832 29714
rect 25780 29650 25832 29656
rect 25056 28422 25084 29650
rect 25412 29640 25464 29646
rect 25412 29582 25464 29588
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 25148 29238 25176 29514
rect 25136 29232 25188 29238
rect 25136 29174 25188 29180
rect 25424 29170 25452 29582
rect 25412 29164 25464 29170
rect 25412 29106 25464 29112
rect 25884 28626 25912 29990
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26160 28626 26188 29106
rect 26528 28694 26556 30126
rect 26608 29572 26660 29578
rect 26608 29514 26660 29520
rect 26620 29306 26648 29514
rect 27540 29306 27568 31350
rect 27908 31142 27936 31622
rect 27896 31136 27948 31142
rect 27896 31078 27948 31084
rect 27908 30734 27936 31078
rect 28000 30802 28028 31826
rect 29196 31822 29224 32438
rect 29184 31816 29236 31822
rect 29012 31764 29184 31770
rect 29012 31758 29236 31764
rect 29012 31742 29224 31758
rect 29012 31482 29040 31742
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 29656 31278 29684 32982
rect 29748 32910 29776 34478
rect 29840 33522 29868 35634
rect 29828 33516 29880 33522
rect 29828 33458 29880 33464
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29932 32434 29960 36314
rect 30116 36242 30144 36518
rect 30484 36242 30512 37266
rect 30576 37194 30604 37266
rect 30564 37188 30616 37194
rect 30564 37130 30616 37136
rect 30576 36854 30604 37130
rect 30564 36848 30616 36854
rect 30564 36790 30616 36796
rect 30104 36236 30156 36242
rect 30024 36196 30104 36224
rect 30024 34950 30052 36196
rect 30104 36178 30156 36184
rect 30472 36236 30524 36242
rect 30472 36178 30524 36184
rect 30576 35766 30604 36790
rect 30564 35760 30616 35766
rect 30392 35720 30564 35748
rect 30012 34944 30064 34950
rect 30012 34886 30064 34892
rect 30104 34944 30156 34950
rect 30104 34886 30156 34892
rect 30116 34610 30144 34886
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 30012 34536 30064 34542
rect 30012 34478 30064 34484
rect 30024 34202 30052 34478
rect 30288 34400 30340 34406
rect 30288 34342 30340 34348
rect 30012 34196 30064 34202
rect 30012 34138 30064 34144
rect 30024 32978 30052 34138
rect 30102 33144 30158 33153
rect 30300 33114 30328 34342
rect 30392 33862 30420 35720
rect 30564 35702 30616 35708
rect 30472 35080 30524 35086
rect 30472 35022 30524 35028
rect 30484 34610 30512 35022
rect 30656 34944 30708 34950
rect 30656 34886 30708 34892
rect 30668 34746 30696 34886
rect 30656 34740 30708 34746
rect 30656 34682 30708 34688
rect 30472 34604 30524 34610
rect 30472 34546 30524 34552
rect 30564 34536 30616 34542
rect 30564 34478 30616 34484
rect 30472 34400 30524 34406
rect 30472 34342 30524 34348
rect 30380 33856 30432 33862
rect 30380 33798 30432 33804
rect 30380 33584 30432 33590
rect 30380 33526 30432 33532
rect 30102 33079 30104 33088
rect 30156 33079 30158 33088
rect 30288 33108 30340 33114
rect 30104 33050 30156 33056
rect 30288 33050 30340 33056
rect 30194 33008 30250 33017
rect 30012 32972 30064 32978
rect 30194 32943 30250 32952
rect 30012 32914 30064 32920
rect 30208 32910 30236 32943
rect 30196 32904 30248 32910
rect 30196 32846 30248 32852
rect 30392 32842 30420 33526
rect 30380 32836 30432 32842
rect 30380 32778 30432 32784
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 29828 32360 29880 32366
rect 30484 32314 30512 34342
rect 30576 32774 30604 34478
rect 30656 33856 30708 33862
rect 30656 33798 30708 33804
rect 30668 33590 30696 33798
rect 30656 33584 30708 33590
rect 30656 33526 30708 33532
rect 30564 32768 30616 32774
rect 30564 32710 30616 32716
rect 30576 32366 30604 32710
rect 29828 32302 29880 32308
rect 29840 31822 29868 32302
rect 30300 32286 30512 32314
rect 30564 32360 30616 32366
rect 30564 32302 30616 32308
rect 30300 32230 30328 32286
rect 29920 32224 29972 32230
rect 29920 32166 29972 32172
rect 30104 32224 30156 32230
rect 30104 32166 30156 32172
rect 30288 32224 30340 32230
rect 30288 32166 30340 32172
rect 30380 32224 30432 32230
rect 30380 32166 30432 32172
rect 29932 31958 29960 32166
rect 29920 31952 29972 31958
rect 29920 31894 29972 31900
rect 30116 31822 30144 32166
rect 30300 32026 30328 32166
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 30104 31816 30156 31822
rect 30104 31758 30156 31764
rect 30288 31680 30340 31686
rect 30288 31622 30340 31628
rect 30300 31414 30328 31622
rect 30288 31408 30340 31414
rect 30288 31350 30340 31356
rect 28908 31272 28960 31278
rect 28908 31214 28960 31220
rect 29644 31272 29696 31278
rect 29644 31214 29696 31220
rect 27988 30796 28040 30802
rect 27988 30738 28040 30744
rect 27896 30728 27948 30734
rect 27896 30670 27948 30676
rect 27620 30592 27672 30598
rect 27620 30534 27672 30540
rect 27632 29850 27660 30534
rect 27620 29844 27672 29850
rect 27620 29786 27672 29792
rect 28000 29578 28028 30738
rect 28920 30666 28948 31214
rect 30392 30938 30420 32166
rect 30472 31816 30524 31822
rect 30524 31764 30604 31770
rect 30472 31758 30604 31764
rect 30484 31742 30604 31758
rect 30668 31754 30696 33526
rect 30748 32768 30800 32774
rect 30748 32710 30800 32716
rect 30760 32434 30788 32710
rect 30748 32428 30800 32434
rect 30748 32370 30800 32376
rect 30576 31346 30604 31742
rect 30656 31748 30708 31754
rect 30656 31690 30708 31696
rect 30564 31340 30616 31346
rect 30564 31282 30616 31288
rect 30380 30932 30432 30938
rect 30380 30874 30432 30880
rect 30576 30802 30604 31282
rect 30564 30796 30616 30802
rect 30564 30738 30616 30744
rect 28908 30660 28960 30666
rect 28908 30602 28960 30608
rect 27988 29572 28040 29578
rect 27988 29514 28040 29520
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 26608 29300 26660 29306
rect 26608 29242 26660 29248
rect 27528 29300 27580 29306
rect 27528 29242 27580 29248
rect 27252 29096 27304 29102
rect 27252 29038 27304 29044
rect 27264 28762 27292 29038
rect 27252 28756 27304 28762
rect 27252 28698 27304 28704
rect 26516 28688 26568 28694
rect 26516 28630 26568 28636
rect 25872 28620 25924 28626
rect 25872 28562 25924 28568
rect 26148 28620 26200 28626
rect 26148 28562 26200 28568
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 24780 27662 24992 27690
rect 25148 27674 25176 28018
rect 25964 28008 26016 28014
rect 25964 27950 26016 27956
rect 25504 27940 25556 27946
rect 25504 27882 25556 27888
rect 25516 27674 25544 27882
rect 25872 27872 25924 27878
rect 25872 27814 25924 27820
rect 24780 27470 24808 27662
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 23848 27056 23900 27062
rect 23848 26998 23900 27004
rect 23296 26784 23348 26790
rect 23296 26726 23348 26732
rect 22836 26580 22888 26586
rect 22836 26522 22888 26528
rect 23308 26450 23336 26726
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 22652 26444 22704 26450
rect 22652 26386 22704 26392
rect 23296 26444 23348 26450
rect 23296 26386 23348 26392
rect 23860 26382 23888 26998
rect 24872 26926 24900 27474
rect 24964 27130 24992 27662
rect 25136 27668 25188 27674
rect 25136 27610 25188 27616
rect 25504 27668 25556 27674
rect 25504 27610 25556 27616
rect 25148 27554 25176 27610
rect 25148 27526 25268 27554
rect 25136 27396 25188 27402
rect 25136 27338 25188 27344
rect 24952 27124 25004 27130
rect 24952 27066 25004 27072
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 23848 26376 23900 26382
rect 23848 26318 23900 26324
rect 24952 26036 25004 26042
rect 24952 25978 25004 25984
rect 24964 25362 24992 25978
rect 25148 25770 25176 27338
rect 25240 26586 25268 27526
rect 25320 27328 25372 27334
rect 25320 27270 25372 27276
rect 25332 27062 25360 27270
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 25228 26580 25280 26586
rect 25228 26522 25280 26528
rect 25516 26450 25544 27610
rect 25688 27124 25740 27130
rect 25688 27066 25740 27072
rect 25700 26994 25728 27066
rect 25688 26988 25740 26994
rect 25688 26930 25740 26936
rect 25504 26444 25556 26450
rect 25504 26386 25556 26392
rect 25516 25838 25544 26386
rect 25700 26234 25728 26930
rect 25884 26450 25912 27814
rect 25976 27334 26004 27950
rect 26160 27538 26188 28562
rect 26148 27532 26200 27538
rect 26148 27474 26200 27480
rect 25964 27328 26016 27334
rect 25964 27270 26016 27276
rect 25872 26444 25924 26450
rect 25872 26386 25924 26392
rect 25700 26206 25820 26234
rect 25792 25974 25820 26206
rect 25780 25968 25832 25974
rect 25780 25910 25832 25916
rect 25504 25832 25556 25838
rect 25504 25774 25556 25780
rect 25136 25764 25188 25770
rect 25136 25706 25188 25712
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22112 24886 22140 25162
rect 22100 24880 22152 24886
rect 22100 24822 22152 24828
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 22296 24410 22324 25298
rect 22836 25288 22888 25294
rect 23388 25288 23440 25294
rect 22888 25236 22968 25242
rect 22836 25230 22968 25236
rect 23388 25230 23440 25236
rect 22848 25214 22968 25230
rect 22940 24954 22968 25214
rect 22928 24948 22980 24954
rect 22928 24890 22980 24896
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22572 24750 22600 24822
rect 22560 24744 22612 24750
rect 22560 24686 22612 24692
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 20352 24268 20404 24274
rect 20352 24210 20404 24216
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19996 23798 20024 24006
rect 20088 23866 20116 24142
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 20364 23730 20392 24210
rect 22572 24206 22600 24686
rect 22560 24200 22612 24206
rect 22560 24142 22612 24148
rect 22940 24070 22968 24890
rect 23400 24750 23428 25230
rect 25228 25220 25280 25226
rect 25228 25162 25280 25168
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23940 24744 23992 24750
rect 23940 24686 23992 24692
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 22928 24064 22980 24070
rect 22928 24006 22980 24012
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 18696 23112 18748 23118
rect 18696 23054 18748 23060
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 15844 22034 15896 22040
rect 16960 22066 17080 22094
rect 17224 22094 17276 22098
rect 17328 22094 17356 22714
rect 18064 22710 18092 22986
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 18156 22710 18184 22918
rect 19628 22778 19656 23598
rect 22940 23186 22968 24006
rect 23216 23730 23244 24550
rect 23400 23730 23428 24686
rect 23676 24274 23704 24686
rect 23664 24268 23716 24274
rect 23664 24210 23716 24216
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23492 23322 23520 23666
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23676 23186 23704 24210
rect 23952 23798 23980 24686
rect 25044 24676 25096 24682
rect 25044 24618 25096 24624
rect 25056 24274 25084 24618
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 24124 24132 24176 24138
rect 24124 24074 24176 24080
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 24136 23730 24164 24074
rect 25240 23866 25268 25162
rect 25516 24886 25544 25774
rect 25976 25770 26004 27270
rect 26160 27062 26188 27474
rect 26976 27464 27028 27470
rect 26976 27406 27028 27412
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 26160 26450 26188 26998
rect 26988 26926 27016 27406
rect 27540 27402 27568 29242
rect 27632 28966 27660 29446
rect 27620 28960 27672 28966
rect 27620 28902 27672 28908
rect 27632 28558 27660 28902
rect 28000 28626 28028 29514
rect 28920 29306 28948 30602
rect 30576 30326 30604 30738
rect 30564 30320 30616 30326
rect 30564 30262 30616 30268
rect 30852 30054 30880 39630
rect 30930 39552 30986 39630
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 31944 37936 31996 37942
rect 31944 37878 31996 37884
rect 32956 37936 33008 37942
rect 32956 37878 33008 37884
rect 31668 37868 31720 37874
rect 31668 37810 31720 37816
rect 31576 37664 31628 37670
rect 31576 37606 31628 37612
rect 31588 37194 31616 37606
rect 31576 37188 31628 37194
rect 31576 37130 31628 37136
rect 31484 37120 31536 37126
rect 31484 37062 31536 37068
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 31116 36780 31168 36786
rect 31116 36722 31168 36728
rect 31036 36378 31064 36722
rect 30932 36372 30984 36378
rect 30932 36314 30984 36320
rect 31024 36372 31076 36378
rect 31024 36314 31076 36320
rect 30944 36174 30972 36314
rect 31128 36242 31156 36722
rect 31300 36576 31352 36582
rect 31300 36518 31352 36524
rect 31116 36236 31168 36242
rect 31116 36178 31168 36184
rect 30932 36168 30984 36174
rect 30932 36110 30984 36116
rect 31312 35204 31340 36518
rect 31392 36100 31444 36106
rect 31392 36042 31444 36048
rect 31404 35766 31432 36042
rect 31392 35760 31444 35766
rect 31392 35702 31444 35708
rect 31392 35216 31444 35222
rect 31312 35176 31392 35204
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 30944 32910 30972 34546
rect 31312 33998 31340 35176
rect 31392 35158 31444 35164
rect 31496 34066 31524 37062
rect 31680 36718 31708 37810
rect 31852 37800 31904 37806
rect 31852 37742 31904 37748
rect 31864 37210 31892 37742
rect 31956 37466 31984 37878
rect 32864 37868 32916 37874
rect 32864 37810 32916 37816
rect 32220 37732 32272 37738
rect 32220 37674 32272 37680
rect 31944 37460 31996 37466
rect 31944 37402 31996 37408
rect 31956 37346 31984 37402
rect 31956 37318 32076 37346
rect 31864 37182 31984 37210
rect 31668 36712 31720 36718
rect 31668 36654 31720 36660
rect 31680 35894 31708 36654
rect 31852 36304 31904 36310
rect 31852 36246 31904 36252
rect 31864 36106 31892 36246
rect 31852 36100 31904 36106
rect 31852 36042 31904 36048
rect 31680 35866 31800 35894
rect 31772 35834 31800 35866
rect 31760 35828 31812 35834
rect 31760 35770 31812 35776
rect 31576 35692 31628 35698
rect 31576 35634 31628 35640
rect 31760 35692 31812 35698
rect 31760 35634 31812 35640
rect 31588 35494 31616 35634
rect 31576 35488 31628 35494
rect 31576 35430 31628 35436
rect 31588 35034 31616 35430
rect 31772 35154 31800 35634
rect 31864 35562 31892 36042
rect 31852 35556 31904 35562
rect 31852 35498 31904 35504
rect 31956 35154 31984 37182
rect 32048 36786 32076 37318
rect 32036 36780 32088 36786
rect 32036 36722 32088 36728
rect 32128 36712 32180 36718
rect 32128 36654 32180 36660
rect 32036 36372 32088 36378
rect 32036 36314 32088 36320
rect 32048 35562 32076 36314
rect 32140 36242 32168 36654
rect 32128 36236 32180 36242
rect 32128 36178 32180 36184
rect 32036 35556 32088 35562
rect 32036 35498 32088 35504
rect 32048 35154 32076 35498
rect 31760 35148 31812 35154
rect 31760 35090 31812 35096
rect 31944 35148 31996 35154
rect 31944 35090 31996 35096
rect 32036 35148 32088 35154
rect 32036 35090 32088 35096
rect 32140 35086 32168 36178
rect 32232 36038 32260 37674
rect 32312 37664 32364 37670
rect 32312 37606 32364 37612
rect 32496 37664 32548 37670
rect 32496 37606 32548 37612
rect 32324 36854 32352 37606
rect 32312 36848 32364 36854
rect 32312 36790 32364 36796
rect 32324 36242 32352 36790
rect 32404 36576 32456 36582
rect 32404 36518 32456 36524
rect 32312 36236 32364 36242
rect 32312 36178 32364 36184
rect 32416 36106 32444 36518
rect 32404 36100 32456 36106
rect 32404 36042 32456 36048
rect 32220 36032 32272 36038
rect 32220 35974 32272 35980
rect 32220 35692 32272 35698
rect 32220 35634 32272 35640
rect 31852 35080 31904 35086
rect 31588 35028 31852 35034
rect 31588 35022 31904 35028
rect 32128 35080 32180 35086
rect 32128 35022 32180 35028
rect 31588 35006 31892 35022
rect 32036 35012 32088 35018
rect 31680 34678 31708 35006
rect 32036 34954 32088 34960
rect 31852 34944 31904 34950
rect 31852 34886 31904 34892
rect 31864 34746 31892 34886
rect 31852 34740 31904 34746
rect 31852 34682 31904 34688
rect 31668 34672 31720 34678
rect 31668 34614 31720 34620
rect 31576 34604 31628 34610
rect 31576 34546 31628 34552
rect 31484 34060 31536 34066
rect 31484 34002 31536 34008
rect 31300 33992 31352 33998
rect 31300 33934 31352 33940
rect 30932 32904 30984 32910
rect 30932 32846 30984 32852
rect 31116 32904 31168 32910
rect 31116 32846 31168 32852
rect 31128 30938 31156 32846
rect 31312 32570 31340 33934
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31300 32564 31352 32570
rect 31300 32506 31352 32512
rect 31404 32502 31432 33458
rect 31588 33454 31616 34546
rect 31576 33448 31628 33454
rect 31576 33390 31628 33396
rect 31588 32978 31616 33390
rect 31864 33046 31892 34682
rect 31944 34604 31996 34610
rect 31944 34546 31996 34552
rect 31956 34202 31984 34546
rect 32048 34542 32076 34954
rect 32232 34746 32260 35634
rect 32312 35624 32364 35630
rect 32312 35566 32364 35572
rect 32220 34740 32272 34746
rect 32220 34682 32272 34688
rect 32324 34626 32352 35566
rect 32232 34610 32352 34626
rect 32508 34610 32536 37606
rect 32876 36582 32904 37810
rect 32968 36922 32996 37878
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 33968 37256 34020 37262
rect 33968 37198 34020 37204
rect 33232 37120 33284 37126
rect 33232 37062 33284 37068
rect 33416 37120 33468 37126
rect 33416 37062 33468 37068
rect 32956 36916 33008 36922
rect 32956 36858 33008 36864
rect 33244 36786 33272 37062
rect 33428 36854 33456 37062
rect 33980 36854 34008 37198
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 34796 36916 34848 36922
rect 34796 36858 34848 36864
rect 33416 36848 33468 36854
rect 33416 36790 33468 36796
rect 33968 36848 34020 36854
rect 34020 36808 34100 36836
rect 33968 36790 34020 36796
rect 33140 36780 33192 36786
rect 33140 36722 33192 36728
rect 33232 36780 33284 36786
rect 33232 36722 33284 36728
rect 32864 36576 32916 36582
rect 32864 36518 32916 36524
rect 32876 36038 32904 36518
rect 33152 36174 33180 36722
rect 33140 36168 33192 36174
rect 33140 36110 33192 36116
rect 32772 36032 32824 36038
rect 32772 35974 32824 35980
rect 32864 36032 32916 36038
rect 32864 35974 32916 35980
rect 32784 35737 32812 35974
rect 33152 35834 33180 36110
rect 33140 35828 33192 35834
rect 33140 35770 33192 35776
rect 33244 35766 33272 36722
rect 33508 36712 33560 36718
rect 33508 36654 33560 36660
rect 33324 36576 33376 36582
rect 33324 36518 33376 36524
rect 33336 36174 33364 36518
rect 33520 36378 33548 36654
rect 33508 36372 33560 36378
rect 33508 36314 33560 36320
rect 33324 36168 33376 36174
rect 33600 36168 33652 36174
rect 33376 36128 33600 36156
rect 33324 36110 33376 36116
rect 33232 35760 33284 35766
rect 32770 35728 32826 35737
rect 33232 35702 33284 35708
rect 32770 35663 32826 35672
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 32770 35592 32826 35601
rect 32770 35527 32772 35536
rect 32824 35527 32826 35536
rect 32772 35498 32824 35504
rect 33048 35488 33100 35494
rect 33048 35430 33100 35436
rect 32678 35184 32734 35193
rect 32678 35119 32680 35128
rect 32732 35119 32734 35128
rect 32680 35090 32732 35096
rect 33060 35018 33088 35430
rect 33336 35222 33364 35634
rect 33324 35216 33376 35222
rect 33324 35158 33376 35164
rect 33232 35080 33284 35086
rect 33324 35080 33376 35086
rect 33232 35022 33284 35028
rect 33322 35048 33324 35057
rect 33376 35048 33378 35057
rect 33048 35012 33100 35018
rect 33048 34954 33100 34960
rect 33060 34678 33088 34954
rect 33244 34746 33272 35022
rect 33322 34983 33378 34992
rect 33232 34740 33284 34746
rect 33232 34682 33284 34688
rect 33048 34672 33100 34678
rect 33048 34614 33100 34620
rect 33244 34610 33272 34682
rect 32220 34604 32352 34610
rect 32272 34598 32352 34604
rect 32496 34604 32548 34610
rect 32220 34546 32272 34552
rect 32496 34546 32548 34552
rect 33232 34604 33284 34610
rect 33232 34546 33284 34552
rect 32036 34536 32088 34542
rect 32036 34478 32088 34484
rect 33244 34474 33272 34546
rect 33232 34468 33284 34474
rect 33232 34410 33284 34416
rect 33048 34400 33100 34406
rect 33048 34342 33100 34348
rect 31944 34196 31996 34202
rect 31944 34138 31996 34144
rect 32772 34060 32824 34066
rect 32772 34002 32824 34008
rect 32784 33590 32812 34002
rect 33060 33658 33088 34342
rect 33048 33652 33100 33658
rect 33048 33594 33100 33600
rect 32772 33584 32824 33590
rect 32772 33526 32824 33532
rect 32404 33312 32456 33318
rect 32404 33254 32456 33260
rect 31852 33040 31904 33046
rect 31852 32982 31904 32988
rect 31576 32972 31628 32978
rect 31576 32914 31628 32920
rect 32416 32910 32444 33254
rect 33336 32978 33364 34983
rect 33428 34746 33456 36128
rect 33652 36128 33916 36156
rect 33600 36110 33652 36116
rect 33600 35692 33652 35698
rect 33600 35634 33652 35640
rect 33612 35290 33640 35634
rect 33600 35284 33652 35290
rect 33600 35226 33652 35232
rect 33888 35154 33916 36128
rect 34072 35766 34100 36808
rect 34808 36310 34836 36858
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34796 36304 34848 36310
rect 34796 36246 34848 36252
rect 34796 36168 34848 36174
rect 34796 36110 34848 36116
rect 34612 36032 34664 36038
rect 34612 35974 34664 35980
rect 34244 35828 34296 35834
rect 34244 35770 34296 35776
rect 33968 35760 34020 35766
rect 33968 35702 34020 35708
rect 34060 35760 34112 35766
rect 34060 35702 34112 35708
rect 33508 35148 33560 35154
rect 33508 35090 33560 35096
rect 33876 35148 33928 35154
rect 33876 35090 33928 35096
rect 33416 34740 33468 34746
rect 33416 34682 33468 34688
rect 33416 34604 33468 34610
rect 33416 34546 33468 34552
rect 33428 34202 33456 34546
rect 33416 34196 33468 34202
rect 33416 34138 33468 34144
rect 33520 33522 33548 35090
rect 33600 35080 33652 35086
rect 33600 35022 33652 35028
rect 33612 34950 33640 35022
rect 33600 34944 33652 34950
rect 33600 34886 33652 34892
rect 33508 33516 33560 33522
rect 33508 33458 33560 33464
rect 33612 33454 33640 34886
rect 33980 34610 34008 35702
rect 34152 35488 34204 35494
rect 34152 35430 34204 35436
rect 33692 34604 33744 34610
rect 33692 34546 33744 34552
rect 33968 34604 34020 34610
rect 33968 34546 34020 34552
rect 33704 33658 33732 34546
rect 34060 34400 34112 34406
rect 34060 34342 34112 34348
rect 33692 33652 33744 33658
rect 33692 33594 33744 33600
rect 34072 33454 34100 34342
rect 34164 33454 34192 35430
rect 34256 34218 34284 35770
rect 34428 35760 34480 35766
rect 34428 35702 34480 35708
rect 34440 34660 34468 35702
rect 34624 35193 34652 35974
rect 34610 35184 34666 35193
rect 34610 35119 34666 35128
rect 34624 34898 34652 35119
rect 34808 35086 34836 36110
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 35624 35488 35676 35494
rect 35624 35430 35676 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35636 35086 35664 35430
rect 34796 35080 34848 35086
rect 35532 35080 35584 35086
rect 34796 35022 34848 35028
rect 35530 35048 35532 35057
rect 35624 35080 35676 35086
rect 35584 35048 35586 35057
rect 35624 35022 35676 35028
rect 35530 34983 35586 34992
rect 34624 34870 34744 34898
rect 34612 34740 34664 34746
rect 34612 34682 34664 34688
rect 34520 34672 34572 34678
rect 34440 34632 34520 34660
rect 34520 34614 34572 34620
rect 34336 34536 34388 34542
rect 34336 34478 34388 34484
rect 34348 34406 34376 34478
rect 34336 34400 34388 34406
rect 34336 34342 34388 34348
rect 34256 34190 34376 34218
rect 34348 33998 34376 34190
rect 34336 33992 34388 33998
rect 34336 33934 34388 33940
rect 33600 33448 33652 33454
rect 33600 33390 33652 33396
rect 34060 33448 34112 33454
rect 34060 33390 34112 33396
rect 34152 33448 34204 33454
rect 34152 33390 34204 33396
rect 33600 33040 33652 33046
rect 33600 32982 33652 32988
rect 33324 32972 33376 32978
rect 33324 32914 33376 32920
rect 32404 32904 32456 32910
rect 32404 32846 32456 32852
rect 31668 32836 31720 32842
rect 31668 32778 31720 32784
rect 33232 32836 33284 32842
rect 33232 32778 33284 32784
rect 31392 32496 31444 32502
rect 31392 32438 31444 32444
rect 31404 31890 31432 32438
rect 31680 32434 31708 32778
rect 32864 32564 32916 32570
rect 32864 32506 32916 32512
rect 32876 32450 32904 32506
rect 31668 32428 31720 32434
rect 31668 32370 31720 32376
rect 32588 32428 32640 32434
rect 32876 32422 33180 32450
rect 32588 32370 32640 32376
rect 31392 31884 31444 31890
rect 31392 31826 31444 31832
rect 31680 31346 31708 32370
rect 32312 32292 32364 32298
rect 32312 32234 32364 32240
rect 32324 31346 32352 32234
rect 32600 32026 32628 32370
rect 32588 32020 32640 32026
rect 32588 31962 32640 31968
rect 32864 31748 32916 31754
rect 32864 31690 32916 31696
rect 32876 31482 32904 31690
rect 32864 31476 32916 31482
rect 32864 31418 32916 31424
rect 31668 31340 31720 31346
rect 31668 31282 31720 31288
rect 32312 31340 32364 31346
rect 32312 31282 32364 31288
rect 33152 31278 33180 32422
rect 32588 31272 32640 31278
rect 32588 31214 32640 31220
rect 33140 31272 33192 31278
rect 33140 31214 33192 31220
rect 31116 30932 31168 30938
rect 31116 30874 31168 30880
rect 32404 30796 32456 30802
rect 32404 30738 32456 30744
rect 31116 30660 31168 30666
rect 31116 30602 31168 30608
rect 31576 30660 31628 30666
rect 31576 30602 31628 30608
rect 31944 30660 31996 30666
rect 31944 30602 31996 30608
rect 30840 30048 30892 30054
rect 30840 29990 30892 29996
rect 29092 29708 29144 29714
rect 29092 29650 29144 29656
rect 28908 29300 28960 29306
rect 28908 29242 28960 29248
rect 27988 28620 28040 28626
rect 27988 28562 28040 28568
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 28920 28150 28948 29242
rect 29000 28960 29052 28966
rect 29000 28902 29052 28908
rect 29012 28558 29040 28902
rect 29104 28694 29132 29650
rect 29552 29504 29604 29510
rect 29552 29446 29604 29452
rect 29920 29504 29972 29510
rect 29920 29446 29972 29452
rect 30104 29504 30156 29510
rect 30104 29446 30156 29452
rect 29092 28688 29144 28694
rect 29092 28630 29144 28636
rect 29276 28620 29328 28626
rect 29276 28562 29328 28568
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 29288 28218 29316 28562
rect 29276 28212 29328 28218
rect 29276 28154 29328 28160
rect 29564 28150 29592 29446
rect 29932 28626 29960 29446
rect 30116 29306 30144 29446
rect 30104 29300 30156 29306
rect 30104 29242 30156 29248
rect 30116 28694 30144 29242
rect 30472 29096 30524 29102
rect 30472 29038 30524 29044
rect 30840 29096 30892 29102
rect 30840 29038 30892 29044
rect 30484 28762 30512 29038
rect 30472 28756 30524 28762
rect 30472 28698 30524 28704
rect 30104 28688 30156 28694
rect 30104 28630 30156 28636
rect 30852 28626 30880 29038
rect 31128 28994 31156 30602
rect 31484 30592 31536 30598
rect 31484 30534 31536 30540
rect 31496 30190 31524 30534
rect 31588 30258 31616 30602
rect 31576 30252 31628 30258
rect 31576 30194 31628 30200
rect 31484 30184 31536 30190
rect 31484 30126 31536 30132
rect 31956 30054 31984 30602
rect 32416 30394 32444 30738
rect 32600 30734 32628 31214
rect 33244 30954 33272 32778
rect 33612 31686 33640 32982
rect 34348 32978 34376 33934
rect 34532 33930 34560 34614
rect 34624 34066 34652 34682
rect 34612 34060 34664 34066
rect 34612 34002 34664 34008
rect 34520 33924 34572 33930
rect 34520 33866 34572 33872
rect 34428 33856 34480 33862
rect 34428 33798 34480 33804
rect 34612 33856 34664 33862
rect 34612 33798 34664 33804
rect 34440 33658 34468 33798
rect 34428 33652 34480 33658
rect 34428 33594 34480 33600
rect 34624 33538 34652 33798
rect 34716 33658 34744 34870
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35716 33992 35768 33998
rect 35360 33940 35716 33946
rect 35360 33934 35768 33940
rect 35256 33924 35308 33930
rect 35256 33866 35308 33872
rect 35360 33918 35756 33934
rect 34704 33652 34756 33658
rect 34704 33594 34756 33600
rect 34440 33510 34652 33538
rect 34704 33516 34756 33522
rect 34440 33017 34468 33510
rect 34704 33458 34756 33464
rect 34520 33380 34572 33386
rect 34520 33322 34572 33328
rect 34426 33008 34482 33017
rect 34336 32972 34388 32978
rect 34426 32943 34482 32952
rect 34336 32914 34388 32920
rect 33968 32496 34020 32502
rect 33968 32438 34020 32444
rect 33980 31822 34008 32438
rect 34428 32428 34480 32434
rect 34532 32416 34560 33322
rect 34612 33312 34664 33318
rect 34612 33254 34664 33260
rect 34624 33153 34652 33254
rect 34610 33144 34666 33153
rect 34716 33114 34744 33458
rect 35268 33454 35296 33866
rect 34796 33448 34848 33454
rect 34796 33390 34848 33396
rect 35256 33448 35308 33454
rect 35256 33390 35308 33396
rect 34610 33079 34666 33088
rect 34704 33108 34756 33114
rect 34704 33050 34756 33056
rect 34480 32388 34560 32416
rect 34428 32370 34480 32376
rect 34612 32360 34664 32366
rect 34612 32302 34664 32308
rect 34520 32292 34572 32298
rect 34520 32234 34572 32240
rect 34152 32224 34204 32230
rect 34152 32166 34204 32172
rect 34164 31890 34192 32166
rect 34152 31884 34204 31890
rect 34152 31826 34204 31832
rect 33968 31816 34020 31822
rect 33968 31758 34020 31764
rect 33600 31680 33652 31686
rect 33600 31622 33652 31628
rect 33060 30926 33272 30954
rect 33060 30870 33088 30926
rect 33048 30864 33100 30870
rect 33048 30806 33100 30812
rect 32588 30728 32640 30734
rect 32588 30670 32640 30676
rect 32404 30388 32456 30394
rect 32404 30330 32456 30336
rect 31944 30048 31996 30054
rect 31944 29990 31996 29996
rect 31760 29640 31812 29646
rect 31760 29582 31812 29588
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 30944 28966 31156 28994
rect 29920 28620 29972 28626
rect 29920 28562 29972 28568
rect 30840 28620 30892 28626
rect 30840 28562 30892 28568
rect 30944 28490 30972 28966
rect 30932 28484 30984 28490
rect 30932 28426 30984 28432
rect 30944 28234 30972 28426
rect 30852 28206 30972 28234
rect 28908 28144 28960 28150
rect 28908 28086 28960 28092
rect 29552 28144 29604 28150
rect 29552 28086 29604 28092
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 27436 27056 27488 27062
rect 27540 27044 27568 27338
rect 27712 27328 27764 27334
rect 27712 27270 27764 27276
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 29184 27328 29236 27334
rect 29184 27270 29236 27276
rect 27488 27016 27568 27044
rect 27436 26998 27488 27004
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 26976 26920 27028 26926
rect 26976 26862 27028 26868
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 26160 26042 26188 26386
rect 26148 26036 26200 26042
rect 26148 25978 26200 25984
rect 26528 25974 26556 26862
rect 27448 26314 27476 26998
rect 27724 26586 27752 27270
rect 28184 27062 28212 27270
rect 28172 27056 28224 27062
rect 28172 26998 28224 27004
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 28460 26450 28488 27270
rect 29196 26926 29224 27270
rect 30024 26926 30052 28018
rect 30104 28008 30156 28014
rect 30104 27950 30156 27956
rect 29000 26920 29052 26926
rect 29000 26862 29052 26868
rect 29184 26920 29236 26926
rect 29184 26862 29236 26868
rect 30012 26920 30064 26926
rect 30012 26862 30064 26868
rect 29012 26450 29040 26862
rect 30116 26790 30144 27950
rect 30472 27940 30524 27946
rect 30472 27882 30524 27888
rect 30484 27538 30512 27882
rect 30656 27872 30708 27878
rect 30656 27814 30708 27820
rect 30472 27532 30524 27538
rect 30472 27474 30524 27480
rect 30564 27396 30616 27402
rect 30564 27338 30616 27344
rect 30576 27062 30604 27338
rect 30668 27062 30696 27814
rect 30852 27418 30880 28206
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 30760 27402 30880 27418
rect 30748 27396 30880 27402
rect 30800 27390 30880 27396
rect 30748 27338 30800 27344
rect 30944 27130 30972 28018
rect 31024 28008 31076 28014
rect 31024 27950 31076 27956
rect 31300 28008 31352 28014
rect 31300 27950 31352 27956
rect 31036 27334 31064 27950
rect 31312 27470 31340 27950
rect 31300 27464 31352 27470
rect 31300 27406 31352 27412
rect 31024 27328 31076 27334
rect 31024 27270 31076 27276
rect 31036 27130 31064 27270
rect 30932 27124 30984 27130
rect 30932 27066 30984 27072
rect 31024 27124 31076 27130
rect 31024 27066 31076 27072
rect 30380 27056 30432 27062
rect 30380 26998 30432 27004
rect 30564 27056 30616 27062
rect 30564 26998 30616 27004
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30104 26784 30156 26790
rect 30104 26726 30156 26732
rect 30116 26450 30144 26726
rect 28448 26444 28500 26450
rect 28448 26386 28500 26392
rect 29000 26444 29052 26450
rect 29000 26386 29052 26392
rect 30104 26444 30156 26450
rect 30104 26386 30156 26392
rect 26700 26308 26752 26314
rect 26700 26250 26752 26256
rect 27436 26308 27488 26314
rect 27436 26250 27488 26256
rect 30012 26308 30064 26314
rect 30012 26250 30064 26256
rect 26516 25968 26568 25974
rect 26516 25910 26568 25916
rect 26712 25838 26740 26250
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 26700 25832 26752 25838
rect 26700 25774 26752 25780
rect 25964 25764 26016 25770
rect 25964 25706 26016 25712
rect 25504 24880 25556 24886
rect 25504 24822 25556 24828
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25884 24410 25912 24754
rect 26252 24750 26280 25774
rect 27448 25294 27476 26250
rect 30024 25974 30052 26250
rect 30392 26246 30420 26998
rect 30944 26432 30972 27066
rect 31312 26994 31340 27406
rect 31404 26994 31432 29106
rect 31772 27946 31800 29582
rect 31956 29170 31984 29990
rect 33060 29714 33088 30806
rect 33612 30734 33640 31622
rect 33600 30728 33652 30734
rect 33600 30670 33652 30676
rect 33980 30394 34008 31758
rect 33508 30388 33560 30394
rect 33508 30330 33560 30336
rect 33968 30388 34020 30394
rect 33968 30330 34020 30336
rect 33048 29708 33100 29714
rect 33048 29650 33100 29656
rect 32496 29504 32548 29510
rect 32496 29446 32548 29452
rect 33416 29504 33468 29510
rect 33416 29446 33468 29452
rect 32508 29238 32536 29446
rect 32496 29232 32548 29238
rect 32496 29174 32548 29180
rect 31944 29164 31996 29170
rect 31944 29106 31996 29112
rect 33140 29096 33192 29102
rect 33140 29038 33192 29044
rect 31852 29028 31904 29034
rect 31852 28970 31904 28976
rect 31864 28558 31892 28970
rect 31852 28552 31904 28558
rect 31852 28494 31904 28500
rect 31864 28014 31892 28494
rect 32680 28484 32732 28490
rect 32680 28426 32732 28432
rect 32692 28150 32720 28426
rect 33152 28150 33180 29038
rect 33428 28626 33456 29446
rect 33520 29238 33548 30330
rect 34164 30258 34192 31826
rect 34532 31346 34560 32234
rect 34624 31958 34652 32302
rect 34612 31952 34664 31958
rect 34612 31894 34664 31900
rect 34624 31346 34652 31894
rect 34808 31414 34836 33390
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35256 32972 35308 32978
rect 35256 32914 35308 32920
rect 35164 32836 35216 32842
rect 35164 32778 35216 32784
rect 35176 32434 35204 32778
rect 35268 32434 35296 32914
rect 35360 32774 35388 33918
rect 35440 33856 35492 33862
rect 35440 33798 35492 33804
rect 35452 32910 35480 33798
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 35440 32904 35492 32910
rect 35440 32846 35492 32852
rect 35348 32768 35400 32774
rect 35348 32710 35400 32716
rect 35164 32428 35216 32434
rect 35164 32370 35216 32376
rect 35256 32428 35308 32434
rect 35256 32370 35308 32376
rect 35360 32230 35388 32710
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 35348 32224 35400 32230
rect 35348 32166 35400 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35440 31884 35492 31890
rect 35440 31826 35492 31832
rect 34796 31408 34848 31414
rect 34796 31350 34848 31356
rect 34520 31340 34572 31346
rect 34520 31282 34572 31288
rect 34612 31340 34664 31346
rect 34612 31282 34664 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34612 30728 34664 30734
rect 34612 30670 34664 30676
rect 35348 30728 35400 30734
rect 35348 30670 35400 30676
rect 34520 30660 34572 30666
rect 34520 30602 34572 30608
rect 34532 30326 34560 30602
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 33876 29708 33928 29714
rect 33876 29650 33928 29656
rect 33508 29232 33560 29238
rect 33508 29174 33560 29180
rect 33416 28620 33468 28626
rect 33416 28562 33468 28568
rect 33428 28218 33456 28562
rect 33784 28484 33836 28490
rect 33784 28426 33836 28432
rect 33416 28212 33468 28218
rect 33416 28154 33468 28160
rect 32680 28144 32732 28150
rect 32680 28086 32732 28092
rect 33140 28144 33192 28150
rect 33140 28086 33192 28092
rect 31852 28008 31904 28014
rect 31852 27950 31904 27956
rect 31760 27940 31812 27946
rect 31760 27882 31812 27888
rect 32128 27668 32180 27674
rect 32128 27610 32180 27616
rect 32140 27062 32168 27610
rect 33152 27402 33180 28086
rect 33232 27668 33284 27674
rect 33232 27610 33284 27616
rect 33140 27396 33192 27402
rect 33140 27338 33192 27344
rect 32128 27056 32180 27062
rect 32128 26998 32180 27004
rect 31300 26988 31352 26994
rect 31300 26930 31352 26936
rect 31392 26988 31444 26994
rect 31392 26930 31444 26936
rect 31024 26444 31076 26450
rect 30944 26404 31024 26432
rect 31024 26386 31076 26392
rect 30380 26240 30432 26246
rect 30380 26182 30432 26188
rect 30392 25974 30420 26182
rect 30012 25968 30064 25974
rect 30012 25910 30064 25916
rect 30380 25968 30432 25974
rect 30380 25910 30432 25916
rect 28080 25900 28132 25906
rect 28080 25842 28132 25848
rect 28264 25900 28316 25906
rect 28264 25842 28316 25848
rect 29644 25900 29696 25906
rect 29644 25842 29696 25848
rect 27804 25832 27856 25838
rect 27804 25774 27856 25780
rect 27436 25288 27488 25294
rect 27488 25236 27568 25242
rect 27436 25230 27568 25236
rect 26608 25220 26660 25226
rect 27448 25214 27568 25230
rect 26608 25162 26660 25168
rect 26056 24744 26108 24750
rect 26056 24686 26108 24692
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 25872 24404 25924 24410
rect 25872 24346 25924 24352
rect 25884 23866 25912 24346
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 26068 23662 26096 24686
rect 26252 24206 26280 24686
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 23756 23656 23808 23662
rect 23756 23598 23808 23604
rect 26056 23656 26108 23662
rect 26056 23598 26108 23604
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 18052 22704 18104 22710
rect 18052 22646 18104 22652
rect 18144 22704 18196 22710
rect 18144 22646 18196 22652
rect 17224 22092 17356 22094
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 16960 21962 16988 22066
rect 17276 22066 17356 22092
rect 17224 22034 17276 22040
rect 18156 21962 18184 22646
rect 19628 22642 19656 22714
rect 19996 22710 20024 22986
rect 19984 22704 20036 22710
rect 19984 22646 20036 22652
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 20548 22574 20576 23054
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20640 22098 20668 22714
rect 21192 22234 21220 22986
rect 21376 22506 21404 23122
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22204 22710 22232 22918
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 22480 22234 22508 23054
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 23584 22778 23612 22986
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 22652 22704 22704 22710
rect 22652 22646 22704 22652
rect 22560 22568 22612 22574
rect 22664 22556 22692 22646
rect 22612 22528 22692 22556
rect 22560 22510 22612 22516
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 20628 22092 20680 22098
rect 20628 22034 20680 22040
rect 22572 21962 22600 22510
rect 23584 22030 23612 22714
rect 23676 22642 23704 23122
rect 23664 22636 23716 22642
rect 23664 22578 23716 22584
rect 23676 22098 23704 22578
rect 23664 22092 23716 22098
rect 23664 22034 23716 22040
rect 23768 22030 23796 23598
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23952 22778 23980 22918
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 24044 22030 24072 22510
rect 25044 22500 25096 22506
rect 25044 22442 25096 22448
rect 25056 22234 25084 22442
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 25424 22098 25452 22578
rect 25504 22432 25556 22438
rect 25504 22374 25556 22380
rect 25412 22092 25464 22098
rect 25412 22034 25464 22040
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 22560 21956 22612 21962
rect 22560 21898 22612 21904
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10796 21146 10824 21422
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10060 20874 10088 20946
rect 11072 20874 11100 21898
rect 16856 20936 16908 20942
rect 18156 20890 18184 21898
rect 16856 20878 16908 20884
rect 10048 20868 10100 20874
rect 10048 20810 10100 20816
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 16028 20868 16080 20874
rect 16028 20810 16080 20816
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 9876 20590 9996 20618
rect 10060 20602 10088 20810
rect 10048 20596 10100 20602
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9876 19854 9904 20590
rect 10048 20538 10100 20544
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 10060 19378 10088 20538
rect 11072 20534 11100 20810
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 15936 20528 15988 20534
rect 16040 20516 16068 20810
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16132 20602 16160 20742
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 15988 20488 16068 20516
rect 15936 20470 15988 20476
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 11072 20058 11100 20334
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 13832 19378 13860 20334
rect 15580 20262 15608 20402
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 7944 18358 7972 18566
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6564 17338 6592 17546
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6932 17270 6960 17682
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 5632 17264 5684 17270
rect 5552 17224 5632 17252
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 5552 16522 5580 17224
rect 5632 17206 5684 17212
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5552 15434 5580 16458
rect 6932 15502 6960 17206
rect 7484 17202 7512 17478
rect 7944 17270 7972 18294
rect 9416 18086 9444 18634
rect 10060 18426 10088 19314
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9416 17270 9444 18022
rect 9876 17882 9904 18158
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8036 16794 8064 17070
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8588 16590 8616 16934
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 9416 16522 9444 17206
rect 9876 17202 9904 17614
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9508 16726 9536 16934
rect 9600 16794 9628 16934
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9876 16590 9904 17138
rect 10060 16658 10088 18362
rect 13832 18290 13860 19314
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 15028 18834 15056 19246
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 15580 18766 15608 20198
rect 16040 19446 16068 20488
rect 16132 19514 16160 20538
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18834 15884 19110
rect 16316 18902 16344 20334
rect 16592 19446 16620 20810
rect 16868 19786 16896 20878
rect 17972 20874 18184 20890
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 17972 20868 18196 20874
rect 17972 20862 18144 20868
rect 17144 20534 17172 20810
rect 17972 20806 18000 20862
rect 18144 20810 18196 20816
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 18064 20398 18092 20742
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14936 18358 14964 18566
rect 14924 18352 14976 18358
rect 14924 18294 14976 18300
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11348 17882 11376 18022
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 11348 17678 11376 17818
rect 14292 17746 14320 18226
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 10520 17134 10548 17614
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 11072 17202 11100 17478
rect 14292 17202 14320 17682
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14568 17270 14596 17546
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 15672 17202 15700 18294
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15570 7236 15846
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5276 14482 5304 14758
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 4632 14362 4660 14418
rect 3332 14340 3384 14346
rect 4632 14334 4752 14362
rect 5552 14346 5580 15370
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5736 14890 5764 15030
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 3332 14282 3384 14288
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 3068 13394 3096 13942
rect 3160 13530 3188 14214
rect 4448 14006 4476 14214
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4724 13938 4752 14334
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5552 14074 5580 14282
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 5644 13870 5672 14758
rect 6748 14618 6776 14826
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6932 14346 6960 15438
rect 7300 15366 7328 16458
rect 10520 16182 10548 17070
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16658 10916 16934
rect 11072 16794 11100 17138
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 14108 16658 14136 17138
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 10508 16176 10560 16182
rect 10508 16118 10560 16124
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7668 15570 7696 15982
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 15162 7328 15302
rect 7668 15162 7696 15506
rect 7760 15162 7788 15914
rect 10520 15706 10548 16118
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10612 15570 10640 16594
rect 15672 16522 15700 17138
rect 16040 16998 16068 17614
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 15570 10916 15846
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7944 14958 7972 15030
rect 8036 14958 8064 15302
rect 8496 15026 8524 15302
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6932 14006 6960 14282
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 7944 13870 7972 14894
rect 8864 14006 8892 14894
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 9232 13938 9260 15302
rect 9692 14482 9720 15302
rect 10060 14958 10088 15370
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10152 15094 10180 15302
rect 10336 15162 10364 15438
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10612 15026 10640 15302
rect 11072 15162 11100 15914
rect 11348 15434 11376 16458
rect 15672 16182 15700 16458
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 14292 15434 14320 16050
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14384 15570 14412 15982
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 14482 9904 14758
rect 10796 14618 10824 14894
rect 11348 14890 11376 15370
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 11348 14482 11376 14826
rect 14292 14482 14320 15370
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 9692 13938 9720 14418
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 14292 13870 14320 14418
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 14292 12850 14320 13806
rect 14568 13394 14596 13806
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 10336 800 10364 12242
rect 15212 12238 15240 12718
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 10674 13768 11630
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13740 10418 13768 10610
rect 13648 10390 13768 10418
rect 13648 9586 13676 10390
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13924 9654 13952 9930
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14108 8566 14136 8842
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14292 8294 14320 8978
rect 15304 8974 15332 16050
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15488 15706 15516 15982
rect 15672 15858 15700 16118
rect 15856 16114 15884 16390
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15580 15830 15700 15858
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15580 15570 15608 15830
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15568 15564 15620 15570
rect 15488 15524 15568 15552
rect 15488 14346 15516 15524
rect 15568 15506 15620 15512
rect 15672 15026 15700 15642
rect 15856 15502 15884 16050
rect 15948 15706 15976 16594
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16224 15434 16252 18634
rect 16316 17116 16344 18838
rect 16868 18766 16896 19722
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17788 19378 17816 19654
rect 18064 19446 18092 20334
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17776 19372 17828 19378
rect 18156 19334 18184 20810
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 19248 20528 19300 20534
rect 19248 20470 19300 20476
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18432 20058 18460 20402
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18432 19514 18460 19994
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 17776 19314 17828 19320
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16500 18426 16528 18566
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16500 17610 16528 18362
rect 16868 17746 16896 18702
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16868 17134 16896 17682
rect 16856 17128 16908 17134
rect 16316 17088 16528 17116
rect 16500 16998 16528 17088
rect 16856 17070 16908 17076
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16408 15570 16436 16934
rect 16500 15570 16528 16934
rect 16868 15570 16896 17070
rect 17144 16250 17172 19314
rect 17972 19306 18184 19334
rect 17972 18698 18000 19306
rect 18340 18970 18368 19382
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17236 18426 17264 18634
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 17972 17592 18000 18634
rect 18340 18358 18368 18906
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18616 18222 18644 19246
rect 19064 18352 19116 18358
rect 19064 18294 19116 18300
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18052 17604 18104 17610
rect 17972 17564 18052 17592
rect 17880 17338 17908 17546
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17592 17264 17644 17270
rect 17972 17218 18000 17564
rect 18052 17546 18104 17552
rect 18616 17542 18644 18158
rect 19076 17882 19104 18294
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 19076 17338 19104 17818
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 17644 17212 18000 17218
rect 17592 17206 18000 17212
rect 17604 17190 18000 17206
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 17788 16590 17816 17070
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15580 14346 15608 14894
rect 15764 14618 15792 14894
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15488 14090 15516 14282
rect 15488 14062 15608 14090
rect 15580 14006 15608 14062
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15764 13326 15792 14554
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15580 12730 15608 13262
rect 15660 12776 15712 12782
rect 15580 12724 15660 12730
rect 15580 12718 15712 12724
rect 15580 12702 15700 12718
rect 15580 12238 15608 12702
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15856 12238 15884 12582
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15396 10062 15424 10746
rect 15948 10130 15976 15370
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13394 16068 13670
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16040 12170 16068 13330
rect 16408 13190 16436 14214
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12918 16436 13126
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 16224 11898 16252 12174
rect 16408 12170 16436 12854
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16040 10810 16068 11834
rect 16408 11830 16436 12106
rect 16396 11824 16448 11830
rect 16396 11766 16448 11772
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16224 11354 16252 11630
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 16132 10062 16160 11154
rect 16224 10606 16252 11290
rect 16408 11082 16436 11766
rect 16500 11694 16528 15506
rect 17328 15434 17356 16458
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 16684 14482 16712 14894
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 17604 14074 17632 14894
rect 17972 14822 18000 15370
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 14074 18000 14758
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18064 14074 18092 14214
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18248 13802 18276 17002
rect 18524 16590 18552 17070
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18432 15910 18460 16526
rect 18984 16114 19012 16594
rect 19168 16574 19196 20266
rect 19260 19786 19288 20470
rect 20732 20398 20760 20742
rect 20824 20398 20852 20742
rect 22112 20534 22140 20810
rect 22572 20534 22600 21898
rect 25516 21894 25544 22374
rect 25976 22234 26004 22578
rect 26068 22556 26096 23598
rect 26252 23186 26280 24142
rect 26516 24132 26568 24138
rect 26516 24074 26568 24080
rect 26528 23866 26556 24074
rect 26516 23860 26568 23866
rect 26516 23802 26568 23808
rect 26620 23746 26648 25162
rect 27436 25152 27488 25158
rect 27436 25094 27488 25100
rect 27448 23798 27476 25094
rect 27540 24886 27568 25214
rect 27528 24880 27580 24886
rect 27528 24822 27580 24828
rect 27540 24206 27568 24822
rect 27816 24750 27844 25774
rect 27804 24744 27856 24750
rect 27804 24686 27856 24692
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 26528 23730 26648 23746
rect 27436 23792 27488 23798
rect 27436 23734 27488 23740
rect 26516 23724 26648 23730
rect 26568 23718 26648 23724
rect 26516 23666 26568 23672
rect 27528 23656 27580 23662
rect 27528 23598 27580 23604
rect 27540 23254 27568 23598
rect 28092 23594 28120 25842
rect 28276 24410 28304 25842
rect 28356 25832 28408 25838
rect 28356 25774 28408 25780
rect 29552 25832 29604 25838
rect 29552 25774 29604 25780
rect 28368 24954 28396 25774
rect 28356 24948 28408 24954
rect 28356 24890 28408 24896
rect 28724 24948 28776 24954
rect 28724 24890 28776 24896
rect 28632 24608 28684 24614
rect 28632 24550 28684 24556
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28276 23866 28304 24346
rect 28644 24274 28672 24550
rect 28632 24268 28684 24274
rect 28632 24210 28684 24216
rect 28736 24206 28764 24890
rect 29564 24886 29592 25774
rect 29656 25362 29684 25842
rect 30196 25832 30248 25838
rect 30196 25774 30248 25780
rect 29644 25356 29696 25362
rect 29644 25298 29696 25304
rect 30208 25294 30236 25774
rect 30196 25288 30248 25294
rect 30196 25230 30248 25236
rect 29552 24880 29604 24886
rect 29552 24822 29604 24828
rect 29368 24744 29420 24750
rect 29368 24686 29420 24692
rect 29380 24274 29408 24686
rect 29368 24268 29420 24274
rect 29368 24210 29420 24216
rect 29564 24206 29592 24822
rect 30392 24818 30420 25910
rect 31116 25832 31168 25838
rect 31116 25774 31168 25780
rect 30656 25696 30708 25702
rect 30656 25638 30708 25644
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30472 25220 30524 25226
rect 30472 25162 30524 25168
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 28908 24200 28960 24206
rect 28908 24142 28960 24148
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 28264 23860 28316 23866
rect 28264 23802 28316 23808
rect 28920 23594 28948 24142
rect 27620 23588 27672 23594
rect 27620 23530 27672 23536
rect 28080 23588 28132 23594
rect 28080 23530 28132 23536
rect 28908 23588 28960 23594
rect 28908 23530 28960 23536
rect 27528 23248 27580 23254
rect 27528 23190 27580 23196
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 26148 23044 26200 23050
rect 26148 22986 26200 22992
rect 26160 22710 26188 22986
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26884 22976 26936 22982
rect 26884 22918 26936 22924
rect 26148 22704 26200 22710
rect 26148 22646 26200 22652
rect 26148 22568 26200 22574
rect 26068 22528 26148 22556
rect 26148 22510 26200 22516
rect 26252 22234 26280 22918
rect 26424 22568 26476 22574
rect 26424 22510 26476 22516
rect 25964 22228 26016 22234
rect 25964 22170 26016 22176
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26436 22166 26464 22510
rect 26424 22160 26476 22166
rect 26424 22102 26476 22108
rect 26896 22030 26924 22918
rect 26988 22574 27016 23122
rect 27632 23118 27660 23530
rect 29564 23118 29592 24142
rect 30392 24138 30420 24754
rect 30380 24132 30432 24138
rect 30380 24074 30432 24080
rect 30484 23798 30512 25162
rect 30472 23792 30524 23798
rect 30472 23734 30524 23740
rect 30196 23656 30248 23662
rect 30196 23598 30248 23604
rect 30208 23186 30236 23598
rect 30196 23180 30248 23186
rect 30196 23122 30248 23128
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 28632 23112 28684 23118
rect 28632 23054 28684 23060
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 27252 23044 27304 23050
rect 27252 22986 27304 22992
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 26988 22098 27016 22510
rect 27080 22438 27108 22714
rect 27264 22710 27292 22986
rect 27896 22976 27948 22982
rect 27896 22918 27948 22924
rect 27252 22704 27304 22710
rect 27252 22646 27304 22652
rect 27068 22432 27120 22438
rect 27068 22374 27120 22380
rect 27908 22234 27936 22918
rect 28644 22778 28672 23054
rect 28632 22772 28684 22778
rect 28632 22714 28684 22720
rect 29012 22642 29040 23054
rect 29368 22976 29420 22982
rect 29368 22918 29420 22924
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 29276 22568 29328 22574
rect 29276 22510 29328 22516
rect 27896 22228 27948 22234
rect 27896 22170 27948 22176
rect 29288 22098 29316 22510
rect 29380 22234 29408 22918
rect 30484 22438 30512 23734
rect 30576 23730 30604 25298
rect 30564 23724 30616 23730
rect 30564 23666 30616 23672
rect 30668 23662 30696 25638
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30852 24274 30880 24550
rect 31128 24342 31156 25774
rect 31404 25226 31432 26930
rect 31484 26920 31536 26926
rect 31484 26862 31536 26868
rect 31496 26586 31524 26862
rect 33152 26858 33180 27338
rect 33244 27130 33272 27610
rect 33232 27124 33284 27130
rect 33232 27066 33284 27072
rect 33692 26920 33744 26926
rect 33692 26862 33744 26868
rect 33140 26852 33192 26858
rect 33140 26794 33192 26800
rect 31484 26580 31536 26586
rect 31484 26522 31536 26528
rect 31496 26042 31524 26522
rect 33232 26444 33284 26450
rect 33232 26386 33284 26392
rect 32128 26308 32180 26314
rect 32128 26250 32180 26256
rect 31484 26036 31536 26042
rect 31484 25978 31536 25984
rect 32140 25838 32168 26250
rect 32404 26240 32456 26246
rect 32404 26182 32456 26188
rect 32416 25974 32444 26182
rect 32404 25968 32456 25974
rect 32404 25910 32456 25916
rect 32128 25832 32180 25838
rect 32128 25774 32180 25780
rect 31760 25696 31812 25702
rect 31760 25638 31812 25644
rect 31392 25220 31444 25226
rect 31392 25162 31444 25168
rect 31208 24812 31260 24818
rect 31208 24754 31260 24760
rect 31220 24410 31248 24754
rect 31208 24404 31260 24410
rect 31208 24346 31260 24352
rect 31116 24336 31168 24342
rect 31116 24278 31168 24284
rect 30840 24268 30892 24274
rect 30840 24210 30892 24216
rect 31772 24206 31800 25638
rect 32140 25294 32168 25774
rect 32128 25288 32180 25294
rect 32128 25230 32180 25236
rect 32140 24750 32168 25230
rect 32036 24744 32088 24750
rect 32036 24686 32088 24692
rect 32128 24744 32180 24750
rect 32128 24686 32180 24692
rect 32048 24274 32076 24686
rect 32140 24274 32168 24686
rect 32036 24268 32088 24274
rect 32036 24210 32088 24216
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 31760 24200 31812 24206
rect 31760 24142 31812 24148
rect 31772 23798 31800 24142
rect 31760 23792 31812 23798
rect 31760 23734 31812 23740
rect 30748 23724 30800 23730
rect 30748 23666 30800 23672
rect 30656 23656 30708 23662
rect 30656 23598 30708 23604
rect 30668 23322 30696 23598
rect 30656 23316 30708 23322
rect 30656 23258 30708 23264
rect 30760 22778 30788 23666
rect 32140 23186 32168 24210
rect 33048 24132 33100 24138
rect 33048 24074 33100 24080
rect 33060 23866 33088 24074
rect 33244 24070 33272 26386
rect 33704 26382 33732 26862
rect 33692 26376 33744 26382
rect 33692 26318 33744 26324
rect 33416 26240 33468 26246
rect 33416 26182 33468 26188
rect 33428 25362 33456 26182
rect 33704 26042 33732 26318
rect 33692 26036 33744 26042
rect 33692 25978 33744 25984
rect 33508 25900 33560 25906
rect 33508 25842 33560 25848
rect 33416 25356 33468 25362
rect 33416 25298 33468 25304
rect 33324 25220 33376 25226
rect 33324 25162 33376 25168
rect 33336 24750 33364 25162
rect 33520 24886 33548 25842
rect 33796 25294 33824 28426
rect 33888 26926 33916 29650
rect 34624 29646 34652 30670
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34624 29306 34652 29582
rect 34612 29300 34664 29306
rect 34612 29242 34664 29248
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 33968 28552 34020 28558
rect 33968 28494 34020 28500
rect 33980 27674 34008 28494
rect 35360 28490 35388 30670
rect 35348 28484 35400 28490
rect 35348 28426 35400 28432
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 33968 27668 34020 27674
rect 33968 27610 34020 27616
rect 33980 27130 34008 27610
rect 33968 27124 34020 27130
rect 33968 27066 34020 27072
rect 33876 26920 33928 26926
rect 33876 26862 33928 26868
rect 33888 26450 33916 26862
rect 34060 26852 34112 26858
rect 34060 26794 34112 26800
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 34072 25906 34100 26794
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34060 25900 34112 25906
rect 34060 25842 34112 25848
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34428 25356 34480 25362
rect 34428 25298 34480 25304
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 34440 24954 34468 25298
rect 34520 25220 34572 25226
rect 34520 25162 34572 25168
rect 34428 24948 34480 24954
rect 34428 24890 34480 24896
rect 33508 24880 33560 24886
rect 33508 24822 33560 24828
rect 33324 24744 33376 24750
rect 33324 24686 33376 24692
rect 33520 24138 33548 24822
rect 34532 24410 34560 25162
rect 35452 25158 35480 31826
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35440 25152 35492 25158
rect 35440 25094 35492 25100
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34520 24404 34572 24410
rect 34520 24346 34572 24352
rect 33508 24132 33560 24138
rect 33508 24074 33560 24080
rect 33232 24064 33284 24070
rect 33232 24006 33284 24012
rect 34060 24064 34112 24070
rect 34060 24006 34112 24012
rect 33048 23860 33100 23866
rect 33048 23802 33100 23808
rect 34072 23730 34100 24006
rect 34532 23866 34560 24346
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 33876 23724 33928 23730
rect 33876 23666 33928 23672
rect 34060 23724 34112 23730
rect 34060 23666 34112 23672
rect 32404 23656 32456 23662
rect 32404 23598 32456 23604
rect 33232 23656 33284 23662
rect 33232 23598 33284 23604
rect 32128 23180 32180 23186
rect 32128 23122 32180 23128
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 30748 22772 30800 22778
rect 30748 22714 30800 22720
rect 30012 22432 30064 22438
rect 30012 22374 30064 22380
rect 30472 22432 30524 22438
rect 30472 22374 30524 22380
rect 29368 22228 29420 22234
rect 29368 22170 29420 22176
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 29276 22092 29328 22098
rect 29276 22034 29328 22040
rect 30024 22030 30052 22374
rect 30760 22098 30788 22714
rect 31496 22710 31524 22918
rect 31484 22704 31536 22710
rect 31484 22646 31536 22652
rect 32140 22642 32168 23122
rect 32416 22710 32444 23598
rect 33244 23050 33272 23598
rect 33232 23044 33284 23050
rect 33232 22986 33284 22992
rect 33416 23044 33468 23050
rect 33416 22986 33468 22992
rect 33428 22710 33456 22986
rect 33888 22778 33916 23666
rect 34428 23656 34480 23662
rect 34428 23598 34480 23604
rect 34440 23322 34468 23598
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34428 23316 34480 23322
rect 34428 23258 34480 23264
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 33876 22772 33928 22778
rect 33876 22714 33928 22720
rect 32404 22704 32456 22710
rect 32404 22646 32456 22652
rect 33416 22704 33468 22710
rect 33416 22646 33468 22652
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 30748 22092 30800 22098
rect 33428 22094 33456 22646
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 30748 22034 30800 22040
rect 33336 22066 33456 22094
rect 26884 22024 26936 22030
rect 26884 21966 26936 21972
rect 30012 22024 30064 22030
rect 30012 21966 30064 21972
rect 26148 21956 26200 21962
rect 26148 21898 26200 21904
rect 27988 21956 28040 21962
rect 27988 21898 28040 21904
rect 25504 21888 25556 21894
rect 25504 21830 25556 21836
rect 23572 21072 23624 21078
rect 23572 21014 23624 21020
rect 22836 20936 22888 20942
rect 22836 20878 22888 20884
rect 22848 20806 22876 20878
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22848 20602 22876 20742
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 23584 20482 23612 21014
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 23676 20602 23704 20946
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 22572 20398 22600 20470
rect 23584 20454 23704 20482
rect 23676 20398 23704 20454
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19536 19922 19564 20198
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19536 18834 19564 19858
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19812 19446 19840 19722
rect 19800 19440 19852 19446
rect 19800 19382 19852 19388
rect 20824 19378 20852 20334
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22296 19854 22324 20198
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19076 16546 19196 16574
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18432 15570 18460 15846
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18616 14482 18644 16050
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18800 15570 18828 15982
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 19076 15162 19104 16546
rect 19352 16182 19380 16934
rect 19536 16250 19564 18770
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19812 18358 19840 18634
rect 20732 18630 20760 19314
rect 20916 18986 20944 19654
rect 21008 19378 21036 19654
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 20824 18958 20944 18986
rect 20824 18698 20852 18958
rect 20904 18896 20956 18902
rect 20904 18838 20956 18844
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20456 16794 20484 17138
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20732 16538 20760 18566
rect 20824 17490 20852 18634
rect 20916 17610 20944 18838
rect 21008 18358 21036 19314
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 21284 18222 21312 18566
rect 22296 18290 22324 19790
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22572 19514 22600 19722
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 23676 19242 23704 20334
rect 24964 20074 24992 20878
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 25148 20534 25176 20742
rect 26160 20602 26188 21898
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27632 21010 27660 21286
rect 28000 21010 28028 21898
rect 28356 21548 28408 21554
rect 28356 21490 28408 21496
rect 29552 21548 29604 21554
rect 29552 21490 29604 21496
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27988 21004 28040 21010
rect 27988 20946 28040 20952
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 26988 20602 27016 20878
rect 27068 20868 27120 20874
rect 27068 20810 27120 20816
rect 26148 20596 26200 20602
rect 26148 20538 26200 20544
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 25412 20392 25464 20398
rect 25412 20334 25464 20340
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 24872 20058 24992 20074
rect 24860 20052 24992 20058
rect 24912 20046 24992 20052
rect 24860 19994 24912 20000
rect 24872 19514 24900 19994
rect 25056 19786 25084 20198
rect 25424 19922 25452 20334
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 26160 19854 26188 20538
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26528 20058 26556 20402
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26988 19922 27016 20538
rect 26976 19916 27028 19922
rect 26976 19858 27028 19864
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 25136 19712 25188 19718
rect 25136 19654 25188 19660
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 25148 19514 25176 19654
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23664 19236 23716 19242
rect 23664 19178 23716 19184
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 21008 17490 21036 17546
rect 20824 17462 21036 17490
rect 21640 17536 21692 17542
rect 21640 17478 21692 17484
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20640 16522 20760 16538
rect 20628 16516 20760 16522
rect 20680 16510 20760 16516
rect 20628 16458 20680 16464
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18420 14340 18472 14346
rect 18420 14282 18472 14288
rect 18432 14006 18460 14282
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 11830 17080 13194
rect 18524 13190 18552 13806
rect 18616 13394 18644 14418
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17880 11830 17908 12038
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16408 10742 16436 11018
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 15488 9722 15516 9998
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15488 9466 15516 9658
rect 16132 9518 16160 9998
rect 16408 9994 16436 10678
rect 16776 10674 16804 11222
rect 17880 11098 17908 11766
rect 17696 11070 17908 11098
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10810 17632 10950
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16408 9654 16436 9930
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 15396 9438 15516 9466
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 15396 8974 15424 9438
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15488 8634 15516 8910
rect 16408 8906 16436 9590
rect 17420 9586 17448 10610
rect 17696 10606 17724 11070
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17880 10266 17908 10950
rect 17972 10742 18000 12106
rect 18064 11762 18092 12718
rect 18524 11762 18552 13126
rect 18616 12782 18644 13330
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18064 11234 18092 11698
rect 18616 11694 18644 12174
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18064 11206 18276 11234
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17880 9654 17908 10202
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 7954 14320 8230
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14292 6458 14320 7890
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14568 7478 14596 7754
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 15488 7426 15516 8570
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15672 7886 15700 8502
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15488 7410 15608 7426
rect 15200 7404 15252 7410
rect 15488 7404 15620 7410
rect 15488 7398 15568 7404
rect 15200 7346 15252 7352
rect 15568 7346 15620 7352
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14108 5234 14136 6326
rect 14844 6254 14872 6666
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 15212 5642 15240 7346
rect 15672 6390 15700 7822
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15396 5710 15424 6054
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 14384 5302 14412 5578
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14108 4690 14136 5170
rect 15580 4690 15608 5578
rect 15672 5302 15700 6326
rect 15764 6118 15792 6734
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15856 5370 15884 5714
rect 15948 5710 15976 8842
rect 16224 8634 16252 8842
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16408 8566 16436 8842
rect 16500 8566 16528 9522
rect 17868 9512 17920 9518
rect 17972 9500 18000 10406
rect 18064 9654 18092 10746
rect 18156 10130 18184 10950
rect 18248 10606 18276 11206
rect 18616 11150 18644 11630
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 18248 10130 18276 10542
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17920 9472 18000 9500
rect 17868 9454 17920 9460
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16684 8430 16712 8978
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16040 7410 16068 7686
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16040 6866 16068 7346
rect 16684 7342 16712 8366
rect 17236 7886 17264 9386
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17420 7478 17448 7754
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16684 6866 16712 7278
rect 16028 6860 16080 6866
rect 16672 6860 16724 6866
rect 16028 6802 16080 6808
rect 16592 6820 16672 6848
rect 16592 5778 16620 6820
rect 16672 6802 16724 6808
rect 17420 6730 17448 7414
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 16960 6390 16988 6666
rect 16948 6384 17000 6390
rect 16948 6326 17000 6332
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 17420 5642 17448 6666
rect 17880 6662 17908 9454
rect 18248 8974 18276 10066
rect 18432 10062 18460 10678
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18432 9722 18460 9998
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18708 8974 18736 10950
rect 18892 10674 18920 12786
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18708 8498 18736 8570
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18340 8090 18368 8298
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 17880 6186 17908 6598
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 17868 6180 17920 6186
rect 17868 6122 17920 6128
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15672 4554 15700 5238
rect 16776 5166 16804 5578
rect 16868 5302 16896 5578
rect 18156 5302 18184 6326
rect 18432 6322 18460 6598
rect 18524 6322 18552 7278
rect 18616 7206 18644 8434
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18800 7954 18828 8366
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18984 7546 19012 13874
rect 19076 10810 19104 15098
rect 19996 15094 20024 15982
rect 20732 15570 20760 16510
rect 20824 16250 20852 17206
rect 20916 16522 20944 17462
rect 21652 17066 21680 17478
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20824 15570 20852 16186
rect 20916 16046 20944 16458
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19996 13938 20024 15030
rect 20640 14346 20668 15438
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 15162 20760 15370
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 21468 14958 21496 15438
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19996 13258 20024 13874
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 19996 12918 20024 13194
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19628 12238 19656 12718
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 19076 10470 19104 10746
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19352 10062 19380 11630
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19536 10130 19564 11018
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19812 10062 19840 12174
rect 19996 11762 20024 12854
rect 21100 12850 21128 13194
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20732 12322 20760 12718
rect 20640 12294 20760 12322
rect 20640 12238 20668 12294
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19996 11082 20024 11698
rect 20272 11558 20300 12174
rect 20732 11694 20760 12174
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19812 9500 19840 9998
rect 19996 9722 20024 11018
rect 20088 10130 20116 11494
rect 21284 11218 21312 14282
rect 21468 14074 21496 14894
rect 21652 14278 21680 17002
rect 21836 16250 21864 17138
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 21928 16658 21956 16934
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21824 16244 21876 16250
rect 21876 16204 21956 16232
rect 21824 16186 21876 16192
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21836 15502 21864 16050
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15094 21864 15438
rect 21928 15366 21956 16204
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21836 14482 21864 15030
rect 21928 15026 21956 15302
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21836 13954 21864 14418
rect 21744 13938 21864 13954
rect 22020 13938 22048 18090
rect 22296 17746 22324 18226
rect 22388 17882 22416 18770
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22572 17882 22600 18158
rect 23676 18086 23704 19178
rect 23768 18222 23796 19246
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24136 18222 24164 18702
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22296 17270 22324 17682
rect 22388 17338 22416 17818
rect 23676 17746 23704 18022
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22296 16658 22324 17206
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22652 16516 22704 16522
rect 22652 16458 22704 16464
rect 22664 16182 22692 16458
rect 22652 16176 22704 16182
rect 22652 16118 22704 16124
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 23296 16108 23348 16114
rect 23296 16050 23348 16056
rect 23124 15570 23152 16050
rect 23308 15706 23336 16050
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 22112 15162 22140 15370
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 21732 13932 21864 13938
rect 21784 13926 21864 13932
rect 22008 13932 22060 13938
rect 21732 13874 21784 13880
rect 22008 13874 22060 13880
rect 21744 13394 21772 13874
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 21560 12170 21588 13194
rect 21744 12918 21772 13330
rect 22020 12986 22048 13874
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 21732 12912 21784 12918
rect 21732 12854 21784 12860
rect 22296 12850 22324 15302
rect 23308 15162 23336 15642
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23676 14958 23704 17682
rect 23768 17678 23796 18158
rect 24136 17678 24164 18158
rect 24780 17882 24808 18702
rect 25148 18222 25176 19450
rect 26068 19310 26096 19654
rect 26160 19514 26188 19790
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 26620 19446 26648 19722
rect 26608 19440 26660 19446
rect 26608 19382 26660 19388
rect 26988 19310 27016 19858
rect 27080 19854 27108 20810
rect 28000 20534 28028 20946
rect 28368 20806 28396 21490
rect 28724 21480 28776 21486
rect 28724 21422 28776 21428
rect 28356 20800 28408 20806
rect 28356 20742 28408 20748
rect 27988 20528 28040 20534
rect 27988 20470 28040 20476
rect 27712 20392 27764 20398
rect 27712 20334 27764 20340
rect 27724 19922 27752 20334
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 27068 19848 27120 19854
rect 27068 19790 27120 19796
rect 26056 19304 26108 19310
rect 26976 19304 27028 19310
rect 26108 19252 26188 19258
rect 26056 19246 26188 19252
rect 26976 19246 27028 19252
rect 26068 19230 26188 19246
rect 26160 18766 26188 19230
rect 26988 18766 27016 19246
rect 27080 19174 27108 19790
rect 28000 19514 28028 20470
rect 28368 19854 28396 20742
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28460 19922 28488 20198
rect 28448 19916 28500 19922
rect 28448 19858 28500 19864
rect 28356 19848 28408 19854
rect 28356 19790 28408 19796
rect 27988 19508 28040 19514
rect 27988 19450 28040 19456
rect 28000 19334 28028 19450
rect 28000 19306 28304 19334
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 27080 18970 27108 19110
rect 27068 18964 27120 18970
rect 27068 18906 27120 18912
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 18358 25636 18566
rect 25596 18352 25648 18358
rect 25596 18294 25648 18300
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 26252 17882 26280 18702
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 24124 17672 24176 17678
rect 24124 17614 24176 17620
rect 25596 17604 25648 17610
rect 25596 17546 25648 17552
rect 25608 17270 25636 17546
rect 26252 17338 26280 17682
rect 26344 17610 26372 18566
rect 26988 18222 27016 18702
rect 28276 18698 28304 19306
rect 27068 18692 27120 18698
rect 27068 18634 27120 18640
rect 28264 18692 28316 18698
rect 28264 18634 28316 18640
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26988 17678 27016 18158
rect 26976 17672 27028 17678
rect 26976 17614 27028 17620
rect 26332 17604 26384 17610
rect 26332 17546 26384 17552
rect 26884 17536 26936 17542
rect 26884 17478 26936 17484
rect 26896 17338 26924 17478
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 26884 17332 26936 17338
rect 26884 17274 26936 17280
rect 25596 17264 25648 17270
rect 25596 17206 25648 17212
rect 25608 16522 25636 17206
rect 26792 17128 26844 17134
rect 26792 17070 26844 17076
rect 26804 16794 26832 17070
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 25596 16516 25648 16522
rect 25596 16458 25648 16464
rect 23952 16182 23980 16458
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 23940 16176 23992 16182
rect 23860 16136 23940 16164
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23768 15094 23796 15982
rect 23860 15434 23888 16136
rect 23940 16118 23992 16124
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24412 15570 24440 15982
rect 25056 15910 25084 16390
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 25056 15502 25084 15846
rect 25516 15570 25544 15982
rect 25700 15978 25728 16730
rect 26148 16652 26200 16658
rect 26200 16612 26280 16640
rect 26148 16594 26200 16600
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 25976 16182 26004 16390
rect 25964 16176 26016 16182
rect 25964 16118 26016 16124
rect 25688 15972 25740 15978
rect 25688 15914 25740 15920
rect 25504 15564 25556 15570
rect 25504 15506 25556 15512
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 23848 15428 23900 15434
rect 23848 15370 23900 15376
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 23860 14346 23888 15370
rect 24400 15088 24452 15094
rect 24400 15030 24452 15036
rect 26148 15088 26200 15094
rect 26148 15030 26200 15036
rect 23940 14884 23992 14890
rect 23940 14826 23992 14832
rect 23952 14618 23980 14826
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 22756 14006 22784 14282
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22572 12850 22600 13466
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 20180 10062 20208 11154
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20076 9512 20128 9518
rect 19812 9472 20076 9500
rect 19812 8634 19840 9472
rect 20076 9454 20128 9460
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19812 8430 19840 8570
rect 20456 8498 20484 8978
rect 20640 8906 20668 9658
rect 20732 9654 20760 10406
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18984 6798 19012 7482
rect 19076 6866 19104 7822
rect 20548 7750 20576 8434
rect 20640 7818 20668 8842
rect 20824 8362 20852 10542
rect 21284 9586 21312 10610
rect 21376 10606 21404 11290
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21560 9994 21588 12106
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 21928 10130 21956 11630
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22112 10742 22140 11086
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 22204 10266 22232 10950
rect 22296 10606 22324 11086
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8498 21220 8842
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18984 6458 19012 6734
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18340 5574 18368 6190
rect 19076 5778 19104 6802
rect 19260 6322 19288 7142
rect 20456 6866 20484 7142
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19536 5778 19564 6666
rect 20456 6322 20484 6802
rect 20548 6662 20576 7686
rect 20640 7478 20668 7754
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 20536 5636 20588 5642
rect 20640 5624 20668 7414
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20916 6390 20944 7278
rect 21284 6798 21312 9522
rect 21928 9042 21956 10066
rect 22296 9518 22324 10542
rect 22572 10266 22600 11086
rect 22848 11082 22876 14214
rect 23952 13938 23980 14554
rect 24412 14482 24440 15030
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 24860 14884 24912 14890
rect 24860 14826 24912 14832
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 24676 14340 24728 14346
rect 24676 14282 24728 14288
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23032 12306 23060 13806
rect 23584 13530 23612 13874
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 24688 13394 24716 14282
rect 24872 13870 24900 14826
rect 25504 14816 25556 14822
rect 25504 14758 25556 14764
rect 25516 14006 25544 14758
rect 25504 14000 25556 14006
rect 25504 13942 25556 13948
rect 25976 13870 26004 14894
rect 26160 14278 26188 15030
rect 26252 14958 26280 16612
rect 26896 16590 26924 17274
rect 27080 16794 27108 18634
rect 28276 18358 28304 18634
rect 28264 18352 28316 18358
rect 28264 18294 28316 18300
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27632 17882 27660 18158
rect 28736 18086 28764 21422
rect 29564 21146 29592 21490
rect 30564 21480 30616 21486
rect 30564 21422 30616 21428
rect 31576 21480 31628 21486
rect 31576 21422 31628 21428
rect 32772 21480 32824 21486
rect 32772 21422 32824 21428
rect 29552 21140 29604 21146
rect 29552 21082 29604 21088
rect 30576 20602 30604 21422
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 31116 21344 31168 21350
rect 31116 21286 31168 21292
rect 31036 21010 31064 21286
rect 31024 21004 31076 21010
rect 31024 20946 31076 20952
rect 30748 20868 30800 20874
rect 30748 20810 30800 20816
rect 30564 20596 30616 20602
rect 30564 20538 30616 20544
rect 30760 20534 30788 20810
rect 31128 20534 31156 21286
rect 31588 21146 31616 21422
rect 31668 21344 31720 21350
rect 31668 21286 31720 21292
rect 31576 21140 31628 21146
rect 31576 21082 31628 21088
rect 30748 20528 30800 20534
rect 30748 20470 30800 20476
rect 31116 20528 31168 20534
rect 31116 20470 31168 20476
rect 30196 19848 30248 19854
rect 30196 19790 30248 19796
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 31116 19848 31168 19854
rect 31116 19790 31168 19796
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 29092 19780 29144 19786
rect 29092 19722 29144 19728
rect 29104 18630 29132 19722
rect 29276 19372 29328 19378
rect 29276 19314 29328 19320
rect 29092 18624 29144 18630
rect 29092 18566 29144 18572
rect 29000 18420 29052 18426
rect 29000 18362 29052 18368
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27804 16992 27856 16998
rect 27804 16934 27856 16940
rect 27068 16788 27120 16794
rect 27068 16730 27120 16736
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26344 15026 26372 15982
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 26252 14414 26280 14894
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24872 13326 24900 13806
rect 26160 13394 26188 14214
rect 26252 14074 26280 14350
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26240 14068 26292 14074
rect 26240 14010 26292 14016
rect 26240 13932 26292 13938
rect 26344 13920 26372 14214
rect 26528 14074 26556 14282
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 26292 13892 26372 13920
rect 26240 13874 26292 13880
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24964 12986 24992 13262
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 26252 12918 26280 13874
rect 26240 12912 26292 12918
rect 26240 12854 26292 12860
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 22928 12096 22980 12102
rect 22928 12038 22980 12044
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 22940 11218 22968 12038
rect 23124 11830 23152 12038
rect 23112 11824 23164 11830
rect 23112 11766 23164 11772
rect 23308 11286 23336 12242
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23860 11898 23888 12038
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 24596 11830 24624 12786
rect 25504 12776 25556 12782
rect 25504 12718 25556 12724
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24400 11688 24452 11694
rect 24400 11630 24452 11636
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 22928 11212 22980 11218
rect 22928 11154 22980 11160
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 23204 11076 23256 11082
rect 23204 11018 23256 11024
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 22848 8922 22876 11018
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22940 9042 22968 10406
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 21468 7954 21496 8910
rect 22848 8894 22968 8922
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21468 7410 21496 7890
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 22112 7342 22140 8366
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21560 6458 21588 6734
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 20588 5596 20668 5624
rect 20536 5578 20588 5584
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 16856 5296 16908 5302
rect 16856 5238 16908 5244
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 18340 5234 18368 5510
rect 20548 5234 20576 5578
rect 21560 5574 21588 6394
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 16776 4826 16804 5102
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 20824 4690 20852 5102
rect 21560 4758 21588 5510
rect 21744 5098 21772 6734
rect 21836 6254 21864 6734
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 21836 5914 21864 6190
rect 22112 6186 22140 7278
rect 22204 7002 22232 7686
rect 22192 6996 22244 7002
rect 22192 6938 22244 6944
rect 22468 6860 22520 6866
rect 22468 6802 22520 6808
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 22204 5386 22232 6258
rect 22480 6254 22508 6802
rect 22940 6798 22968 8894
rect 23032 8566 23060 9998
rect 23216 9654 23244 11018
rect 23308 10538 23336 11222
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 23400 10062 23428 11018
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23400 9042 23428 9590
rect 23584 9586 23612 10066
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23676 9178 23704 10610
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23572 9036 23624 9042
rect 23572 8978 23624 8984
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 23400 7970 23428 8978
rect 23584 8430 23612 8978
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 23308 7942 23428 7970
rect 23308 7886 23336 7942
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23308 7478 23336 7822
rect 23296 7472 23348 7478
rect 23296 7414 23348 7420
rect 23400 7206 23428 7822
rect 23584 7546 23612 8366
rect 23676 7954 23704 9114
rect 23860 8974 23888 10746
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23860 8498 23888 8910
rect 23952 8548 23980 10406
rect 24412 10130 24440 11630
rect 24688 11354 24716 11630
rect 25056 11558 25084 12038
rect 25516 11898 25544 12718
rect 26056 12708 26108 12714
rect 26056 12650 26108 12656
rect 26068 12306 26096 12650
rect 26056 12300 26108 12306
rect 26056 12242 26108 12248
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25964 11824 26016 11830
rect 25964 11766 26016 11772
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 25056 11150 25084 11494
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 25148 10674 25176 10950
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24688 10130 24716 10406
rect 25148 10266 25176 10610
rect 25332 10606 25360 11154
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 25976 9994 26004 11766
rect 26068 10606 26096 12242
rect 26252 11830 26280 12854
rect 26620 12170 26648 16186
rect 27080 15434 27108 16730
rect 27816 16658 27844 16934
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27540 16182 27568 16594
rect 27528 16176 27580 16182
rect 27528 16118 27580 16124
rect 27908 15570 27936 18022
rect 29012 17746 29040 18362
rect 29000 17740 29052 17746
rect 29000 17682 29052 17688
rect 28172 17604 28224 17610
rect 28172 17546 28224 17552
rect 28724 17604 28776 17610
rect 28724 17546 28776 17552
rect 28184 16250 28212 17546
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28184 15910 28212 16186
rect 28540 16040 28592 16046
rect 28736 16028 28764 17546
rect 28816 17264 28868 17270
rect 28816 17206 28868 17212
rect 28592 16000 28764 16028
rect 28540 15982 28592 15988
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28736 15570 28764 16000
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 27068 15428 27120 15434
rect 27068 15370 27120 15376
rect 27620 15360 27672 15366
rect 27620 15302 27672 15308
rect 27632 15094 27660 15302
rect 27620 15088 27672 15094
rect 27620 15030 27672 15036
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27816 14346 27844 15030
rect 27804 14340 27856 14346
rect 27804 14282 27856 14288
rect 27908 13802 27936 15506
rect 28828 15502 28856 17206
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 29012 16182 29040 17138
rect 29288 16522 29316 19314
rect 29460 19168 29512 19174
rect 29460 19110 29512 19116
rect 29276 16516 29328 16522
rect 29276 16458 29328 16464
rect 29092 16244 29144 16250
rect 29092 16186 29144 16192
rect 29000 16176 29052 16182
rect 29000 16118 29052 16124
rect 28908 16040 28960 16046
rect 28908 15982 28960 15988
rect 28920 15706 28948 15982
rect 28908 15700 28960 15706
rect 28908 15642 28960 15648
rect 29012 15570 29040 16118
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28080 15360 28132 15366
rect 28080 15302 28132 15308
rect 28092 14618 28120 15302
rect 28828 15162 28856 15438
rect 29104 15434 29132 16186
rect 29288 16046 29316 16458
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29092 15428 29144 15434
rect 29092 15370 29144 15376
rect 28816 15156 28868 15162
rect 28816 15098 28868 15104
rect 28080 14612 28132 14618
rect 28080 14554 28132 14560
rect 28092 14074 28120 14554
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 29288 13870 29316 15982
rect 28908 13864 28960 13870
rect 28908 13806 28960 13812
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 27896 13796 27948 13802
rect 27896 13738 27948 13744
rect 28080 13456 28132 13462
rect 28080 13398 28132 13404
rect 27712 13252 27764 13258
rect 27712 13194 27764 13200
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 26976 12776 27028 12782
rect 26976 12718 27028 12724
rect 26608 12164 26660 12170
rect 26608 12106 26660 12112
rect 26332 12096 26384 12102
rect 26332 12038 26384 12044
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26148 10668 26200 10674
rect 26148 10610 26200 10616
rect 26056 10600 26108 10606
rect 26056 10542 26108 10548
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9654 24992 9862
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 25136 9648 25188 9654
rect 25136 9590 25188 9596
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24688 9178 24716 9454
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24584 8900 24636 8906
rect 24584 8842 24636 8848
rect 24032 8560 24084 8566
rect 23952 8520 24032 8548
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23768 7818 23796 8434
rect 23952 7954 23980 8520
rect 24032 8502 24084 8508
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23940 7948 23992 7954
rect 23940 7890 23992 7896
rect 23756 7812 23808 7818
rect 23756 7754 23808 7760
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 24044 7478 24072 8366
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 22940 6390 22968 6734
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 23400 6254 23428 7142
rect 24136 6866 24164 7890
rect 24596 7478 24624 8842
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 23112 6248 23164 6254
rect 23112 6190 23164 6196
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 22296 5778 22324 6190
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 23124 5710 23152 6190
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 22284 5636 22336 5642
rect 22284 5578 22336 5584
rect 22112 5358 22232 5386
rect 22112 5166 22140 5358
rect 22296 5234 22324 5578
rect 23124 5370 23152 5646
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23308 5302 23336 6054
rect 24412 5778 24440 6190
rect 24400 5772 24452 5778
rect 24400 5714 24452 5720
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23296 5296 23348 5302
rect 23296 5238 23348 5244
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21548 4752 21600 4758
rect 21548 4694 21600 4700
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 21744 4622 21772 5034
rect 22112 4690 22140 5102
rect 23860 5030 23888 5646
rect 24688 5302 24716 6258
rect 24872 5710 24900 8910
rect 25148 7954 25176 9590
rect 26068 9042 26096 10542
rect 26160 9722 26188 10610
rect 26252 10606 26280 11086
rect 26344 10810 26372 12038
rect 26620 11014 26648 12106
rect 26988 11286 27016 12718
rect 27356 12102 27384 12786
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27436 12096 27488 12102
rect 27436 12038 27488 12044
rect 27448 11830 27476 12038
rect 27724 11898 27752 13194
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 27436 11824 27488 11830
rect 27436 11766 27488 11772
rect 26976 11280 27028 11286
rect 26976 11222 27028 11228
rect 27724 11218 27752 11834
rect 28092 11694 28120 13398
rect 28920 13394 28948 13806
rect 28908 13388 28960 13394
rect 28908 13330 28960 13336
rect 29000 13252 29052 13258
rect 29000 13194 29052 13200
rect 29012 12986 29040 13194
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 28356 12640 28408 12646
rect 28356 12582 28408 12588
rect 28368 12306 28396 12582
rect 28356 12300 28408 12306
rect 28356 12242 28408 12248
rect 28448 12164 28500 12170
rect 28448 12106 28500 12112
rect 28460 11830 28488 12106
rect 29000 12096 29052 12102
rect 29000 12038 29052 12044
rect 29012 11898 29040 12038
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 28448 11824 28500 11830
rect 28448 11766 28500 11772
rect 28080 11688 28132 11694
rect 28080 11630 28132 11636
rect 28460 11218 28488 11766
rect 27712 11212 27764 11218
rect 27712 11154 27764 11160
rect 28448 11212 28500 11218
rect 28448 11154 28500 11160
rect 26608 11008 26660 11014
rect 26608 10950 26660 10956
rect 26332 10804 26384 10810
rect 26332 10746 26384 10752
rect 26620 10674 26648 10950
rect 26608 10668 26660 10674
rect 26608 10610 26660 10616
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26976 10600 27028 10606
rect 26976 10542 27028 10548
rect 26148 9716 26200 9722
rect 26148 9658 26200 9664
rect 26056 9036 26108 9042
rect 26056 8978 26108 8984
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25148 7818 25176 7890
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 25136 7812 25188 7818
rect 25136 7754 25188 7760
rect 24964 6866 24992 7754
rect 25148 7478 25176 7754
rect 25608 7546 25636 8910
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25976 8090 26004 8774
rect 26068 8378 26096 8978
rect 26160 8974 26188 9658
rect 26252 9654 26280 10542
rect 26700 10532 26752 10538
rect 26700 10474 26752 10480
rect 26712 9654 26740 10474
rect 26792 10464 26844 10470
rect 26792 10406 26844 10412
rect 26804 9654 26832 10406
rect 26988 10062 27016 10542
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26240 9648 26292 9654
rect 26240 9590 26292 9596
rect 26700 9648 26752 9654
rect 26700 9590 26752 9596
rect 26792 9648 26844 9654
rect 26792 9590 26844 9596
rect 26712 9178 26740 9590
rect 26988 9518 27016 9998
rect 26976 9512 27028 9518
rect 26976 9454 27028 9460
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 26712 8566 26740 9114
rect 26988 9042 27016 9454
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27632 8566 27660 8774
rect 28000 8634 28028 10610
rect 28460 10606 28488 11154
rect 29012 11082 29040 11834
rect 29000 11076 29052 11082
rect 29000 11018 29052 11024
rect 28632 10736 28684 10742
rect 28632 10678 28684 10684
rect 28448 10600 28500 10606
rect 28448 10542 28500 10548
rect 28644 9722 28672 10678
rect 28724 10600 28776 10606
rect 28724 10542 28776 10548
rect 28736 10266 28764 10542
rect 28724 10260 28776 10266
rect 28724 10202 28776 10208
rect 28632 9716 28684 9722
rect 28632 9658 28684 9664
rect 28356 9580 28408 9586
rect 28356 9522 28408 9528
rect 28724 9580 28776 9586
rect 28724 9522 28776 9528
rect 28368 8974 28396 9522
rect 28736 9178 28764 9522
rect 29288 9518 29316 13806
rect 29276 9512 29328 9518
rect 29276 9454 29328 9460
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28724 9172 28776 9178
rect 28724 9114 28776 9120
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 26700 8560 26752 8566
rect 26700 8502 26752 8508
rect 27620 8560 27672 8566
rect 27620 8502 27672 8508
rect 27528 8424 27580 8430
rect 26068 8362 26280 8378
rect 27528 8366 27580 8372
rect 26068 8356 26292 8362
rect 26068 8350 26240 8356
rect 26240 8298 26292 8304
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 25688 7948 25740 7954
rect 25688 7890 25740 7896
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 25608 6798 25636 7482
rect 25320 6792 25372 6798
rect 25320 6734 25372 6740
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 25148 5778 25176 6054
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 24412 4690 24440 5102
rect 24964 5030 24992 5646
rect 25148 5522 25176 5714
rect 25056 5494 25176 5522
rect 24492 5024 24544 5030
rect 24492 4966 24544 4972
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24504 4690 24532 4966
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 24964 2650 24992 4966
rect 25056 4622 25084 5494
rect 25044 4616 25096 4622
rect 25044 4558 25096 4564
rect 25332 4554 25360 6734
rect 25700 6458 25728 7890
rect 25976 6866 26004 8026
rect 27540 7954 27568 8366
rect 27632 7954 27660 8502
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27540 7818 27568 7890
rect 27528 7812 27580 7818
rect 27356 7772 27528 7800
rect 26976 7200 27028 7206
rect 26976 7142 27028 7148
rect 26988 7002 27016 7142
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 25964 6860 26016 6866
rect 25964 6802 26016 6808
rect 27356 6798 27384 7772
rect 27528 7754 27580 7760
rect 27632 7410 27660 7890
rect 27620 7404 27672 7410
rect 27620 7346 27672 7352
rect 27528 7336 27580 7342
rect 27724 7290 27752 8298
rect 27908 7750 27936 8434
rect 28368 8430 28396 8910
rect 28736 8566 28764 9114
rect 28828 9042 28856 9318
rect 28816 9036 28868 9042
rect 28816 8978 28868 8984
rect 29472 8906 29500 19110
rect 30208 18426 30236 19790
rect 30300 18970 30328 19790
rect 30380 19780 30432 19786
rect 30380 19722 30432 19728
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 30392 18834 30420 19722
rect 30472 19508 30524 19514
rect 30472 19450 30524 19456
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 30484 17610 30512 19450
rect 31128 19378 31156 19790
rect 31116 19372 31168 19378
rect 31116 19314 31168 19320
rect 30840 18692 30892 18698
rect 30840 18634 30892 18640
rect 30852 17610 30880 18634
rect 30932 18284 30984 18290
rect 30932 18226 30984 18232
rect 30472 17604 30524 17610
rect 30472 17546 30524 17552
rect 30840 17604 30892 17610
rect 30840 17546 30892 17552
rect 30852 17354 30880 17546
rect 30668 17326 30880 17354
rect 30668 17270 30696 17326
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 29552 17196 29604 17202
rect 29552 17138 29604 17144
rect 29564 16794 29592 17138
rect 29828 17128 29880 17134
rect 29828 17070 29880 17076
rect 29552 16788 29604 16794
rect 29552 16730 29604 16736
rect 29564 15366 29592 16730
rect 29840 16454 29868 17070
rect 30668 16590 30696 17206
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 29828 16448 29880 16454
rect 29828 16390 29880 16396
rect 29920 16448 29972 16454
rect 29920 16390 29972 16396
rect 29932 15910 29960 16390
rect 30668 16182 30696 16526
rect 30656 16176 30708 16182
rect 30656 16118 30708 16124
rect 29920 15904 29972 15910
rect 29920 15846 29972 15852
rect 30668 15450 30696 16118
rect 30840 16040 30892 16046
rect 30840 15982 30892 15988
rect 30576 15434 30696 15450
rect 30564 15428 30696 15434
rect 30616 15422 30696 15428
rect 30564 15370 30616 15376
rect 29552 15360 29604 15366
rect 29552 15302 29604 15308
rect 30472 15360 30524 15366
rect 30472 15302 30524 15308
rect 30484 15162 30512 15302
rect 30472 15156 30524 15162
rect 30472 15098 30524 15104
rect 30668 15094 30696 15422
rect 30852 15366 30880 15982
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30656 15088 30708 15094
rect 30656 15030 30708 15036
rect 30668 14346 30696 15030
rect 30852 14958 30880 15302
rect 30840 14952 30892 14958
rect 30840 14894 30892 14900
rect 30656 14340 30708 14346
rect 30656 14282 30708 14288
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29552 13864 29604 13870
rect 29552 13806 29604 13812
rect 29564 13258 29592 13806
rect 29552 13252 29604 13258
rect 29552 13194 29604 13200
rect 29656 12986 29684 13874
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 29644 12980 29696 12986
rect 29644 12922 29696 12928
rect 29656 12442 29684 12922
rect 29920 12912 29972 12918
rect 30116 12900 30144 13262
rect 30300 12918 30328 13806
rect 30668 13326 30696 14282
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30748 13184 30800 13190
rect 30748 13126 30800 13132
rect 29972 12872 30144 12900
rect 29920 12854 29972 12860
rect 29644 12436 29696 12442
rect 29644 12378 29696 12384
rect 30116 12186 30144 12872
rect 30288 12912 30340 12918
rect 30288 12854 30340 12860
rect 30760 12850 30788 13126
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 30564 12776 30616 12782
rect 30564 12718 30616 12724
rect 30576 12306 30604 12718
rect 30564 12300 30616 12306
rect 30564 12242 30616 12248
rect 30024 12170 30144 12186
rect 30012 12164 30144 12170
rect 30064 12158 30144 12164
rect 30012 12106 30064 12112
rect 30024 11898 30052 12106
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 30024 10742 30052 11834
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30380 11212 30432 11218
rect 30380 11154 30432 11160
rect 30392 10810 30420 11154
rect 30380 10804 30432 10810
rect 30380 10746 30432 10752
rect 30852 10742 30880 11494
rect 30012 10736 30064 10742
rect 30012 10678 30064 10684
rect 30840 10736 30892 10742
rect 30840 10678 30892 10684
rect 30380 10464 30432 10470
rect 30380 10406 30432 10412
rect 29644 10056 29696 10062
rect 29644 9998 29696 10004
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 29564 9042 29592 9454
rect 29656 9178 29684 9998
rect 29828 9920 29880 9926
rect 29828 9862 29880 9868
rect 29840 9586 29868 9862
rect 30208 9722 30236 9998
rect 30392 9994 30420 10406
rect 30380 9988 30432 9994
rect 30380 9930 30432 9936
rect 30196 9716 30248 9722
rect 30196 9658 30248 9664
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 29736 9512 29788 9518
rect 29736 9454 29788 9460
rect 29644 9172 29696 9178
rect 29644 9114 29696 9120
rect 29552 9036 29604 9042
rect 29552 8978 29604 8984
rect 29460 8900 29512 8906
rect 29460 8842 29512 8848
rect 29748 8566 29776 9454
rect 30196 9104 30248 9110
rect 30196 9046 30248 9052
rect 28724 8560 28776 8566
rect 28724 8502 28776 8508
rect 29736 8560 29788 8566
rect 29736 8502 29788 8508
rect 30208 8430 30236 9046
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 29460 8424 29512 8430
rect 29460 8366 29512 8372
rect 30196 8424 30248 8430
rect 30196 8366 30248 8372
rect 27988 8288 28040 8294
rect 27988 8230 28040 8236
rect 28000 7818 28028 8230
rect 27988 7812 28040 7818
rect 27988 7754 28040 7760
rect 27896 7744 27948 7750
rect 27896 7686 27948 7692
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 27908 7546 27936 7686
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 28460 7478 28488 7686
rect 27804 7472 27856 7478
rect 27804 7414 27856 7420
rect 28448 7472 28500 7478
rect 28448 7414 28500 7420
rect 27580 7284 27752 7290
rect 27528 7278 27752 7284
rect 27540 7262 27752 7278
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 27344 6792 27396 6798
rect 27344 6734 27396 6740
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 26068 5778 26096 6734
rect 27160 6112 27212 6118
rect 27160 6054 27212 6060
rect 26056 5772 26108 5778
rect 26056 5714 26108 5720
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25424 5234 25452 5646
rect 27172 5302 27200 6054
rect 27356 5710 27384 6734
rect 27724 6254 27752 7262
rect 27816 7002 27844 7414
rect 28172 7404 28224 7410
rect 28172 7346 28224 7352
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 27436 6248 27488 6254
rect 27436 6190 27488 6196
rect 27712 6248 27764 6254
rect 27712 6190 27764 6196
rect 27448 5846 27476 6190
rect 27436 5840 27488 5846
rect 27436 5782 27488 5788
rect 27816 5778 27844 6938
rect 28184 6866 28212 7346
rect 28172 6860 28224 6866
rect 28172 6802 28224 6808
rect 28184 6254 28212 6802
rect 28540 6384 28592 6390
rect 28540 6326 28592 6332
rect 28080 6248 28132 6254
rect 28080 6190 28132 6196
rect 28172 6248 28224 6254
rect 28172 6190 28224 6196
rect 28092 5778 28120 6190
rect 27804 5772 27856 5778
rect 27804 5714 27856 5720
rect 28080 5772 28132 5778
rect 28080 5714 28132 5720
rect 27344 5704 27396 5710
rect 27344 5646 27396 5652
rect 28184 5370 28212 6190
rect 28552 5710 28580 6326
rect 29472 6186 29500 8366
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 29932 7886 29960 8230
rect 30208 7954 30236 8366
rect 30196 7948 30248 7954
rect 30116 7908 30196 7936
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 29736 7472 29788 7478
rect 29736 7414 29788 7420
rect 29748 6662 29776 7414
rect 29932 6914 29960 7822
rect 30116 7546 30144 7908
rect 30196 7890 30248 7896
rect 30196 7744 30248 7750
rect 30196 7686 30248 7692
rect 30104 7540 30156 7546
rect 30104 7482 30156 7488
rect 30012 7336 30064 7342
rect 30012 7278 30064 7284
rect 29840 6886 29960 6914
rect 29736 6656 29788 6662
rect 29736 6598 29788 6604
rect 29748 6458 29776 6598
rect 29736 6452 29788 6458
rect 29736 6394 29788 6400
rect 29460 6180 29512 6186
rect 29460 6122 29512 6128
rect 28540 5704 28592 5710
rect 28540 5646 28592 5652
rect 28552 5370 28580 5646
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 28540 5364 28592 5370
rect 28540 5306 28592 5312
rect 27160 5296 27212 5302
rect 27160 5238 27212 5244
rect 25412 5228 25464 5234
rect 25412 5170 25464 5176
rect 25320 4548 25372 4554
rect 25320 4490 25372 4496
rect 28184 4146 28212 5306
rect 29564 5234 29592 5510
rect 29748 5302 29776 6394
rect 29840 5642 29868 6886
rect 30024 6866 30052 7278
rect 30208 7154 30236 7686
rect 30300 7410 30328 9522
rect 30392 8956 30420 9930
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30472 8968 30524 8974
rect 30392 8928 30472 8956
rect 30472 8910 30524 8916
rect 30564 8900 30616 8906
rect 30564 8842 30616 8848
rect 30656 8900 30708 8906
rect 30760 8888 30788 9522
rect 30708 8860 30788 8888
rect 30656 8842 30708 8848
rect 30576 7818 30604 8842
rect 30668 7954 30696 8842
rect 30840 8832 30892 8838
rect 30840 8774 30892 8780
rect 30852 8430 30880 8774
rect 30944 8650 30972 18226
rect 31128 12850 31156 19314
rect 31300 19304 31352 19310
rect 31404 19292 31432 19790
rect 31680 19334 31708 21286
rect 32784 21146 32812 21422
rect 32956 21344 33008 21350
rect 32956 21286 33008 21292
rect 32772 21140 32824 21146
rect 32772 21082 32824 21088
rect 31760 21004 31812 21010
rect 31760 20946 31812 20952
rect 31772 20398 31800 20946
rect 32784 20602 32812 21082
rect 32968 20874 32996 21286
rect 32864 20868 32916 20874
rect 32864 20810 32916 20816
rect 32956 20868 33008 20874
rect 32956 20810 33008 20816
rect 32876 20602 32904 20810
rect 32772 20596 32824 20602
rect 32772 20538 32824 20544
rect 32864 20596 32916 20602
rect 32864 20538 32916 20544
rect 33336 20534 33364 22066
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 33416 20936 33468 20942
rect 33416 20878 33468 20884
rect 33968 20936 34020 20942
rect 33968 20878 34020 20884
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 33324 20528 33376 20534
rect 33324 20470 33376 20476
rect 31760 20392 31812 20398
rect 31760 20334 31812 20340
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 31772 19530 31800 20334
rect 31772 19502 31892 19530
rect 31680 19310 31800 19334
rect 31680 19306 31812 19310
rect 31352 19264 31432 19292
rect 31760 19304 31812 19306
rect 31300 19246 31352 19252
rect 31760 19246 31812 19252
rect 31312 18970 31340 19246
rect 31300 18964 31352 18970
rect 31300 18906 31352 18912
rect 31864 18834 31892 19502
rect 31944 19372 31996 19378
rect 31944 19314 31996 19320
rect 31852 18828 31904 18834
rect 31852 18770 31904 18776
rect 31208 18216 31260 18222
rect 31208 18158 31260 18164
rect 31760 18216 31812 18222
rect 31760 18158 31812 18164
rect 31220 16998 31248 18158
rect 31576 18148 31628 18154
rect 31576 18090 31628 18096
rect 31208 16992 31260 16998
rect 31208 16934 31260 16940
rect 31392 15428 31444 15434
rect 31392 15370 31444 15376
rect 31300 15020 31352 15026
rect 31300 14962 31352 14968
rect 31116 12844 31168 12850
rect 31116 12786 31168 12792
rect 31024 12776 31076 12782
rect 31024 12718 31076 12724
rect 31036 12170 31064 12718
rect 31024 12164 31076 12170
rect 31024 12106 31076 12112
rect 31208 11620 31260 11626
rect 31208 11562 31260 11568
rect 31116 11552 31168 11558
rect 31116 11494 31168 11500
rect 31128 11354 31156 11494
rect 31116 11348 31168 11354
rect 31116 11290 31168 11296
rect 31220 10606 31248 11562
rect 31208 10600 31260 10606
rect 31208 10542 31260 10548
rect 31220 10130 31248 10542
rect 31208 10124 31260 10130
rect 31208 10066 31260 10072
rect 31312 9586 31340 14962
rect 31404 14482 31432 15370
rect 31588 15366 31616 18090
rect 31772 17270 31800 18158
rect 31864 17746 31892 18770
rect 31956 18358 31984 19314
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 31944 18352 31996 18358
rect 31944 18294 31996 18300
rect 31956 17882 31984 18294
rect 32128 18216 32180 18222
rect 32128 18158 32180 18164
rect 31944 17876 31996 17882
rect 31944 17818 31996 17824
rect 31852 17740 31904 17746
rect 31852 17682 31904 17688
rect 31864 17626 31892 17682
rect 31864 17598 31984 17626
rect 31760 17264 31812 17270
rect 31760 17206 31812 17212
rect 31956 17202 31984 17598
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 32140 17134 32168 18158
rect 33048 17672 33100 17678
rect 33048 17614 33100 17620
rect 33060 17134 33088 17614
rect 32128 17128 32180 17134
rect 32128 17070 32180 17076
rect 32404 17128 32456 17134
rect 32404 17070 32456 17076
rect 33048 17128 33100 17134
rect 33048 17070 33100 17076
rect 31944 16992 31996 16998
rect 31996 16940 32076 16946
rect 31944 16934 32076 16940
rect 31956 16918 32076 16934
rect 31680 16782 31984 16810
rect 31680 16522 31708 16782
rect 31760 16720 31812 16726
rect 31760 16662 31812 16668
rect 31668 16516 31720 16522
rect 31668 16458 31720 16464
rect 31576 15360 31628 15366
rect 31576 15302 31628 15308
rect 31392 14476 31444 14482
rect 31392 14418 31444 14424
rect 31680 14074 31708 16458
rect 31772 16114 31800 16662
rect 31956 16590 31984 16782
rect 32048 16658 32076 16918
rect 32140 16726 32168 17070
rect 32128 16720 32180 16726
rect 32128 16662 32180 16668
rect 32416 16658 32444 17070
rect 33060 16658 33088 17070
rect 32036 16652 32088 16658
rect 32036 16594 32088 16600
rect 32404 16652 32456 16658
rect 32404 16594 32456 16600
rect 33048 16652 33100 16658
rect 33048 16594 33100 16600
rect 31944 16584 31996 16590
rect 31944 16526 31996 16532
rect 31760 16108 31812 16114
rect 31760 16050 31812 16056
rect 31772 14822 31800 16050
rect 33152 16046 33180 19246
rect 33244 19174 33272 20334
rect 33232 19168 33284 19174
rect 33232 19110 33284 19116
rect 33324 18828 33376 18834
rect 33324 18770 33376 18776
rect 33336 17882 33364 18770
rect 33428 18222 33456 20878
rect 33508 20868 33560 20874
rect 33508 20810 33560 20816
rect 33520 20534 33548 20810
rect 33980 20806 34008 20878
rect 33968 20800 34020 20806
rect 33968 20742 34020 20748
rect 33508 20528 33560 20534
rect 33508 20470 33560 20476
rect 34164 20466 34192 20878
rect 34980 20868 35032 20874
rect 34980 20810 35032 20816
rect 35440 20868 35492 20874
rect 35440 20810 35492 20816
rect 34428 20800 34480 20806
rect 34428 20742 34480 20748
rect 34440 20466 34468 20742
rect 34992 20534 35020 20810
rect 35452 20602 35480 20810
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35440 20596 35492 20602
rect 35440 20538 35492 20544
rect 34980 20528 35032 20534
rect 34980 20470 35032 20476
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 34428 20460 34480 20466
rect 34428 20402 34480 20408
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34164 19514 34192 20402
rect 34532 19922 34560 20402
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34520 19916 34572 19922
rect 34520 19858 34572 19864
rect 34532 19514 34560 19858
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 34152 19508 34204 19514
rect 34152 19450 34204 19456
rect 34520 19508 34572 19514
rect 34520 19450 34572 19456
rect 34716 19310 34744 19722
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18986 35388 19790
rect 35452 19378 35480 20538
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35440 19372 35492 19378
rect 35440 19314 35492 19320
rect 35268 18958 35388 18986
rect 35268 18766 35296 18958
rect 35348 18896 35400 18902
rect 35348 18838 35400 18844
rect 35256 18760 35308 18766
rect 35256 18702 35308 18708
rect 33600 18692 33652 18698
rect 33600 18634 33652 18640
rect 34796 18692 34848 18698
rect 34796 18634 34848 18640
rect 33612 18358 33640 18634
rect 33784 18624 33836 18630
rect 33784 18566 33836 18572
rect 33600 18352 33652 18358
rect 33600 18294 33652 18300
rect 33416 18216 33468 18222
rect 33416 18158 33468 18164
rect 33324 17876 33376 17882
rect 33324 17818 33376 17824
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33428 16998 33456 17614
rect 33612 17354 33640 18294
rect 33796 17746 33824 18566
rect 34808 17746 34836 18634
rect 35268 18222 35296 18702
rect 35360 18426 35388 18838
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35256 18216 35308 18222
rect 35256 18158 35308 18164
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 33784 17740 33836 17746
rect 33784 17682 33836 17688
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 34060 17536 34112 17542
rect 34060 17478 34112 17484
rect 33520 17326 33640 17354
rect 34072 17338 34100 17478
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 33520 17202 33548 17326
rect 33508 17196 33560 17202
rect 33508 17138 33560 17144
rect 33416 16992 33468 16998
rect 33416 16934 33468 16940
rect 33508 16992 33560 16998
rect 33508 16934 33560 16940
rect 31944 16040 31996 16046
rect 31944 15982 31996 15988
rect 32772 16040 32824 16046
rect 32772 15982 32824 15988
rect 33140 16040 33192 16046
rect 33140 15982 33192 15988
rect 31956 15638 31984 15982
rect 32220 15904 32272 15910
rect 32220 15846 32272 15852
rect 31944 15632 31996 15638
rect 31944 15574 31996 15580
rect 32036 15632 32088 15638
rect 32036 15574 32088 15580
rect 31956 15502 31984 15574
rect 31944 15496 31996 15502
rect 31944 15438 31996 15444
rect 31760 14816 31812 14822
rect 31760 14758 31812 14764
rect 31772 14482 31800 14758
rect 32048 14482 32076 15574
rect 32232 15570 32260 15846
rect 32220 15564 32272 15570
rect 32220 15506 32272 15512
rect 32128 15496 32180 15502
rect 32128 15438 32180 15444
rect 32140 14618 32168 15438
rect 32784 15162 32812 15982
rect 33428 15502 33456 16934
rect 33520 16794 33548 16934
rect 33508 16788 33560 16794
rect 33508 16730 33560 16736
rect 33520 16250 33548 16730
rect 33508 16244 33560 16250
rect 33508 16186 33560 16192
rect 33508 15564 33560 15570
rect 33508 15506 33560 15512
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 32772 15156 32824 15162
rect 32772 15098 32824 15104
rect 32864 14952 32916 14958
rect 32864 14894 32916 14900
rect 32128 14612 32180 14618
rect 32128 14554 32180 14560
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 32036 14476 32088 14482
rect 32036 14418 32088 14424
rect 31668 14068 31720 14074
rect 31668 14010 31720 14016
rect 32588 14068 32640 14074
rect 32588 14010 32640 14016
rect 32036 13932 32088 13938
rect 32036 13874 32088 13880
rect 31392 12300 31444 12306
rect 31392 12242 31444 12248
rect 31404 11218 31432 12242
rect 31668 11688 31720 11694
rect 31668 11630 31720 11636
rect 31760 11688 31812 11694
rect 31760 11630 31812 11636
rect 31392 11212 31444 11218
rect 31392 11154 31444 11160
rect 31680 11014 31708 11630
rect 31668 11008 31720 11014
rect 31668 10950 31720 10956
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31300 9580 31352 9586
rect 31300 9522 31352 9528
rect 31496 9178 31524 10610
rect 31772 10266 31800 11630
rect 31852 11008 31904 11014
rect 31852 10950 31904 10956
rect 31864 10742 31892 10950
rect 31852 10736 31904 10742
rect 31852 10678 31904 10684
rect 31864 10266 31892 10678
rect 31760 10260 31812 10266
rect 31760 10202 31812 10208
rect 31852 10260 31904 10266
rect 31852 10202 31904 10208
rect 31864 10062 31892 10202
rect 31852 10056 31904 10062
rect 31680 10004 31852 10010
rect 31680 9998 31904 10004
rect 31680 9982 31892 9998
rect 31484 9172 31536 9178
rect 31484 9114 31536 9120
rect 31680 9042 31708 9982
rect 32048 9654 32076 13874
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 32416 13530 32444 13806
rect 32404 13524 32456 13530
rect 32404 13466 32456 13472
rect 32128 13252 32180 13258
rect 32128 13194 32180 13200
rect 32140 12918 32168 13194
rect 32416 12918 32444 13466
rect 32128 12912 32180 12918
rect 32128 12854 32180 12860
rect 32404 12912 32456 12918
rect 32404 12854 32456 12860
rect 32600 12850 32628 14010
rect 32876 14006 32904 14894
rect 33324 14340 33376 14346
rect 33324 14282 33376 14288
rect 32772 14000 32824 14006
rect 32772 13942 32824 13948
rect 32864 14000 32916 14006
rect 32864 13942 32916 13948
rect 32588 12844 32640 12850
rect 32588 12786 32640 12792
rect 32784 12442 32812 13942
rect 33336 13274 33364 14282
rect 33428 13938 33456 15438
rect 33520 14618 33548 15506
rect 33612 15094 33640 17326
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 34072 16182 34100 17274
rect 34244 17128 34296 17134
rect 34244 17070 34296 17076
rect 34256 16250 34284 17070
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 36452 16652 36504 16658
rect 36452 16594 36504 16600
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 34244 16244 34296 16250
rect 34244 16186 34296 16192
rect 34060 16176 34112 16182
rect 34060 16118 34112 16124
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34520 15360 34572 15366
rect 34520 15302 34572 15308
rect 33600 15088 33652 15094
rect 33600 15030 33652 15036
rect 33612 14958 33640 15030
rect 33600 14952 33652 14958
rect 33600 14894 33652 14900
rect 34428 14952 34480 14958
rect 34428 14894 34480 14900
rect 33508 14612 33560 14618
rect 33508 14554 33560 14560
rect 33520 13954 33548 14554
rect 33612 14346 33640 14894
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34348 14346 34376 14758
rect 33600 14340 33652 14346
rect 33600 14282 33652 14288
rect 34336 14340 34388 14346
rect 34336 14282 34388 14288
rect 33520 13938 33640 13954
rect 34348 13938 34376 14282
rect 33416 13932 33468 13938
rect 33520 13932 33652 13938
rect 33520 13926 33600 13932
rect 33416 13874 33468 13880
rect 33600 13874 33652 13880
rect 34336 13932 34388 13938
rect 34336 13874 34388 13880
rect 33876 13728 33928 13734
rect 33876 13670 33928 13676
rect 33336 13258 33824 13274
rect 33888 13258 33916 13670
rect 34440 13394 34468 14894
rect 34532 14414 34560 15302
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 34612 15156 34664 15162
rect 34612 15098 34664 15104
rect 34520 14408 34572 14414
rect 34520 14350 34572 14356
rect 34428 13388 34480 13394
rect 34428 13330 34480 13336
rect 34624 13258 34652 15098
rect 34704 14952 34756 14958
rect 34704 14894 34756 14900
rect 34716 14482 34744 14894
rect 35440 14816 35492 14822
rect 35440 14758 35492 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35452 14482 35480 14758
rect 34704 14476 34756 14482
rect 34704 14418 34756 14424
rect 35440 14476 35492 14482
rect 35440 14418 35492 14424
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35348 13388 35400 13394
rect 35348 13330 35400 13336
rect 33324 13252 33824 13258
rect 33376 13246 33824 13252
rect 33324 13194 33376 13200
rect 33612 13190 33640 13246
rect 33600 13184 33652 13190
rect 33600 13126 33652 13132
rect 33692 13184 33744 13190
rect 33692 13126 33744 13132
rect 33048 12776 33100 12782
rect 33048 12718 33100 12724
rect 32772 12436 32824 12442
rect 32772 12378 32824 12384
rect 32128 11756 32180 11762
rect 32128 11698 32180 11704
rect 32140 11354 32168 11698
rect 32128 11348 32180 11354
rect 32128 11290 32180 11296
rect 32140 10062 32168 11290
rect 33060 11218 33088 12718
rect 33612 12170 33640 13126
rect 33704 12918 33732 13126
rect 33796 12918 33824 13246
rect 33876 13252 33928 13258
rect 33876 13194 33928 13200
rect 34612 13252 34664 13258
rect 34612 13194 34664 13200
rect 34612 12980 34664 12986
rect 34612 12922 34664 12928
rect 33692 12912 33744 12918
rect 33692 12854 33744 12860
rect 33784 12912 33836 12918
rect 33784 12854 33836 12860
rect 34624 12238 34652 12922
rect 35360 12646 35388 13330
rect 35452 13190 35480 14418
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 35440 13184 35492 13190
rect 35440 13126 35492 13132
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 35348 12640 35400 12646
rect 35348 12582 35400 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12238 35388 12582
rect 34520 12232 34572 12238
rect 34520 12174 34572 12180
rect 34612 12232 34664 12238
rect 34612 12174 34664 12180
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 33600 12164 33652 12170
rect 33600 12106 33652 12112
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 32692 10674 32720 11154
rect 33612 11014 33640 12106
rect 33968 11144 34020 11150
rect 33968 11086 34020 11092
rect 33600 11008 33652 11014
rect 33600 10950 33652 10956
rect 33612 10742 33640 10950
rect 33600 10736 33652 10742
rect 33600 10678 33652 10684
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 32680 10668 32732 10674
rect 32680 10610 32732 10616
rect 32404 10532 32456 10538
rect 32404 10474 32456 10480
rect 32416 10198 32444 10474
rect 32508 10266 32536 10610
rect 32496 10260 32548 10266
rect 32496 10202 32548 10208
rect 32404 10192 32456 10198
rect 32404 10134 32456 10140
rect 32508 10062 32536 10202
rect 32692 10062 32720 10610
rect 33416 10600 33468 10606
rect 33416 10542 33468 10548
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 32036 9648 32088 9654
rect 32036 9590 32088 9596
rect 31392 9036 31444 9042
rect 31392 8978 31444 8984
rect 31668 9036 31720 9042
rect 31668 8978 31720 8984
rect 31208 8968 31260 8974
rect 31208 8910 31260 8916
rect 30944 8622 31064 8650
rect 30840 8424 30892 8430
rect 30840 8366 30892 8372
rect 30656 7948 30708 7954
rect 30656 7890 30708 7896
rect 30564 7812 30616 7818
rect 30564 7754 30616 7760
rect 30576 7410 30604 7754
rect 31036 7478 31064 8622
rect 31220 8566 31248 8910
rect 31300 8900 31352 8906
rect 31300 8842 31352 8848
rect 31208 8560 31260 8566
rect 31208 8502 31260 8508
rect 31312 8362 31340 8842
rect 31404 8362 31432 8978
rect 32140 8974 32168 9998
rect 32312 9988 32364 9994
rect 32312 9930 32364 9936
rect 32324 9654 32352 9930
rect 32508 9722 32536 9998
rect 32692 9722 32720 9998
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 33428 9654 33456 10542
rect 32312 9648 32364 9654
rect 32312 9590 32364 9596
rect 33416 9648 33468 9654
rect 33416 9590 33468 9596
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 31576 8832 31628 8838
rect 31628 8792 31708 8820
rect 31576 8774 31628 8780
rect 31680 8566 31708 8792
rect 32692 8566 32720 9522
rect 32784 9178 32812 9522
rect 33048 9444 33100 9450
rect 33048 9386 33100 9392
rect 32772 9172 32824 9178
rect 32772 9114 32824 9120
rect 31668 8560 31720 8566
rect 31668 8502 31720 8508
rect 32680 8560 32732 8566
rect 32680 8502 32732 8508
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 32128 8424 32180 8430
rect 32128 8366 32180 8372
rect 31300 8356 31352 8362
rect 31300 8298 31352 8304
rect 31392 8356 31444 8362
rect 31392 8298 31444 8304
rect 31852 7880 31904 7886
rect 31852 7822 31904 7828
rect 31864 7478 31892 7822
rect 31024 7472 31076 7478
rect 31024 7414 31076 7420
rect 31852 7472 31904 7478
rect 31852 7414 31904 7420
rect 32140 7410 32168 8366
rect 32508 8294 32536 8434
rect 33060 8362 33088 9386
rect 33140 9376 33192 9382
rect 33140 9318 33192 9324
rect 33152 9042 33180 9318
rect 33428 9042 33456 9590
rect 33140 9036 33192 9042
rect 33140 8978 33192 8984
rect 33416 9036 33468 9042
rect 33468 8996 33548 9024
rect 33416 8978 33468 8984
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33428 8498 33456 8774
rect 33520 8498 33548 8996
rect 33612 8906 33640 10678
rect 33980 10470 34008 11086
rect 34244 11008 34296 11014
rect 34244 10950 34296 10956
rect 34428 11008 34480 11014
rect 34428 10950 34480 10956
rect 34256 10742 34284 10950
rect 34440 10810 34468 10950
rect 34428 10804 34480 10810
rect 34428 10746 34480 10752
rect 34244 10736 34296 10742
rect 34244 10678 34296 10684
rect 34532 10606 34560 12174
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34704 11280 34756 11286
rect 34704 11222 34756 11228
rect 34520 10600 34572 10606
rect 34520 10542 34572 10548
rect 33968 10464 34020 10470
rect 33968 10406 34020 10412
rect 34428 10464 34480 10470
rect 34428 10406 34480 10412
rect 33692 10260 33744 10266
rect 33692 10202 33744 10208
rect 33704 9586 33732 10202
rect 34440 10130 34468 10406
rect 34612 10260 34664 10266
rect 34612 10202 34664 10208
rect 34428 10124 34480 10130
rect 34428 10066 34480 10072
rect 34624 9994 34652 10202
rect 34716 10062 34744 11222
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 34796 10600 34848 10606
rect 34796 10542 34848 10548
rect 34808 10266 34836 10542
rect 35348 10464 35400 10470
rect 35348 10406 35400 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 10260 34848 10266
rect 34796 10202 34848 10208
rect 34704 10056 34756 10062
rect 34704 9998 34756 10004
rect 34796 10056 34848 10062
rect 34796 9998 34848 10004
rect 34612 9988 34664 9994
rect 34612 9930 34664 9936
rect 33784 9920 33836 9926
rect 33784 9862 33836 9868
rect 34060 9920 34112 9926
rect 34060 9862 34112 9868
rect 34244 9920 34296 9926
rect 34244 9862 34296 9868
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 33796 9450 33824 9862
rect 33784 9444 33836 9450
rect 33784 9386 33836 9392
rect 34072 9382 34100 9862
rect 34256 9586 34284 9862
rect 34624 9654 34652 9930
rect 34612 9648 34664 9654
rect 34612 9590 34664 9596
rect 34244 9580 34296 9586
rect 34244 9522 34296 9528
rect 34060 9376 34112 9382
rect 34060 9318 34112 9324
rect 34244 9376 34296 9382
rect 34244 9318 34296 9324
rect 34256 9178 34284 9318
rect 34244 9172 34296 9178
rect 34244 9114 34296 9120
rect 34624 9042 34652 9590
rect 34716 9382 34744 9998
rect 34808 9518 34836 9998
rect 35360 9586 35388 10406
rect 35452 10266 35480 11154
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 35440 10260 35492 10266
rect 35440 10202 35492 10208
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 35348 9580 35400 9586
rect 35348 9522 35400 9528
rect 34796 9512 34848 9518
rect 34796 9454 34848 9460
rect 34704 9376 34756 9382
rect 34704 9318 34756 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34612 9036 34664 9042
rect 34612 8978 34664 8984
rect 34060 8968 34112 8974
rect 34060 8910 34112 8916
rect 33600 8900 33652 8906
rect 33652 8860 33732 8888
rect 33600 8842 33652 8848
rect 33704 8634 33732 8860
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 33416 8492 33468 8498
rect 33416 8434 33468 8440
rect 33508 8492 33560 8498
rect 33508 8434 33560 8440
rect 33048 8356 33100 8362
rect 33048 8298 33100 8304
rect 32496 8288 32548 8294
rect 33428 8242 33456 8434
rect 33704 8294 33732 8570
rect 32496 8230 32548 8236
rect 33244 8214 33456 8242
rect 33692 8288 33744 8294
rect 33692 8230 33744 8236
rect 32956 7812 33008 7818
rect 32956 7754 33008 7760
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 30564 7404 30616 7410
rect 30564 7346 30616 7352
rect 32128 7404 32180 7410
rect 32128 7346 32180 7352
rect 30208 7126 30328 7154
rect 30300 6934 30328 7126
rect 30288 6928 30340 6934
rect 30576 6914 30604 7346
rect 31760 7336 31812 7342
rect 31760 7278 31812 7284
rect 30288 6870 30340 6876
rect 30392 6886 30604 6914
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 29920 6112 29972 6118
rect 29920 6054 29972 6060
rect 29828 5636 29880 5642
rect 29828 5578 29880 5584
rect 29932 5302 29960 6054
rect 30024 5370 30052 6802
rect 30104 6248 30156 6254
rect 30104 6190 30156 6196
rect 30116 5370 30144 6190
rect 30300 5778 30328 6870
rect 30392 6730 30420 6886
rect 31772 6866 31800 7278
rect 32140 6866 32168 7346
rect 32496 7200 32548 7206
rect 32496 7142 32548 7148
rect 30656 6860 30708 6866
rect 30576 6820 30656 6848
rect 30576 6730 30604 6820
rect 30656 6802 30708 6808
rect 31760 6860 31812 6866
rect 31760 6802 31812 6808
rect 32128 6860 32180 6866
rect 32128 6802 32180 6808
rect 30380 6724 30432 6730
rect 30380 6666 30432 6672
rect 30564 6724 30616 6730
rect 30564 6666 30616 6672
rect 30380 6384 30432 6390
rect 30380 6326 30432 6332
rect 30288 5772 30340 5778
rect 30208 5732 30288 5760
rect 30012 5364 30064 5370
rect 30012 5306 30064 5312
rect 30104 5364 30156 5370
rect 30104 5306 30156 5312
rect 29736 5296 29788 5302
rect 29736 5238 29788 5244
rect 29920 5296 29972 5302
rect 29920 5238 29972 5244
rect 30208 5234 30236 5732
rect 30288 5714 30340 5720
rect 30392 5658 30420 6326
rect 30472 6248 30524 6254
rect 30472 6190 30524 6196
rect 30484 5914 30512 6190
rect 32140 6118 32168 6802
rect 32220 6792 32272 6798
rect 32220 6734 32272 6740
rect 32232 6322 32260 6734
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 32128 6112 32180 6118
rect 32128 6054 32180 6060
rect 32312 6112 32364 6118
rect 32312 6054 32364 6060
rect 30472 5908 30524 5914
rect 30472 5850 30524 5856
rect 32324 5778 32352 6054
rect 32312 5772 32364 5778
rect 32312 5714 32364 5720
rect 30300 5630 30420 5658
rect 31116 5704 31168 5710
rect 31116 5646 31168 5652
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 30196 5228 30248 5234
rect 30196 5170 30248 5176
rect 29460 4548 29512 4554
rect 29460 4490 29512 4496
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 29472 4078 29500 4490
rect 30300 4214 30328 5630
rect 30380 5296 30432 5302
rect 30380 5238 30432 5244
rect 30392 4758 30420 5238
rect 31128 5234 31156 5646
rect 32324 5370 32352 5714
rect 32312 5364 32364 5370
rect 32312 5306 32364 5312
rect 32508 5302 32536 7142
rect 32968 6848 32996 7754
rect 33048 6860 33100 6866
rect 32968 6820 33048 6848
rect 33048 6802 33100 6808
rect 32588 6724 32640 6730
rect 32588 6666 32640 6672
rect 32600 6390 32628 6666
rect 32588 6384 32640 6390
rect 32588 6326 32640 6332
rect 33060 6254 33088 6802
rect 32680 6248 32732 6254
rect 32680 6190 32732 6196
rect 33048 6248 33100 6254
rect 33048 6190 33100 6196
rect 32496 5296 32548 5302
rect 32496 5238 32548 5244
rect 30840 5228 30892 5234
rect 30840 5170 30892 5176
rect 31024 5228 31076 5234
rect 31024 5170 31076 5176
rect 31116 5228 31168 5234
rect 31116 5170 31168 5176
rect 30472 5092 30524 5098
rect 30472 5034 30524 5040
rect 30380 4752 30432 4758
rect 30380 4694 30432 4700
rect 30484 4622 30512 5034
rect 30656 5024 30708 5030
rect 30656 4966 30708 4972
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30380 4480 30432 4486
rect 30380 4422 30432 4428
rect 30392 4282 30420 4422
rect 30380 4276 30432 4282
rect 30380 4218 30432 4224
rect 30288 4208 30340 4214
rect 30288 4150 30340 4156
rect 29460 4072 29512 4078
rect 29460 4014 29512 4020
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30012 3528 30064 3534
rect 30012 3470 30064 3476
rect 30024 2990 30052 3470
rect 30484 3126 30512 3878
rect 30668 3602 30696 4966
rect 30852 4690 30880 5170
rect 30840 4684 30892 4690
rect 30840 4626 30892 4632
rect 31036 4554 31064 5170
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 32324 4758 32352 4966
rect 32312 4752 32364 4758
rect 32312 4694 32364 4700
rect 31944 4684 31996 4690
rect 31944 4626 31996 4632
rect 31024 4548 31076 4554
rect 31024 4490 31076 4496
rect 31300 4480 31352 4486
rect 31300 4422 31352 4428
rect 31312 4214 31340 4422
rect 31956 4282 31984 4626
rect 32036 4616 32088 4622
rect 32036 4558 32088 4564
rect 31760 4276 31812 4282
rect 31760 4218 31812 4224
rect 31944 4276 31996 4282
rect 31944 4218 31996 4224
rect 31300 4208 31352 4214
rect 31300 4150 31352 4156
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 30760 3754 30788 4082
rect 30760 3726 30972 3754
rect 31772 3738 31800 4218
rect 32048 4214 32076 4558
rect 32312 4480 32364 4486
rect 32312 4422 32364 4428
rect 32496 4480 32548 4486
rect 32496 4422 32548 4428
rect 32324 4282 32352 4422
rect 32312 4276 32364 4282
rect 32312 4218 32364 4224
rect 32404 4276 32456 4282
rect 32404 4218 32456 4224
rect 32036 4208 32088 4214
rect 32036 4150 32088 4156
rect 31852 4072 31904 4078
rect 31852 4014 31904 4020
rect 30656 3596 30708 3602
rect 30656 3538 30708 3544
rect 30944 3466 30972 3726
rect 31760 3732 31812 3738
rect 31760 3674 31812 3680
rect 31864 3602 31892 4014
rect 31852 3596 31904 3602
rect 31852 3538 31904 3544
rect 30932 3460 30984 3466
rect 30932 3402 30984 3408
rect 30944 3126 30972 3402
rect 30472 3120 30524 3126
rect 30472 3062 30524 3068
rect 30932 3120 30984 3126
rect 30932 3062 30984 3068
rect 32048 2990 32076 4150
rect 32416 4078 32444 4218
rect 32508 4146 32536 4422
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 32692 4078 32720 6190
rect 33060 4078 33088 6190
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 33152 5234 33180 5714
rect 33244 5710 33272 8214
rect 33324 7812 33376 7818
rect 33324 7754 33376 7760
rect 33336 6662 33364 7754
rect 33704 7478 33732 8230
rect 34072 7886 34100 8910
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 34256 8566 34284 8774
rect 34244 8560 34296 8566
rect 34244 8502 34296 8508
rect 34624 8090 34652 8978
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34980 8968 35032 8974
rect 34980 8910 35032 8916
rect 34612 8084 34664 8090
rect 34612 8026 34664 8032
rect 34060 7880 34112 7886
rect 34060 7822 34112 7828
rect 34072 7478 34100 7822
rect 34336 7744 34388 7750
rect 34336 7686 34388 7692
rect 33692 7472 33744 7478
rect 33692 7414 33744 7420
rect 34060 7472 34112 7478
rect 34060 7414 34112 7420
rect 33704 6798 33732 7414
rect 34348 7410 34376 7686
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 34520 7268 34572 7274
rect 34520 7210 34572 7216
rect 34152 6928 34204 6934
rect 34152 6870 34204 6876
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33600 6384 33652 6390
rect 33600 6326 33652 6332
rect 33612 5914 33640 6326
rect 33704 6202 33732 6734
rect 34060 6724 34112 6730
rect 34060 6666 34112 6672
rect 33784 6384 33836 6390
rect 34072 6338 34100 6666
rect 34164 6390 34192 6870
rect 34336 6792 34388 6798
rect 34336 6734 34388 6740
rect 34348 6390 34376 6734
rect 33836 6332 34100 6338
rect 33784 6326 34100 6332
rect 34152 6384 34204 6390
rect 34152 6326 34204 6332
rect 34336 6384 34388 6390
rect 34336 6326 34388 6332
rect 33796 6310 34100 6326
rect 33704 6174 34008 6202
rect 33692 6112 33744 6118
rect 33692 6054 33744 6060
rect 33784 6112 33836 6118
rect 33784 6054 33836 6060
rect 33704 5914 33732 6054
rect 33600 5908 33652 5914
rect 33600 5850 33652 5856
rect 33692 5908 33744 5914
rect 33692 5850 33744 5856
rect 33704 5760 33732 5850
rect 33796 5846 33824 6054
rect 33784 5840 33836 5846
rect 33784 5782 33836 5788
rect 33612 5732 33732 5760
rect 33232 5704 33284 5710
rect 33232 5646 33284 5652
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 33140 5228 33192 5234
rect 33140 5170 33192 5176
rect 33244 5030 33272 5646
rect 33324 5636 33376 5642
rect 33324 5578 33376 5584
rect 33336 5302 33364 5578
rect 33324 5296 33376 5302
rect 33324 5238 33376 5244
rect 33428 5234 33456 5646
rect 33416 5228 33468 5234
rect 33416 5170 33468 5176
rect 33232 5024 33284 5030
rect 33232 4966 33284 4972
rect 33244 4706 33272 4966
rect 33152 4678 33272 4706
rect 33152 4622 33180 4678
rect 33140 4616 33192 4622
rect 33140 4558 33192 4564
rect 33232 4616 33284 4622
rect 33232 4558 33284 4564
rect 33324 4616 33376 4622
rect 33324 4558 33376 4564
rect 32404 4072 32456 4078
rect 32404 4014 32456 4020
rect 32680 4072 32732 4078
rect 32680 4014 32732 4020
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 32956 3732 33008 3738
rect 32956 3674 33008 3680
rect 32968 3534 32996 3674
rect 32956 3528 33008 3534
rect 32956 3470 33008 3476
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 32416 3126 32444 3334
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 33060 2990 33088 4014
rect 33244 3602 33272 4558
rect 33336 4282 33364 4558
rect 33428 4554 33456 5170
rect 33416 4548 33468 4554
rect 33416 4490 33468 4496
rect 33428 4282 33456 4490
rect 33324 4276 33376 4282
rect 33324 4218 33376 4224
rect 33416 4276 33468 4282
rect 33416 4218 33468 4224
rect 33612 3942 33640 5732
rect 33784 5704 33836 5710
rect 33784 5646 33836 5652
rect 33692 4616 33744 4622
rect 33692 4558 33744 4564
rect 33704 4214 33732 4558
rect 33692 4208 33744 4214
rect 33692 4150 33744 4156
rect 33600 3936 33652 3942
rect 33600 3878 33652 3884
rect 33612 3670 33640 3878
rect 33600 3664 33652 3670
rect 33600 3606 33652 3612
rect 33232 3596 33284 3602
rect 33232 3538 33284 3544
rect 33796 3482 33824 5646
rect 33980 4146 34008 6174
rect 34072 5166 34100 6310
rect 34532 5642 34560 7210
rect 34624 6662 34652 8026
rect 34808 6662 34836 8910
rect 34992 8634 35020 8910
rect 36464 8906 36492 16594
rect 36636 16516 36688 16522
rect 36636 16458 36688 16464
rect 36648 16425 36676 16458
rect 36634 16416 36690 16425
rect 36634 16351 36690 16360
rect 35992 8900 36044 8906
rect 35992 8842 36044 8848
rect 36452 8900 36504 8906
rect 36452 8842 36504 8848
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 36004 7954 36032 8842
rect 35992 7948 36044 7954
rect 35992 7890 36044 7896
rect 35440 7880 35492 7886
rect 35440 7822 35492 7828
rect 35452 7478 35480 7822
rect 36176 7812 36228 7818
rect 36176 7754 36228 7760
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 35440 7472 35492 7478
rect 35440 7414 35492 7420
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34612 6656 34664 6662
rect 34612 6598 34664 6604
rect 34796 6656 34848 6662
rect 34796 6598 34848 6604
rect 34624 5914 34652 6598
rect 34808 6254 34836 6598
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34796 6248 34848 6254
rect 34796 6190 34848 6196
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 35072 5636 35124 5642
rect 35072 5578 35124 5584
rect 35084 5302 35112 5578
rect 35072 5296 35124 5302
rect 35072 5238 35124 5244
rect 34704 5228 34756 5234
rect 34704 5170 34756 5176
rect 34888 5228 34940 5234
rect 34888 5170 34940 5176
rect 34060 5160 34112 5166
rect 34060 5102 34112 5108
rect 34428 5160 34480 5166
rect 34428 5102 34480 5108
rect 34336 5092 34388 5098
rect 34336 5034 34388 5040
rect 34348 4554 34376 5034
rect 34440 4690 34468 5102
rect 34716 4758 34744 5170
rect 34900 5114 34928 5170
rect 34808 5086 34928 5114
rect 34808 5030 34836 5086
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 34704 4752 34756 4758
rect 34704 4694 34756 4700
rect 34808 4706 34836 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34428 4684 34480 4690
rect 34428 4626 34480 4632
rect 34336 4548 34388 4554
rect 34336 4490 34388 4496
rect 33968 4140 34020 4146
rect 33968 4082 34020 4088
rect 33704 3466 33824 3482
rect 33692 3460 33824 3466
rect 33744 3454 33824 3460
rect 33692 3402 33744 3408
rect 33980 3126 34008 4082
rect 34716 3466 34744 4694
rect 34808 4678 34928 4706
rect 34900 4622 34928 4678
rect 35360 4622 35388 5850
rect 36188 5574 36216 7754
rect 36726 6216 36782 6225
rect 36726 6151 36728 6160
rect 36780 6151 36782 6160
rect 36728 6122 36780 6128
rect 36176 5568 36228 5574
rect 36176 5510 36228 5516
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 35532 5024 35584 5030
rect 35532 4966 35584 4972
rect 34888 4616 34940 4622
rect 34888 4558 34940 4564
rect 35348 4616 35400 4622
rect 35348 4558 35400 4564
rect 35544 4554 35572 4966
rect 35532 4548 35584 4554
rect 35532 4490 35584 4496
rect 35348 4480 35400 4486
rect 35348 4422 35400 4428
rect 35360 4214 35388 4422
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 35348 4208 35400 4214
rect 35348 4150 35400 4156
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34704 3460 34756 3466
rect 34704 3402 34756 3408
rect 34716 3194 34744 3402
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 33968 3120 34020 3126
rect 33968 3062 34020 3068
rect 30012 2984 30064 2990
rect 30012 2926 30064 2932
rect 32036 2984 32088 2990
rect 32036 2926 32088 2932
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23216 800 23244 2382
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 10322 0 10378 800
rect 23202 0 23258 800
<< via2 >>
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 846 36896 902 36952
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 1122 29280 1178 29336
rect 846 25372 848 25392
rect 848 25372 900 25392
rect 900 25372 902 25392
rect 846 25336 902 25372
rect 846 23724 902 23760
rect 846 23704 848 23724
rect 848 23704 900 23724
rect 900 23704 902 23724
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 5630 30096 5686 30152
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 5630 26732 5632 26752
rect 5632 26732 5684 26752
rect 5684 26732 5686 26752
rect 5630 26696 5686 26732
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 9126 30132 9128 30152
rect 9128 30132 9180 30152
rect 9180 30132 9182 30152
rect 9126 30096 9182 30132
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 7102 26732 7104 26752
rect 7104 26732 7156 26752
rect 7156 26732 7158 26752
rect 7102 26696 7158 26732
rect 25502 36660 25504 36680
rect 25504 36660 25556 36680
rect 25556 36660 25558 36680
rect 25502 36624 25558 36660
rect 23570 35692 23626 35728
rect 23570 35672 23572 35692
rect 23572 35672 23624 35692
rect 23624 35672 23626 35692
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 1398 17720 1454 17776
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1306 14320 1362 14376
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 24766 35536 24822 35592
rect 28814 36624 28870 36680
rect 30102 33108 30158 33144
rect 30102 33088 30104 33108
rect 30104 33088 30156 33108
rect 30156 33088 30158 33108
rect 30194 32952 30250 33008
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 32770 35672 32826 35728
rect 32770 35556 32826 35592
rect 32770 35536 32772 35556
rect 32772 35536 32824 35556
rect 32824 35536 32826 35556
rect 32678 35148 32734 35184
rect 32678 35128 32680 35148
rect 32680 35128 32732 35148
rect 32732 35128 32734 35148
rect 33322 35028 33324 35048
rect 33324 35028 33376 35048
rect 33376 35028 33378 35048
rect 33322 34992 33378 35028
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34610 35128 34666 35184
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35530 35028 35532 35048
rect 35532 35028 35584 35048
rect 35584 35028 35586 35048
rect 35530 34992 35586 35028
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34426 32952 34482 33008
rect 34610 33088 34666 33144
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 36634 16360 36690 16416
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 36726 6180 36782 6216
rect 36726 6160 36728 6180
rect 36728 6160 36780 6180
rect 36780 6160 36782 6180
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 841 36954 907 36957
rect 798 36952 907 36954
rect 798 36896 846 36952
rect 902 36896 907 36952
rect 798 36891 907 36896
rect 798 36848 858 36891
rect 0 36758 858 36848
rect 0 36728 800 36758
rect 25497 36682 25563 36685
rect 28809 36682 28875 36685
rect 25497 36680 28875 36682
rect 25497 36624 25502 36680
rect 25558 36624 28814 36680
rect 28870 36624 28875 36680
rect 25497 36622 28875 36624
rect 25497 36619 25563 36622
rect 28809 36619 28875 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 23565 35730 23631 35733
rect 32765 35730 32831 35733
rect 23565 35728 32831 35730
rect 23565 35672 23570 35728
rect 23626 35672 32770 35728
rect 32826 35672 32831 35728
rect 23565 35670 32831 35672
rect 23565 35667 23631 35670
rect 32765 35667 32831 35670
rect 24761 35594 24827 35597
rect 32765 35594 32831 35597
rect 24761 35592 32831 35594
rect 24761 35536 24766 35592
rect 24822 35536 32770 35592
rect 32826 35536 32831 35592
rect 24761 35534 32831 35536
rect 24761 35531 24827 35534
rect 32765 35531 32831 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 32673 35186 32739 35189
rect 34605 35186 34671 35189
rect 32673 35184 34671 35186
rect 32673 35128 32678 35184
rect 32734 35128 34610 35184
rect 34666 35128 34671 35184
rect 32673 35126 34671 35128
rect 32673 35123 32739 35126
rect 34605 35123 34671 35126
rect 33317 35050 33383 35053
rect 35525 35050 35591 35053
rect 33317 35048 35591 35050
rect 33317 34992 33322 35048
rect 33378 34992 35530 35048
rect 35586 34992 35591 35048
rect 33317 34990 35591 34992
rect 33317 34987 33383 34990
rect 35525 34987 35591 34990
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 30097 33146 30163 33149
rect 34605 33146 34671 33149
rect 30097 33144 34671 33146
rect 30097 33088 30102 33144
rect 30158 33088 34610 33144
rect 34666 33088 34671 33144
rect 30097 33086 34671 33088
rect 30097 33083 30163 33086
rect 34605 33083 34671 33086
rect 30189 33010 30255 33013
rect 34421 33010 34487 33013
rect 30189 33008 34487 33010
rect 30189 32952 30194 33008
rect 30250 32952 34426 33008
rect 34482 32952 34487 33008
rect 30189 32950 34487 32952
rect 30189 32947 30255 32950
rect 34421 32947 34487 32950
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 5625 30154 5691 30157
rect 9121 30154 9187 30157
rect 5625 30152 9187 30154
rect 5625 30096 5630 30152
rect 5686 30096 9126 30152
rect 9182 30096 9187 30152
rect 5625 30094 9187 30096
rect 5625 30091 5691 30094
rect 9121 30091 9187 30094
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 4870 29408 5186 29409
rect 0 29338 800 29368
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 1117 29338 1183 29341
rect 0 29336 1183 29338
rect 0 29280 1122 29336
rect 1178 29280 1183 29336
rect 0 29278 1183 29280
rect 0 29248 800 29278
rect 1117 29275 1183 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 5625 26754 5691 26757
rect 7097 26754 7163 26757
rect 5625 26752 7163 26754
rect 5625 26696 5630 26752
rect 5686 26696 7102 26752
rect 7158 26696 7163 26752
rect 5625 26694 7163 26696
rect 5625 26691 5691 26694
rect 7097 26691 7163 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 841 25394 907 25397
rect 798 25392 907 25394
rect 798 25336 846 25392
rect 902 25336 907 25392
rect 798 25331 907 25336
rect 798 25288 858 25331
rect 0 25198 858 25288
rect 0 25168 800 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 4870 23968 5186 23969
rect 0 23898 800 23928
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 0 23808 858 23898
rect 798 23765 858 23808
rect 798 23760 907 23765
rect 798 23704 846 23760
rect 902 23704 907 23760
rect 798 23702 907 23704
rect 841 23699 907 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 36629 16418 36695 16421
rect 37408 16418 38208 16448
rect 36629 16416 38208 16418
rect 36629 16360 36634 16416
rect 36690 16360 38208 16416
rect 36629 16358 38208 16360
rect 36629 16355 36695 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 37408 16328 38208 16358
rect 35590 16287 35906 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 0 14378 800 14408
rect 1301 14378 1367 14381
rect 0 14376 1367 14378
rect 0 14320 1306 14376
rect 1362 14320 1367 14376
rect 0 14318 1367 14320
rect 0 14288 800 14318
rect 1301 14315 1367 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 36721 6218 36787 6221
rect 37408 6218 38208 6248
rect 36721 6216 38208 6218
rect 36721 6160 36726 6216
rect 36782 6160 38208 6216
rect 36721 6158 38208 6160
rect 36721 6155 36787 6158
rect 37408 6128 38208 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 38128
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 38112 5188 38128
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 37568 35248 38128
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 38112 35908 38128
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 4910 6048 5146 6284
rect 34970 36024 35206 36260
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 37124 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 37124 36920
rect 1056 36642 37124 36684
rect 1056 36260 37124 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 37124 36260
rect 1056 35982 37124 36024
rect 1056 6284 37124 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 37124 6284
rect 1056 6006 37124 6048
rect 1056 5624 37124 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 37124 5624
rect 1056 5346 37124 5388
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 0
transform -1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 0
transform 1 0 9936 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 0
transform -1 0 10672 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 0
transform 1 0 35512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 0
transform -1 0 31188 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0534_
timestamp 0
transform -1 0 10948 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0535_
timestamp 0
transform 1 0 9660 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0536_
timestamp 0
transform 1 0 9568 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0537_
timestamp 0
transform -1 0 4416 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0538_
timestamp 0
transform 1 0 5704 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0539_
timestamp 0
transform 1 0 5704 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0540_
timestamp 0
transform 1 0 5336 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0541_
timestamp 0
transform 1 0 9476 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0542_
timestamp 0
transform -1 0 10396 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0543_
timestamp 0
transform 1 0 6348 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0544_
timestamp 0
transform 1 0 6164 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0545_
timestamp 0
transform 1 0 32752 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0546_
timestamp 0
transform -1 0 34868 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _0547_
timestamp 0
transform 1 0 32660 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _0548_
timestamp 0
transform 1 0 34684 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0549_
timestamp 0
transform -1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0550_
timestamp 0
transform -1 0 34500 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0551_
timestamp 0
transform 1 0 31372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0552_
timestamp 0
transform 1 0 29532 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0553_
timestamp 0
transform -1 0 29440 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _0554_
timestamp 0
transform -1 0 32016 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _0555_
timestamp 0
transform 1 0 28612 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _0556_
timestamp 0
transform -1 0 31004 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0557_
timestamp 0
transform 1 0 31372 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0558_
timestamp 0
transform -1 0 29992 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0559_
timestamp 0
transform -1 0 2392 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0560_
timestamp 0
transform 1 0 3312 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0561_
timestamp 0
transform 1 0 1840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0562_
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0563_
timestamp 0
transform 1 0 3496 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0564_
timestamp 0
transform -1 0 4784 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 0
transform 1 0 4784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0566_
timestamp 0
transform 1 0 1932 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0567_
timestamp 0
transform 1 0 2484 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0568_
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0569_
timestamp 0
transform -1 0 3496 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _0570_
timestamp 0
transform 1 0 2760 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _0571_
timestamp 0
transform -1 0 4232 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0572_
timestamp 0
transform -1 0 3128 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0573_
timestamp 0
transform -1 0 2484 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 0
transform 1 0 2024 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0575_
timestamp 0
transform -1 0 4416 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0576_
timestamp 0
transform 1 0 3864 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0577_
timestamp 0
transform -1 0 4140 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0578_
timestamp 0
transform -1 0 5060 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0579_
timestamp 0
transform 1 0 3772 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0580_
timestamp 0
transform 1 0 4416 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0581_
timestamp 0
transform 1 0 5060 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0582_
timestamp 0
transform -1 0 5888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0583_
timestamp 0
transform 1 0 5244 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0584_
timestamp 0
transform 1 0 5520 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0585_
timestamp 0
transform 1 0 6348 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0586_
timestamp 0
transform 1 0 6348 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0587_
timestamp 0
transform -1 0 6256 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0588_
timestamp 0
transform 1 0 5336 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0589_
timestamp 0
transform 1 0 5244 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 0
transform -1 0 6348 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0591_
timestamp 0
transform 1 0 5796 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0592_
timestamp 0
transform 1 0 7452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0593_
timestamp 0
transform -1 0 7452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0594_
timestamp 0
transform -1 0 7268 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0595_
timestamp 0
transform 1 0 5152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0596_
timestamp 0
transform -1 0 6808 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0597_
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 0
transform 1 0 4324 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0599_
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0600_
timestamp 0
transform -1 0 6256 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0601_
timestamp 0
transform -1 0 6808 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 0
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0603_
timestamp 0
transform 1 0 4968 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0604_
timestamp 0
transform -1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 0
transform 1 0 2300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 0
transform -1 0 2116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0607_
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0608_
timestamp 0
transform -1 0 5796 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0609_
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0610_
timestamp 0
transform 1 0 4324 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0611_
timestamp 0
transform -1 0 6992 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0612_
timestamp 0
transform -1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0613_
timestamp 0
transform 1 0 5796 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0614_
timestamp 0
transform -1 0 7544 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0615_
timestamp 0
transform 1 0 7268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0616_
timestamp 0
transform 1 0 5888 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0617_
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 0
transform 1 0 6440 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0619_
timestamp 0
transform 1 0 7728 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _0620_
timestamp 0
transform 1 0 7636 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0621_
timestamp 0
transform 1 0 6900 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0622_
timestamp 0
transform -1 0 8832 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 0
transform 1 0 9016 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 0
transform 1 0 8188 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _0625_
timestamp 0
transform -1 0 9660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0626_
timestamp 0
transform 1 0 8832 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0627_
timestamp 0
transform 1 0 9016 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0628_
timestamp 0
transform -1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0629_
timestamp 0
transform 1 0 9752 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 0
transform 1 0 10120 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0631_
timestamp 0
transform -1 0 10212 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0632_
timestamp 0
transform 1 0 10304 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0633_
timestamp 0
transform 1 0 10212 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0634_
timestamp 0
transform 1 0 10672 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0635_
timestamp 0
transform -1 0 9568 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0636_
timestamp 0
transform 1 0 9476 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0637_
timestamp 0
transform 1 0 9752 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0638_
timestamp 0
transform 1 0 8188 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 0
transform 1 0 8188 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0640_
timestamp 0
transform 1 0 9108 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0641_
timestamp 0
transform 1 0 7360 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0642_
timestamp 0
transform -1 0 9660 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0643_
timestamp 0
transform -1 0 9292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0644_
timestamp 0
transform 1 0 9752 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0645_
timestamp 0
transform -1 0 11408 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0646_
timestamp 0
transform -1 0 10212 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0647_
timestamp 0
transform 1 0 10396 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0648_
timestamp 0
transform 1 0 9200 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0649_
timestamp 0
transform 1 0 9936 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0650_
timestamp 0
transform 1 0 10856 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0651_
timestamp 0
transform -1 0 11040 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0652_
timestamp 0
transform -1 0 10856 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0653_
timestamp 0
transform 1 0 8188 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0654_
timestamp 0
transform 1 0 9476 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0655_
timestamp 0
transform -1 0 8740 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0656_
timestamp 0
transform 1 0 8004 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0657_
timestamp 0
transform 1 0 7912 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0658_
timestamp 0
transform 1 0 7728 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0659_
timestamp 0
transform -1 0 9016 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0660_
timestamp 0
transform -1 0 8372 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 0
transform 1 0 9752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0662_
timestamp 0
transform 1 0 9016 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0663_
timestamp 0
transform 1 0 8924 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0664_
timestamp 0
transform 1 0 10672 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0665_
timestamp 0
transform 1 0 10028 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0666_
timestamp 0
transform 1 0 30176 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0667_
timestamp 0
transform 1 0 29992 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _0668_
timestamp 0
transform 1 0 34684 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__and3_1  _0669_
timestamp 0
transform -1 0 32568 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0670_
timestamp 0
transform -1 0 30544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0671_
timestamp 0
transform 1 0 30636 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0672_
timestamp 0
transform -1 0 31648 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _0673_
timestamp 0
transform -1 0 30728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_1  _0674_
timestamp 0
transform 1 0 31924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0675_
timestamp 0
transform -1 0 32660 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0676_
timestamp 0
transform -1 0 31372 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0677_
timestamp 0
transform -1 0 34040 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _0678_
timestamp 0
transform -1 0 33764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 0
transform -1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0680_
timestamp 0
transform 1 0 34868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0681_
timestamp 0
transform -1 0 35328 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0682_
timestamp 0
transform -1 0 35788 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0683_
timestamp 0
transform -1 0 33672 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0684_
timestamp 0
transform 1 0 33488 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0685_
timestamp 0
transform -1 0 34592 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0686_
timestamp 0
transform -1 0 33396 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 0
transform 1 0 29532 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0688_
timestamp 0
transform 1 0 33120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0689_
timestamp 0
transform 1 0 28980 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _0690_
timestamp 0
transform -1 0 30360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0691_
timestamp 0
transform -1 0 31832 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0692_
timestamp 0
transform 1 0 30636 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0693_
timestamp 0
transform 1 0 29900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0694_
timestamp 0
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0695_
timestamp 0
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0696_
timestamp 0
transform 1 0 30268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _0697_
timestamp 0
transform 1 0 31740 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0698_
timestamp 0
transform 1 0 31280 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 0
transform -1 0 31280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0700_
timestamp 0
transform 1 0 33672 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 0
transform -1 0 31740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0702_
timestamp 0
transform -1 0 32016 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0703_
timestamp 0
transform -1 0 34684 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0704_
timestamp 0
transform 1 0 34684 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0705_
timestamp 0
transform -1 0 34224 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _0706_
timestamp 0
transform 1 0 34684 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0707_
timestamp 0
transform -1 0 35604 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _0708_
timestamp 0
transform -1 0 34316 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 0
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0710_
timestamp 0
transform 1 0 27140 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 0
transform 1 0 27508 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0713_
timestamp 0
transform 1 0 28520 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 0
transform 1 0 28796 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 0
transform -1 0 26864 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0717_
timestamp 0
transform 1 0 26128 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0718_
timestamp 0
transform 1 0 27968 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0719_
timestamp 0
transform 1 0 29256 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0720_
timestamp 0
transform 1 0 30360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0721_
timestamp 0
transform -1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0722_
timestamp 0
transform -1 0 32936 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0723_
timestamp 0
transform -1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0724_
timestamp 0
transform 1 0 34684 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0725_
timestamp 0
transform -1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0726_
timestamp 0
transform -1 0 34132 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0727_
timestamp 0
transform 1 0 32476 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0728_
timestamp 0
transform -1 0 32476 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0729_
timestamp 0
transform 1 0 32108 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0730_
timestamp 0
transform 1 0 28612 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0731_
timestamp 0
transform 1 0 29164 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 0
transform 1 0 27600 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0733_
timestamp 0
transform 1 0 26956 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0734_
timestamp 0
transform 1 0 25392 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0735_
timestamp 0
transform -1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 0
transform 1 0 25024 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0737_
timestamp 0
transform 1 0 23460 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 0
transform 1 0 24656 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0739_
timestamp 0
transform 1 0 24748 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 0
transform 1 0 25484 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0741_
timestamp 0
transform -1 0 26036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0742_
timestamp 0
transform -1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0743_
timestamp 0
transform 1 0 23368 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 0
transform 1 0 23368 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0745_
timestamp 0
transform 1 0 22908 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0746_
timestamp 0
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0747_
timestamp 0
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 0
transform 1 0 22540 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0749_
timestamp 0
transform -1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0750_
timestamp 0
transform -1 0 21804 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0751_
timestamp 0
transform 1 0 20240 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0752_
timestamp 0
transform 1 0 22816 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0753_
timestamp 0
transform 1 0 21344 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0754_
timestamp 0
transform -1 0 21344 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0755_
timestamp 0
transform -1 0 21252 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 0
transform 1 0 20700 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0757_
timestamp 0
transform -1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0758_
timestamp 0
transform -1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0759_
timestamp 0
transform 1 0 23276 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 0
transform 1 0 23368 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0761_
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0762_
timestamp 0
transform -1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0763_
timestamp 0
transform -1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 0
transform 1 0 25760 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0765_
timestamp 0
transform -1 0 28796 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 0
transform 1 0 28152 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0767_
timestamp 0
transform 1 0 30268 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 0
transform 1 0 31096 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 0
transform 1 0 32292 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0770_
timestamp 0
transform -1 0 34408 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0771_
timestamp 0
transform 1 0 34132 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0772_
timestamp 0
transform -1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0773_
timestamp 0
transform -1 0 35512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0774_
timestamp 0
transform 1 0 33212 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp 0
transform -1 0 34040 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0776_
timestamp 0
transform 1 0 31372 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0777_
timestamp 0
transform 1 0 30912 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 0
transform 1 0 31188 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0779_
timestamp 0
transform -1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0780_
timestamp 0
transform -1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0781_
timestamp 0
transform 1 0 28244 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0782_
timestamp 0
transform 1 0 26680 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0783_
timestamp 0
transform 1 0 25576 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0784_
timestamp 0
transform -1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0785_
timestamp 0
transform -1 0 23736 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 0
transform 1 0 22908 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0787_
timestamp 0
transform -1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0788_
timestamp 0
transform -1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0789_
timestamp 0
transform -1 0 20700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0790_
timestamp 0
transform -1 0 20424 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0791_
timestamp 0
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 0
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0793_
timestamp 0
transform 1 0 18124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0794_
timestamp 0
transform -1 0 19596 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0795_
timestamp 0
transform -1 0 18400 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0796_
timestamp 0
transform -1 0 18032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0797_
timestamp 0
transform -1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0798_
timestamp 0
transform -1 0 15456 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0799_
timestamp 0
transform -1 0 16008 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0800_
timestamp 0
transform -1 0 16100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0801_
timestamp 0
transform -1 0 15824 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0802_
timestamp 0
transform -1 0 15824 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 0
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 0
transform 1 0 15732 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0805_
timestamp 0
transform -1 0 16192 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0806_
timestamp 0
transform -1 0 16192 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0807_
timestamp 0
transform -1 0 16100 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0808_
timestamp 0
transform -1 0 15824 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 0
transform 1 0 15916 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0810_
timestamp 0
transform -1 0 16376 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 0
transform 1 0 16100 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0812_
timestamp 0
transform -1 0 16100 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 0
transform 1 0 15640 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0814_
timestamp 0
transform -1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0815_
timestamp 0
transform -1 0 18584 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0816_
timestamp 0
transform 1 0 17756 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0817_
timestamp 0
transform 1 0 17940 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 0
transform 1 0 18676 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0819_
timestamp 0
transform -1 0 18860 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0820_
timestamp 0
transform 1 0 17756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 0
transform 1 0 17572 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0822_
timestamp 0
transform -1 0 19504 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0823_
timestamp 0
transform -1 0 18584 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0824_
timestamp 0
transform 1 0 17204 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0825_
timestamp 0
transform 1 0 17112 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0826_
timestamp 0
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0827_
timestamp 0
transform -1 0 18952 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0828_
timestamp 0
transform 1 0 20148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 0
transform 1 0 22172 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0830_
timestamp 0
transform 1 0 20148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0831_
timestamp 0
transform -1 0 22172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0832_
timestamp 0
transform -1 0 21896 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0834_
timestamp 0
transform -1 0 24288 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0835_
timestamp 0
transform -1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0836_
timestamp 0
transform -1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0837_
timestamp 0
transform -1 0 29164 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _0838_
timestamp 0
transform -1 0 32660 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _0839_
timestamp 0
transform -1 0 32016 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__and3_1  _0840_
timestamp 0
transform -1 0 27508 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0841_
timestamp 0
transform 1 0 26956 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0842_
timestamp 0
transform 1 0 28060 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _0843_
timestamp 0
transform -1 0 27600 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _0844_
timestamp 0
transform -1 0 28612 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_1  _0845_
timestamp 0
transform 1 0 27968 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0846_
timestamp 0
transform -1 0 29440 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0847_
timestamp 0
transform -1 0 28980 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0848_
timestamp 0
transform 1 0 29348 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _0849_
timestamp 0
transform -1 0 29348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 0
transform -1 0 28244 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0851_
timestamp 0
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0852_
timestamp 0
transform 1 0 31464 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0853_
timestamp 0
transform -1 0 29808 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0854_
timestamp 0
transform 1 0 30268 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0855_
timestamp 0
transform 1 0 27508 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0856_
timestamp 0
transform -1 0 30452 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0857_
timestamp 0
transform -1 0 30176 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _0858_
timestamp 0
transform -1 0 31372 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_2  _0859_
timestamp 0
transform 1 0 32016 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0860_
timestamp 0
transform 1 0 32108 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0861_
timestamp 0
transform -1 0 31832 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0862_
timestamp 0
transform 1 0 32108 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0863_
timestamp 0
transform 1 0 32568 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0864_
timestamp 0
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 0
transform -1 0 33580 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0866_
timestamp 0
transform -1 0 35880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0867_
timestamp 0
transform -1 0 33672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _0868_
timestamp 0
transform -1 0 33856 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0869_
timestamp 0
transform 1 0 33764 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 0
transform 1 0 33672 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0871_
timestamp 0
transform 1 0 33028 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 0
transform -1 0 30268 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0873_
timestamp 0
transform -1 0 33028 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0874_
timestamp 0
transform -1 0 34868 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 0
transform -1 0 35972 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0876_
timestamp 0
transform -1 0 34408 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 0
transform -1 0 35328 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0878_
timestamp 0
transform -1 0 35236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _0879_
timestamp 0
transform -1 0 34960 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 0
transform -1 0 32016 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0881_
timestamp 0
transform -1 0 35052 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0882_
timestamp 0
transform 1 0 24932 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0883_
timestamp 0
transform 1 0 25024 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0884_
timestamp 0
transform 1 0 25208 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0885_
timestamp 0
transform 1 0 27416 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 0
transform 1 0 26956 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0887_
timestamp 0
transform 1 0 27692 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0888_
timestamp 0
transform 1 0 27232 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0889_
timestamp 0
transform -1 0 29440 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp 0
transform 1 0 29532 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0891_
timestamp 0
transform -1 0 31924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0892_
timestamp 0
transform 1 0 31372 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0893_
timestamp 0
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0894_
timestamp 0
transform 1 0 32844 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0895_
timestamp 0
transform -1 0 33764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 0
transform 1 0 33212 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0897_
timestamp 0
transform 1 0 32936 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0898_
timestamp 0
transform -1 0 34408 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 0
transform 1 0 34316 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0900_
timestamp 0
transform -1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0901_
timestamp 0
transform -1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 0
transform 1 0 31372 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0903_
timestamp 0
transform 1 0 30820 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0904_
timestamp 0
transform 1 0 28336 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0905_
timestamp 0
transform -1 0 28704 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0907_
timestamp 0
transform 1 0 25300 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0908_
timestamp 0
transform 1 0 25484 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0909_
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0910_
timestamp 0
transform -1 0 23368 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0911_
timestamp 0
transform -1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0912_
timestamp 0
transform 1 0 22080 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0913_
timestamp 0
transform 1 0 21804 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp 0
transform 1 0 22816 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0915_
timestamp 0
transform -1 0 24288 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0916_
timestamp 0
transform 1 0 25668 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0917_
timestamp 0
transform 1 0 24932 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp 0
transform -1 0 28244 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0919_
timestamp 0
transform 1 0 28244 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 0
transform -1 0 30912 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0921_
timestamp 0
transform -1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0922_
timestamp 0
transform 1 0 29072 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0923_
timestamp 0
transform -1 0 31188 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0924_
timestamp 0
transform -1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0925_
timestamp 0
transform 1 0 28152 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0926_
timestamp 0
transform -1 0 28152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0927_
timestamp 0
transform 1 0 26220 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp 0
transform 1 0 25576 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0929_
timestamp 0
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0930_
timestamp 0
transform 1 0 22356 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0931_
timestamp 0
transform -1 0 22264 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0932_
timestamp 0
transform -1 0 21068 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0933_
timestamp 0
transform -1 0 19136 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0934_
timestamp 0
transform -1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0935_
timestamp 0
transform -1 0 21436 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 0
transform 1 0 18308 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0937_
timestamp 0
transform 1 0 17296 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 0
transform -1 0 17480 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 0
transform 1 0 15640 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 0
transform 1 0 15456 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0941_
timestamp 0
transform -1 0 17848 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 0
transform 1 0 16836 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0943_
timestamp 0
transform 1 0 15548 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0944_
timestamp 0
transform 1 0 14536 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 0
transform 1 0 13064 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0947_
timestamp 0
transform 1 0 13524 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 0
transform -1 0 13892 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0951_
timestamp 0
transform 1 0 12972 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 0
transform 1 0 12604 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0953_
timestamp 0
transform 1 0 12512 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 0
transform 1 0 12788 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0955_
timestamp 0
transform -1 0 15364 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 0
transform 1 0 14812 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0957_
timestamp 0
transform -1 0 17480 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp 0
transform 1 0 16284 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0959_
timestamp 0
transform -1 0 18308 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 0
transform 1 0 18492 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0961_
timestamp 0
transform 1 0 19504 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0962_
timestamp 0
transform 1 0 19688 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0963_
timestamp 0
transform 1 0 20884 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0964_
timestamp 0
transform -1 0 23092 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0965_
timestamp 0
transform -1 0 23920 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0966_
timestamp 0
transform 1 0 24564 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0967_
timestamp 0
transform 1 0 25852 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp 0
transform 1 0 25852 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp 0
transform 1 0 24380 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp 0
transform 1 0 23092 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 0
transform 1 0 23092 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0972_
timestamp 0
transform 1 0 22080 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 0
transform 1 0 21804 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0974_
timestamp 0
transform 1 0 21804 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0975_
timestamp 0
transform 1 0 20332 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0976_
timestamp 0
transform 1 0 19228 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0977_
timestamp 0
transform 1 0 17848 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0978_
timestamp 0
transform 1 0 16744 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0979_
timestamp 0
transform 1 0 16652 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0980_
timestamp 0
transform 1 0 14444 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0981_
timestamp 0
transform 1 0 13340 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp 0
transform 1 0 12696 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0983_
timestamp 0
transform 1 0 12696 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp 0
transform 1 0 11868 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0985_
timestamp 0
transform -1 0 13524 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0986_
timestamp 0
transform 1 0 12052 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0987_
timestamp 0
transform 1 0 13156 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0988_
timestamp 0
transform 1 0 14168 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0989_
timestamp 0
transform 1 0 15640 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 0
transform 1 0 16652 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0991_
timestamp 0
transform 1 0 15732 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0992_
timestamp 0
transform -1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0993_
timestamp 0
transform 1 0 17480 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp 0
transform 1 0 16652 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 0
transform -1 0 18308 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 0
transform 1 0 19228 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0997_
timestamp 0
transform 1 0 19688 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 0
transform 1 0 19228 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp 0
transform 1 0 18216 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 0
transform 1 0 17940 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 0
transform 1 0 18216 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp 0
transform -1 0 20056 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1003_
timestamp 0
transform -1 0 21528 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 0
transform 1 0 20884 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp 0
transform 1 0 23644 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 0
transform -1 0 25300 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1007_
timestamp 0
transform 1 0 23184 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 0
transform -1 0 26128 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1009_
timestamp 0
transform 1 0 25760 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1010_
timestamp 0
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1011_
timestamp 0
transform 1 0 28336 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1012_
timestamp 0
transform 1 0 29532 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1013_
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1014_
timestamp 0
transform 1 0 3128 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1015_
timestamp 0
transform -1 0 3496 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1016_
timestamp 0
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1017_
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1018_
timestamp 0
transform -1 0 3496 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 0
transform -1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1020_
timestamp 0
transform -1 0 2392 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1021_
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1022_
timestamp 0
transform -1 0 4324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1023_
timestamp 0
transform 1 0 4324 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1024_
timestamp 0
transform 1 0 4508 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1025_
timestamp 0
transform -1 0 4416 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1026_
timestamp 0
transform 1 0 5060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1027_
timestamp 0
transform -1 0 4416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1028_
timestamp 0
transform -1 0 2484 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1029_
timestamp 0
transform -1 0 3220 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1030_
timestamp 0
transform -1 0 2024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1031_
timestamp 0
transform 1 0 2392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1032_
timestamp 0
transform -1 0 2484 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1033_
timestamp 0
transform -1 0 30820 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1034_
timestamp 0
transform -1 0 6256 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1035_
timestamp 0
transform -1 0 5980 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1036_
timestamp 0
transform -1 0 5520 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1037_
timestamp 0
transform 1 0 5520 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1038_
timestamp 0
transform 1 0 7084 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1039_
timestamp 0
transform 1 0 7728 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1040_
timestamp 0
transform -1 0 7544 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 0
transform -1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 0
transform -1 0 9568 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1043_
timestamp 0
transform -1 0 9476 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1044_
timestamp 0
transform 1 0 9200 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1045_
timestamp 0
transform 1 0 9936 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1046_
timestamp 0
transform -1 0 11132 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1047_
timestamp 0
transform 1 0 10488 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1048_
timestamp 0
transform 1 0 10212 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1049_
timestamp 0
transform -1 0 10948 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1050_
timestamp 0
transform -1 0 11316 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1051_
timestamp 0
transform -1 0 10304 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1052_
timestamp 0
transform -1 0 9200 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 0
transform -1 0 10028 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1054_
timestamp 0
transform -1 0 8740 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1055_
timestamp 0
transform -1 0 7728 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _1056_
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1057_
timestamp 0
transform 1 0 1840 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1058_
timestamp 0
transform 1 0 1380 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1059_
timestamp 0
transform 1 0 1840 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1060_
timestamp 0
transform 1 0 3404 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1061_
timestamp 0
transform 1 0 5152 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1062_
timestamp 0
transform -1 0 6716 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1063_
timestamp 0
transform -1 0 8188 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1064_
timestamp 0
transform 1 0 6808 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1065_
timestamp 0
transform 1 0 4140 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1066_
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1067_
timestamp 0
transform 1 0 4968 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1068_
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1069_
timestamp 0
transform 1 0 3128 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1070_
timestamp 0
transform 1 0 3128 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1071_
timestamp 0
transform -1 0 6440 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1072_
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1073_
timestamp 0
transform -1 0 10028 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1074_
timestamp 0
transform 1 0 6992 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1075_
timestamp 0
transform -1 0 11408 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1076_
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1077_
timestamp 0
transform 1 0 10488 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1078_
timestamp 0
transform 1 0 10304 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1079_
timestamp 0
transform 1 0 6992 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1080_
timestamp 0
transform 1 0 7912 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1081_
timestamp 0
transform 1 0 10304 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1082_
timestamp 0
transform 1 0 10304 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1083_
timestamp 0
transform 1 0 8740 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1084_
timestamp 0
transform 1 0 7452 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1085_
timestamp 0
transform 1 0 6716 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1086_
timestamp 0
transform 1 0 8096 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1087_
timestamp 0
transform 1 0 9660 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1088_
timestamp 0
transform 1 0 30176 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1089_
timestamp 0
transform 1 0 29992 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1090_
timestamp 0
transform 1 0 28428 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1091_
timestamp 0
transform 1 0 30176 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1092_
timestamp 0
transform 1 0 32108 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1093_
timestamp 0
transform -1 0 35420 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1094_
timestamp 0
transform 1 0 33948 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 0
transform 1 0 32292 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1096_
timestamp 0
transform 1 0 28152 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 0
transform 1 0 29532 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1098_
timestamp 0
transform 1 0 28428 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1099_
timestamp 0
transform 1 0 29532 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 0
transform 1 0 31372 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 0
transform -1 0 33856 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 0
transform 1 0 34500 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 0
transform 1 0 32660 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1104_
timestamp 0
transform 1 0 32108 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 0
transform 1 0 26956 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 0
transform 1 0 25668 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 0
transform 1 0 26036 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 0
transform -1 0 28336 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 0
transform 1 0 26956 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 0
transform -1 0 28704 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 0
transform -1 0 28796 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 0
transform -1 0 29072 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 0
transform -1 0 30360 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1115_
timestamp 0
transform -1 0 31372 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1116_
timestamp 0
transform -1 0 32384 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1117_
timestamp 0
transform -1 0 34224 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 0
transform -1 0 34592 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 0
transform 1 0 33396 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 0
transform 1 0 34408 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 0
transform 1 0 32568 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 0
transform 1 0 31740 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 0
transform -1 0 31740 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1124_
timestamp 0
transform 1 0 29532 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 0
transform 1 0 28612 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 0
transform 1 0 27508 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 0
transform 1 0 27048 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 0
transform 1 0 26220 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 0
transform 1 0 24932 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1131_
timestamp 0
transform 1 0 23184 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1132_
timestamp 0
transform 1 0 22540 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1133_
timestamp 0
transform 1 0 24380 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 0
transform 1 0 24380 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 0
transform 1 0 24288 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 0
transform -1 0 24288 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1139_
timestamp 0
transform 1 0 21528 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1140_
timestamp 0
transform 1 0 21896 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1141_
timestamp 0
transform -1 0 23644 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 0
transform 1 0 20608 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1143_
timestamp 0
transform 1 0 20700 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 0
transform -1 0 21436 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 0
transform -1 0 20792 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 0
transform 1 0 19044 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1147_
timestamp 0
transform -1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1148_
timestamp 0
transform 1 0 20608 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1149_
timestamp 0
transform 1 0 19504 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1151_
timestamp 0
transform 1 0 19780 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 0
transform -1 0 25484 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 0
transform 1 0 22264 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1155_
timestamp 0
transform 1 0 22264 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1156_
timestamp 0
transform -1 0 25944 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 0
transform -1 0 26588 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 0
transform -1 0 26864 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 0
transform 1 0 24748 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 0
transform -1 0 28796 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 0
transform 1 0 27324 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 0
transform -1 0 31372 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 0
transform -1 0 31556 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1164_
timestamp 0
transform -1 0 33304 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1165_
timestamp 0
transform -1 0 34132 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 0
transform 1 0 34684 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 0
transform 1 0 34040 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 0
transform 1 0 32568 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 0
transform 1 0 32016 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 0
transform 1 0 33948 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 0
transform 1 0 32108 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 0
transform -1 0 32016 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 0
transform 1 0 30084 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 0
transform 1 0 29532 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 0
transform 1 0 27508 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 0
transform 1 0 25024 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 0
transform 1 0 24840 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 0
transform 1 0 23736 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 0
transform 1 0 22356 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 0
transform 1 0 21804 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 0
transform 1 0 22172 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 0
transform 1 0 20792 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 0
transform 1 0 18952 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 0
transform 1 0 18584 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 0
transform -1 0 20056 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1188_
timestamp 0
transform -1 0 19136 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 0
transform 1 0 16652 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 0
transform 1 0 16560 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 0
transform 1 0 15272 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 0
transform 1 0 14076 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 0
transform 1 0 13800 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 0
transform 1 0 14260 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 0
transform 1 0 13800 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1197_
timestamp 0
transform 1 0 13616 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1199_
timestamp 0
transform 1 0 13892 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1200_
timestamp 0
transform 1 0 14352 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 0
transform 1 0 14260 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 0
transform -1 0 15916 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1203_
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 0
transform 1 0 14260 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 0
transform 1 0 14628 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 0
transform 1 0 14076 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 0
transform 1 0 13800 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 0
transform -1 0 16836 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1210_
timestamp 0
transform 1 0 16836 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 0
transform 1 0 16652 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 0
transform 1 0 16928 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 0
transform 1 0 17296 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 0
transform 1 0 16836 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1215_
timestamp 0
transform -1 0 18492 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1216_
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1217_
timestamp 0
transform -1 0 18676 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 0
transform 1 0 16744 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 0
transform -1 0 18308 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 0
transform -1 0 18124 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1221_
timestamp 0
transform 1 0 16100 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1222_
timestamp 0
transform 1 0 16008 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1223_
timestamp 0
transform -1 0 21528 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1224_
timestamp 0
transform -1 0 21528 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1225_
timestamp 0
transform -1 0 21252 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1226_
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1227_
timestamp 0
transform 1 0 18952 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1228_
timestamp 0
transform -1 0 23644 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 0
transform -1 0 23184 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1230_
timestamp 0
transform -1 0 25484 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1231_
timestamp 0
transform 1 0 23368 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1232_
timestamp 0
transform -1 0 28060 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1233_
timestamp 0
transform 1 0 27416 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1234_
timestamp 0
transform 1 0 26772 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1235_
timestamp 0
transform 1 0 26680 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1236_
timestamp 0
transform 1 0 27140 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1237_
timestamp 0
transform 1 0 29808 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1238_
timestamp 0
transform 1 0 29808 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 0
transform -1 0 30636 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1240_
timestamp 0
transform 1 0 29808 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1241_
timestamp 0
transform 1 0 31648 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1242_
timestamp 0
transform 1 0 33212 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1243_
timestamp 0
transform 1 0 33672 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 0
transform 1 0 33948 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1245_
timestamp 0
transform 1 0 31464 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1246_
timestamp 0
transform 1 0 33120 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1247_
timestamp 0
transform 1 0 32568 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1248_
timestamp 0
transform 1 0 30452 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1249_
timestamp 0
transform 1 0 33672 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1250_
timestamp 0
transform 1 0 24380 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1251_
timestamp 0
transform 1 0 24380 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1252_
timestamp 0
transform 1 0 24564 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1253_
timestamp 0
transform -1 0 27416 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1254_
timestamp 0
transform 1 0 26956 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1255_
timestamp 0
transform 1 0 25852 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1256_
timestamp 0
transform 1 0 26956 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1257_
timestamp 0
transform -1 0 30820 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1258_
timestamp 0
transform -1 0 29992 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1259_
timestamp 0
transform -1 0 31924 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1260_
timestamp 0
transform 1 0 30176 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1261_
timestamp 0
transform -1 0 34224 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1262_
timestamp 0
transform 1 0 32200 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1263_
timestamp 0
transform 1 0 32108 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1264_
timestamp 0
transform 1 0 32200 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1265_
timestamp 0
transform 1 0 32108 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1266_
timestamp 0
transform 1 0 32660 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1267_
timestamp 0
transform 1 0 32752 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1268_
timestamp 0
transform 1 0 32660 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1269_
timestamp 0
transform 1 0 32108 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1270_
timestamp 0
transform 1 0 30176 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1271_
timestamp 0
transform 1 0 29532 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1272_
timestamp 0
transform 1 0 28980 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1273_
timestamp 0
transform 1 0 27140 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1274_
timestamp 0
transform 1 0 26220 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1275_
timestamp 0
transform 1 0 24932 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1276_
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1277_
timestamp 0
transform 1 0 23644 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1278_
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1279_
timestamp 0
transform 1 0 20516 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1280_
timestamp 0
transform 1 0 19872 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1281_
timestamp 0
transform 1 0 19964 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1282_
timestamp 0
transform -1 0 23828 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1283_
timestamp 0
transform -1 0 25668 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1284_
timestamp 0
transform -1 0 26220 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 0
transform 1 0 24840 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 0
transform -1 0 28796 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 0
transform -1 0 28796 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1288_
timestamp 0
transform -1 0 31004 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1289_
timestamp 0
transform -1 0 31372 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1290_
timestamp 0
transform 1 0 29716 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1291_
timestamp 0
transform 1 0 29900 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1292_
timestamp 0
transform 1 0 28980 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1293_
timestamp 0
transform 1 0 27600 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1294_
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1295_
timestamp 0
transform 1 0 25208 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1296_
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1297_
timestamp 0
transform 1 0 23736 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1298_
timestamp 0
transform 1 0 21896 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1299_
timestamp 0
transform 1 0 20700 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1300_
timestamp 0
transform 1 0 19596 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1301_
timestamp 0
transform 1 0 17756 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1302_
timestamp 0
transform -1 0 20332 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1303_
timestamp 0
transform 1 0 18492 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1304_
timestamp 0
transform 1 0 17664 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1305_
timestamp 0
transform 1 0 16928 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1306_
timestamp 0
transform 1 0 17112 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1307_
timestamp 0
transform 1 0 14904 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1308_
timestamp 0
transform 1 0 14444 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1309_
timestamp 0
transform -1 0 18216 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1310_
timestamp 0
transform 1 0 16376 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1311_
timestamp 0
transform 1 0 15272 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 0
transform 1 0 14076 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 0
transform 1 0 12236 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 0
transform 1 0 12144 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1315_
timestamp 0
transform 1 0 12144 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1316_
timestamp 0
transform 1 0 11776 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1317_
timestamp 0
transform 1 0 12788 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1318_
timestamp 0
transform -1 0 15916 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1319_
timestamp 0
transform 1 0 12144 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1320_
timestamp 0
transform 1 0 11684 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1321_
timestamp 0
transform 1 0 11500 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1322_
timestamp 0
transform 1 0 11592 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1323_
timestamp 0
transform -1 0 15548 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1324_
timestamp 0
transform 1 0 13892 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1325_
timestamp 0
transform -1 0 17572 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1326_
timestamp 0
transform 1 0 14720 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1327_
timestamp 0
transform -1 0 18492 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1328_
timestamp 0
transform -1 0 19136 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1329_
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1330_
timestamp 0
transform 1 0 19228 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1331_
timestamp 0
transform 1 0 20424 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1332_
timestamp 0
transform -1 0 23644 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1333_
timestamp 0
transform -1 0 24012 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1334_
timestamp 0
transform -1 0 25484 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1335_
timestamp 0
transform -1 0 26220 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1336_
timestamp 0
transform 1 0 24380 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 0
transform 1 0 24012 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1338_
timestamp 0
transform 1 0 22172 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1339_
timestamp 0
transform 1 0 22632 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1340_
timestamp 0
transform 1 0 21528 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1341_
timestamp 0
transform 1 0 20792 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1342_
timestamp 0
transform 1 0 20700 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1343_
timestamp 0
transform 1 0 19872 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1344_
timestamp 0
transform 1 0 18032 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1345_
timestamp 0
transform 1 0 17296 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1346_
timestamp 0
transform 1 0 15456 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1347_
timestamp 0
transform 1 0 15272 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1348_
timestamp 0
transform 1 0 14168 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1349_
timestamp 0
transform 1 0 12880 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1350_
timestamp 0
transform 1 0 11776 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1351_
timestamp 0
transform 1 0 11500 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1352_
timestamp 0
transform 1 0 11776 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1353_
timestamp 0
transform -1 0 13708 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1354_
timestamp 0
transform 1 0 11408 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1355_
timestamp 0
transform -1 0 13800 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1356_
timestamp 0
transform -1 0 14720 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1357_
timestamp 0
transform -1 0 16560 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1358_
timestamp 0
transform 1 0 14720 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1359_
timestamp 0
transform 1 0 15180 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1360_
timestamp 0
transform 1 0 14168 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1361_
timestamp 0
transform 1 0 13984 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1362_
timestamp 0
transform 1 0 15640 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1363_
timestamp 0
transform -1 0 18860 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1364_
timestamp 0
transform -1 0 19872 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1365_
timestamp 0
transform 1 0 19320 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1366_
timestamp 0
transform 1 0 18768 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1367_
timestamp 0
transform 1 0 17296 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1368_
timestamp 0
transform 1 0 17204 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1369_
timestamp 0
transform 1 0 17204 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1370_
timestamp 0
transform -1 0 20608 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1371_
timestamp 0
transform -1 0 21896 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1372_
timestamp 0
transform 1 0 19964 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1373_
timestamp 0
transform -1 0 23644 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1374_
timestamp 0
transform -1 0 25484 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1375_
timestamp 0
transform 1 0 22080 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1376_
timestamp 0
transform -1 0 26220 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1377_
timestamp 0
transform 1 0 26220 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1378_
timestamp 0
transform 1 0 28152 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1379_
timestamp 0
transform 1 0 1564 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1380_
timestamp 0
transform -1 0 3220 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1381_
timestamp 0
transform 1 0 1564 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1382_
timestamp 0
transform -1 0 4784 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1383_
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1384_
timestamp 0
transform 1 0 1656 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1385_
timestamp 0
transform 1 0 4048 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1386_
timestamp 0
transform -1 0 6992 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1387_
timestamp 0
transform -1 0 6256 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1388_
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1389_
timestamp 0
transform 1 0 2024 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1390_
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1391_
timestamp 0
transform 1 0 29532 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1392_
timestamp 0
transform 1 0 5152 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1393_
timestamp 0
transform 1 0 4968 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1394_
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1395_
timestamp 0
transform 1 0 6900 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1396_
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1397_
timestamp 0
transform 1 0 9844 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1398_
timestamp 0
transform 1 0 10580 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1399_
timestamp 0
transform 1 0 10580 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1400_
timestamp 0
transform 1 0 9568 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1401_
timestamp 0
transform 1 0 7728 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1402_
timestamp 0
transform 1 0 6256 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _1917_
timestamp 0
transform -1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform 1 0 7084 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 0
transform 1 0 9292 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 0
transform 1 0 28796 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 0
transform 1 0 21252 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 0
transform 1 0 23276 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 0
transform 1 0 7268 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 0
transform 1 0 9476 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 0
transform 1 0 21068 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 0
transform 1 0 23460 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_A_in_serial_clk
timestamp 0
transform 1 0 25024 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_B_in_serial_clk
timestamp 0
transform -1 0 25852 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 6256 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform 1 0 7728 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform -1 0 6256 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 6992 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_A_in_serial_clk
timestamp 0
transform -1 0 17664 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_B_in_serial_clk
timestamp 0
transform -1 0 15916 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_A_in_serial_clk
timestamp 0
transform -1 0 16560 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_B_in_serial_clk
timestamp 0
transform -1 0 14904 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_A_in_serial_clk
timestamp 0
transform -1 0 23092 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_B_in_serial_clk
timestamp 0
transform -1 0 20608 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_A_in_serial_clk
timestamp 0
transform 1 0 22540 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_B_in_serial_clk
timestamp 0
transform -1 0 22080 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_A_in_serial_clk
timestamp 0
transform -1 0 17388 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_B_in_serial_clk
timestamp 0
transform 1 0 14812 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_A_in_serial_clk
timestamp 0
transform -1 0 17756 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_B_in_serial_clk
timestamp 0
transform -1 0 15640 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_A_in_serial_clk
timestamp 0
transform 1 0 21896 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_B_in_serial_clk
timestamp 0
transform 1 0 20332 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_A_in_serial_clk
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_B_in_serial_clk
timestamp 0
transform 1 0 20516 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_A_in_serial_clk
timestamp 0
transform -1 0 28520 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_B_in_serial_clk
timestamp 0
transform 1 0 25760 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_A_in_serial_clk
timestamp 0
transform 1 0 27416 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_B_in_serial_clk
timestamp 0
transform 1 0 25668 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_A_in_serial_clk
timestamp 0
transform -1 0 33120 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_B_in_serial_clk
timestamp 0
transform 1 0 31556 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_A_in_serial_clk
timestamp 0
transform 1 0 32660 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_B_in_serial_clk
timestamp 0
transform 1 0 30912 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_A_in_serial_clk
timestamp 0
transform 1 0 26956 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_B_in_serial_clk
timestamp 0
transform 1 0 25852 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_A_in_serial_clk
timestamp 0
transform -1 0 28244 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_B_in_serial_clk
timestamp 0
transform -1 0 27968 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_A_in_serial_clk
timestamp 0
transform 1 0 33488 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_B_in_serial_clk
timestamp 0
transform 1 0 31372 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_A_in_serial_clk
timestamp 0
transform -1 0 33488 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_B_in_serial_clk
timestamp 0
transform 1 0 32108 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_4  clkload0
timestamp 0
transform 1 0 4600 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_4  clkload1
timestamp 0
transform 1 0 3772 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload2
timestamp 0
transform 1 0 7268 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload3
timestamp 0
transform -1 0 17296 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  clkload4
timestamp 0
transform 1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  clkload5
timestamp 0
transform -1 0 14720 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  clkload6
timestamp 0
transform -1 0 21712 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  clkload7
timestamp 0
transform -1 0 26956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__bufinv_16  clkload8
timestamp 0
transform 1 0 27232 0 1 9792
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_8  clkload9
timestamp 0
transform 1 0 32936 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload10
timestamp 0
transform 1 0 32660 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload11
timestamp 0
transform -1 0 29164 0 -1 17408
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload12
timestamp 0
transform 1 0 26680 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload13
timestamp 0
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload14
timestamp 0
transform 1 0 32292 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload15
timestamp 0
transform 1 0 14904 0 1 26112
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  clkload16
timestamp 0
transform 1 0 15916 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload17
timestamp 0
transform -1 0 21712 0 -1 26112
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_6  clkload18
timestamp 0
transform 1 0 19228 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload19
timestamp 0
transform 1 0 14812 0 1 32640
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_6  clkload20
timestamp 0
transform 1 0 20148 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload21
timestamp 0
transform 1 0 20608 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload22
timestamp 0
transform -1 0 26772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload23
timestamp 0
transform 1 0 24380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload24
timestamp 0
transform 1 0 31096 0 1 25024
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload25
timestamp 0
transform 1 0 31004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_6  clkload26
timestamp 0
transform -1 0 25852 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload27
timestamp 0
transform 1 0 26036 0 1 32640
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_6  clkload28
timestamp 0
transform 1 0 31372 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload29
timestamp 0
transform 1 0 33120 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_16  clone2
timestamp 0
transform 1 0 29532 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone24
timestamp 0
transform -1 0 30636 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__nand2b_2  clone29
timestamp 0
transform 1 0 32108 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_16  clone31
timestamp 0
transform -1 0 21436 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone624
timestamp 0
transform 1 0 27140 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  clone626
timestamp 0
transform -1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  clone627
timestamp 0
transform 1 0 29808 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clone630
timestamp 0
transform -1 0 24196 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone631
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone712
timestamp 0
transform 1 0 20332 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  clone714
timestamp 0
transform -1 0 20700 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  clone716
timestamp 0
transform -1 0 21528 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  clone718
timestamp 0
transform -1 0 18952 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clone719
timestamp 0
transform -1 0 21068 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone724
timestamp 0
transform -1 0 31556 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  clone753
timestamp 0
transform 1 0 29716 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  clone792
timestamp 0
transform 1 0 30452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clone793
timestamp 0
transform -1 0 29716 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone829
timestamp 0
transform -1 0 23644 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone831
timestamp 0
transform -1 0 23644 0 -1 35904
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 0
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 0
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 0
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 0
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 0
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 0
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 0
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 0
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 0
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 0
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 0
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 0
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_377
timestamp 0
transform 1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_385
timestamp 0
transform 1 0 36524 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 0
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 0
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 0
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 0
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 0
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 0
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 0
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 0
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 0
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_305
timestamp 0
transform 1 0 29164 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_313
timestamp 0
transform 1 0 29900 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_357
timestamp 0
transform 1 0 33948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_369
timestamp 0
transform 1 0 35052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_381
timestamp 0
transform 1 0 36156 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_387
timestamp 0
transform 1 0 36708 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 0
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 0
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 0
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 0
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 0
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 0
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 0
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 0
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 0
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 0
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 0
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 0
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_334
timestamp 0
transform 1 0 31832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 0
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 0
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_377
timestamp 0
transform 1 0 35788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_385
timestamp 0
transform 1 0 36524 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 0
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 0
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 0
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 0
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 0
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 0
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 0
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 0
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_351
timestamp 0
transform 1 0 33396 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 0
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_385
timestamp 0
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_174
timestamp 0
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_186
timestamp 0
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 0
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 0
transform 1 0 20700 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_226
timestamp 0
transform 1 0 21896 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_238
timestamp 0
transform 1 0 23000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 0
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 0
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 0
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 0
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 0
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 0
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_309
timestamp 0
transform 1 0 29532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_322
timestamp 0
transform 1 0 30728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 0
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 0
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_385
timestamp 0
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 0
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_184
timestamp 0
transform 1 0 18032 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_192
timestamp 0
transform 1 0 18768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214
timestamp 0
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 0
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_265
timestamp 0
transform 1 0 25484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 0
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_301
timestamp 0
transform 1 0 28796 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_320
timestamp 0
transform 1 0 30544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 0
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_342
timestamp 0
transform 1 0 32568 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_371
timestamp 0
transform 1 0 35236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_383
timestamp 0
transform 1 0 36340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_387
timestamp 0
transform 1 0 36708 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 0
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 0
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_217
timestamp 0
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_265
timestamp 0
transform 1 0 25484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 0
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 0
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_309
timestamp 0
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_315
timestamp 0
transform 1 0 30084 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_335
timestamp 0
transform 1 0 31924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_369
timestamp 0
transform 1 0 35052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_381
timestamp 0
transform 1 0 36156 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_387
timestamp 0
transform 1 0 36708 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 0
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 0
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_175
timestamp 0
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_188
timestamp 0
transform 1 0 18400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_201
timestamp 0
transform 1 0 19596 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 0
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_234
timestamp 0
transform 1 0 22632 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_262
timestamp 0
transform 1 0 25208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 0
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 0
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_292
timestamp 0
transform 1 0 27968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_314
timestamp 0
transform 1 0 29992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_351
timestamp 0
transform 1 0 33396 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_377
timestamp 0
transform 1 0 35788 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_149
timestamp 0
transform 1 0 14812 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_162
timestamp 0
transform 1 0 16008 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_168
timestamp 0
transform 1 0 16560 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 0
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 0
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_238
timestamp 0
transform 1 0 23000 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 0
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp 0
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_291
timestamp 0
transform 1 0 27876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 0
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 0
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 0
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_313
timestamp 0
transform 1 0 29900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_320
timestamp 0
transform 1 0 30544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_327
timestamp 0
transform 1 0 31188 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_332
timestamp 0
transform 1 0 31648 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_338
timestamp 0
transform 1 0 32200 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_373
timestamp 0
transform 1 0 35420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_385
timestamp 0
transform 1 0 36524 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_149
timestamp 0
transform 1 0 14812 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 0
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_189
timestamp 0
transform 1 0 18492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 0
transform 1 0 19228 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 0
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 0
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp 0
transform 1 0 22356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 0
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_290
timestamp 0
transform 1 0 27784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_324
timestamp 0
transform 1 0 30912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_330
timestamp 0
transform 1 0 31464 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 0
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_385
timestamp 0
transform 1 0 36524 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_163
timestamp 0
transform 1 0 16100 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 0
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 0
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_273
timestamp 0
transform 1 0 26220 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_296
timestamp 0
transform 1 0 28336 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_357
timestamp 0
transform 1 0 33948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 0
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_385
timestamp 0
transform 1 0 36524 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 0
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 0
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 0
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 0
transform 1 0 18032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_197
timestamp 0
transform 1 0 19228 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_205
timestamp 0
transform 1 0 19964 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 0
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 0
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_239
timestamp 0
transform 1 0 23092 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_254
timestamp 0
transform 1 0 24472 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_262
timestamp 0
transform 1 0 25208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_285
timestamp 0
transform 1 0 27324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_307
timestamp 0
transform 1 0 29348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 0
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_352
timestamp 0
transform 1 0 33488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_377
timestamp 0
transform 1 0 35788 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_385
timestamp 0
transform 1 0 36524 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 0
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_160
timestamp 0
transform 1 0 15824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 0
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 0
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_222
timestamp 0
transform 1 0 21528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 0
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_274
timestamp 0
transform 1 0 26312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_301
timestamp 0
transform 1 0 28796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 0
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_369
timestamp 0
transform 1 0 35052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_381
timestamp 0
transform 1 0 36156 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_387
timestamp 0
transform 1 0 36708 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_133
timestamp 0
transform 1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_156
timestamp 0
transform 1 0 15456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_173
timestamp 0
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 0
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_249
timestamp 0
transform 1 0 24012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_273
timestamp 0
transform 1 0 26220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 0
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_370
timestamp 0
transform 1 0 35144 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_382
timestamp 0
transform 1 0 36248 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 0
transform 1 0 14628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_160
timestamp 0
transform 1 0 15824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_183
timestamp 0
transform 1 0 17940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 0
transform 1 0 20424 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_232
timestamp 0
transform 1 0 22448 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 0
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_273
timestamp 0
transform 1 0 26220 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_281
timestamp 0
transform 1 0 26956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_309
timestamp 0
transform 1 0 29532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 0
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_375
timestamp 0
transform 1 0 35604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_387
timestamp 0
transform 1 0 36708 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 0
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_187
timestamp 0
transform 1 0 18308 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 0
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_246
timestamp 0
transform 1 0 23736 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_254
timestamp 0
transform 1 0 24472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_266
timestamp 0
transform 1 0 25576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_270
timestamp 0
transform 1 0 25944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_285
timestamp 0
transform 1 0 27324 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_321
timestamp 0
transform 1 0 30636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_337
timestamp 0
transform 1 0 32108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_383
timestamp 0
transform 1 0 36340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_387
timestamp 0
transform 1 0 36708 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 0
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 0
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_265
timestamp 0
transform 1 0 25484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_271
timestamp 0
transform 1 0 26036 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 0
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 0
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 0
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_377
timestamp 0
transform 1 0 35788 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_385
timestamp 0
transform 1 0 36524 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_177
timestamp 0
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_210
timestamp 0
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 0
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 0
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 0
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_281
timestamp 0
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_304
timestamp 0
transform 1 0 29072 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_316
timestamp 0
transform 1 0 30176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_320
timestamp 0
transform 1 0 30544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_324
timestamp 0
transform 1 0 30912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 0
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 0
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 0
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 0
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 0
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_385
timestamp 0
transform 1 0 36524 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_149
timestamp 0
transform 1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_164
timestamp 0
transform 1 0 16192 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 0
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 0
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_242
timestamp 0
transform 1 0 23368 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 0
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 0
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_329
timestamp 0
transform 1 0 31372 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_341
timestamp 0
transform 1 0 32476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_377
timestamp 0
transform 1 0 35788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_385
timestamp 0
transform 1 0 36524 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 0
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_137
timestamp 0
transform 1 0 13708 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_143
timestamp 0
transform 1 0 14260 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 0
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_177
timestamp 0
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 0
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 0
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_237
timestamp 0
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 0
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 0
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_290
timestamp 0
transform 1 0 27784 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_330
timestamp 0
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_349
timestamp 0
transform 1 0 33212 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_371
timestamp 0
transform 1 0 35236 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_383
timestamp 0
transform 1 0 36340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_387
timestamp 0
transform 1 0 36708 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 0
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 0
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 0
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_149
timestamp 0
transform 1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_164
timestamp 0
transform 1 0 16192 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 0
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 0
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 0
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_234
timestamp 0
transform 1 0 22632 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 0
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 0
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 0
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_289
timestamp 0
transform 1 0 27692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 0
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 0
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 0
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_317
timestamp 0
transform 1 0 30268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 0
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_374
timestamp 0
transform 1 0 35512 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_386
timestamp 0
transform 1 0 36616 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_6
timestamp 0
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 0
transform 1 0 2760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_40
timestamp 0
transform 1 0 4784 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_77
timestamp 0
transform 1 0 8188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_85
timestamp 0
transform 1 0 8924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_91
timestamp 0
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp 0
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_137
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 0
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 0
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_200
timestamp 0
transform 1 0 19504 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 0
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_249
timestamp 0
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_257
timestamp 0
transform 1 0 24748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 0
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_290
timestamp 0
transform 1 0 27784 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_318
timestamp 0
transform 1 0 30360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 0
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_346
timestamp 0
transform 1 0 32936 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_359
timestamp 0
transform 1 0 34132 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_371
timestamp 0
transform 1 0 35236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_383
timestamp 0
transform 1 0 36340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_387
timestamp 0
transform 1 0 36708 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_10
timestamp 0
transform 1 0 2024 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 0
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 0
transform 1 0 4048 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 0
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_62
timestamp 0
transform 1 0 6808 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_74
timestamp 0
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 0
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_115
timestamp 0
transform 1 0 11684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_127
timestamp 0
transform 1 0 12788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_161
timestamp 0
transform 1 0 15916 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_169
timestamp 0
transform 1 0 16652 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 0
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 0
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_293
timestamp 0
transform 1 0 28060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 0
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 0
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_353
timestamp 0
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 0
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_377
timestamp 0
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_385
timestamp 0
transform 1 0 36524 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_21
timestamp 0
transform 1 0 3036 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_79
timestamp 0
transform 1 0 8372 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_101
timestamp 0
transform 1 0 10396 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 0
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 0
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 0
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_193
timestamp 0
transform 1 0 18860 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 0
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 0
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_225
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_246
timestamp 0
transform 1 0 23736 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_258
timestamp 0
transform 1 0 24840 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 0
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 0
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_281
timestamp 0
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_302
timestamp 0
transform 1 0 28888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_310
timestamp 0
transform 1 0 29624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_331
timestamp 0
transform 1 0 31556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 0
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_337
timestamp 0
transform 1 0 32108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_341
timestamp 0
transform 1 0 32476 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_382
timestamp 0
transform 1 0 36248 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 0
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_36
timestamp 0
transform 1 0 4416 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_48
timestamp 0
transform 1 0 5520 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_60
timestamp 0
transform 1 0 6624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_95
timestamp 0
transform 1 0 9844 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_123
timestamp 0
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 0
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 0
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 0
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 0
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 0
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_277
timestamp 0
transform 1 0 26588 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_285
timestamp 0
transform 1 0 27324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 0
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_350
timestamp 0
transform 1 0 33304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 0
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 0
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_377
timestamp 0
transform 1 0 35788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_385
timestamp 0
transform 1 0 36524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_11
timestamp 0
transform 1 0 2116 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_23
timestamp 0
transform 1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 0
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 0
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 0
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_63
timestamp 0
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_70
timestamp 0
transform 1 0 7544 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_82
timestamp 0
transform 1 0 8648 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_94
timestamp 0
transform 1 0 9752 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 0
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 0
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 0
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_189
timestamp 0
transform 1 0 18492 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 0
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 0
transform 1 0 21252 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_233
timestamp 0
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 0
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 0
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_292
timestamp 0
transform 1 0 27968 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 0
transform 1 0 28520 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_331
timestamp 0
transform 1 0 31556 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_346
timestamp 0
transform 1 0 32936 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_358
timestamp 0
transform 1 0 34040 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_370
timestamp 0
transform 1 0 35144 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_382
timestamp 0
transform 1 0 36248 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_14
timestamp 0
transform 1 0 2392 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 0
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_43
timestamp 0
transform 1 0 5060 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_67
timestamp 0
transform 1 0 7268 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_75
timestamp 0
transform 1 0 8004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_88
timestamp 0
transform 1 0 9200 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_100
timestamp 0
transform 1 0 10304 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_123
timestamp 0
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 0
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_161
timestamp 0
transform 1 0 15916 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 0
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_230
timestamp 0
transform 1 0 22264 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 0
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 0
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 0
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 0
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 0
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_377
timestamp 0
transform 1 0 35788 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_383
timestamp 0
transform 1 0 36340 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_26
timestamp 0
transform 1 0 3496 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 0
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_97
timestamp 0
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 0
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 0
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_200
timestamp 0
transform 1 0 19504 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 0
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 0
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_245
timestamp 0
transform 1 0 23644 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_257
timestamp 0
transform 1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_314
timestamp 0
transform 1 0 29992 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_377
timestamp 0
transform 1 0 35788 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_385
timestamp 0
transform 1 0 36524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_11
timestamp 0
transform 1 0 2116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 0
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_47
timestamp 0
transform 1 0 5428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_55
timestamp 0
transform 1 0 6164 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 0
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_100
timestamp 0
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_111
timestamp 0
transform 1 0 11316 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_123
timestamp 0
transform 1 0 12420 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp 0
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_166
timestamp 0
transform 1 0 16376 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_174
timestamp 0
transform 1 0 17112 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_209
timestamp 0
transform 1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_232
timestamp 0
transform 1 0 22448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_240
timestamp 0
transform 1 0 23184 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 0
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_277
timestamp 0
transform 1 0 26588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 0
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 0
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_335
timestamp 0
transform 1 0 31924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_345
timestamp 0
transform 1 0 32844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 0
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 0
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 0
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_385
timestamp 0
transform 1 0 36524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_6
timestamp 0
transform 1 0 1656 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 0
transform 1 0 14444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_192
timestamp 0
transform 1 0 18768 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_204
timestamp 0
transform 1 0 19872 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 0
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_229
timestamp 0
transform 1 0 22172 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 0
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 0
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_321
timestamp 0
transform 1 0 30636 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_337
timestamp 0
transform 1 0 32108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_341
timestamp 0
transform 1 0 32476 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_362
timestamp 0
transform 1 0 34408 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_374
timestamp 0
transform 1 0 35512 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_386
timestamp 0
transform 1 0 36616 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 0
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 0
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 0
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 0
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 0
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_229
timestamp 0
transform 1 0 22172 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 0
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 0
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_277
timestamp 0
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_285
timestamp 0
transform 1 0 27324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 0
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_329
timestamp 0
transform 1 0 31372 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_335
timestamp 0
transform 1 0 31924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 0
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_374
timestamp 0
transform 1 0 35512 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_386
timestamp 0
transform 1 0 36616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_30
timestamp 0
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_97
timestamp 0
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 0
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_190
timestamp 0
transform 1 0 18584 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_202
timestamp 0
transform 1 0 19688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_206
timestamp 0
transform 1 0 20056 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 0
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 0
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_237
timestamp 0
transform 1 0 22908 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_250
timestamp 0
transform 1 0 24104 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_258
timestamp 0
transform 1 0 24840 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_281
timestamp 0
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_289
timestamp 0
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 0
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_349
timestamp 0
transform 1 0 33212 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_357
timestamp 0
transform 1 0 33948 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_378
timestamp 0
transform 1 0 35880 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_386
timestamp 0
transform 1 0 36616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 0
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_17
timestamp 0
transform 1 0 2668 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 0
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 0
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 0
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 0
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 0
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_93
timestamp 0
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_99
timestamp 0
transform 1 0 10212 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_111
timestamp 0
transform 1 0 11316 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_123
timestamp 0
transform 1 0 12420 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 0
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 0
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 0
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_217
timestamp 0
transform 1 0 21068 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_229
timestamp 0
transform 1 0 22172 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 0
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 0
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 0
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 0
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 0
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 0
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 0
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_377
timestamp 0
transform 1 0 35788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_385
timestamp 0
transform 1 0 36524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp 0
transform 1 0 1748 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 0
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_91
timestamp 0
transform 1 0 9476 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_137
timestamp 0
transform 1 0 13708 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_177
timestamp 0
transform 1 0 17388 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_190
timestamp 0
transform 1 0 18584 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_202
timestamp 0
transform 1 0 19688 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 0
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_265
timestamp 0
transform 1 0 25484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 0
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_301
timestamp 0
transform 1 0 28796 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_309
timestamp 0
transform 1 0 29532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_331
timestamp 0
transform 1 0 31556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 0
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 0
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_371
timestamp 0
transform 1 0 35236 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_383
timestamp 0
transform 1 0 36340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_387
timestamp 0
transform 1 0 36708 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 0
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_33
timestamp 0
transform 1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_37
timestamp 0
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_70
timestamp 0
transform 1 0 7544 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_76
timestamp 0
transform 1 0 8096 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_93
timestamp 0
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_117
timestamp 0
transform 1 0 11868 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_129
timestamp 0
transform 1 0 12972 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_137
timestamp 0
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 0
transform 1 0 14812 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 0
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 0
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_222
timestamp 0
transform 1 0 21528 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_240
timestamp 0
transform 1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 0
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_277
timestamp 0
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 0
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_329
timestamp 0
transform 1 0 31372 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 0
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_385
timestamp 0
transform 1 0 36524 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_15
timestamp 0
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_21
timestamp 0
transform 1 0 3036 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_42
timestamp 0
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 0
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_63
timestamp 0
transform 1 0 6900 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_75
timestamp 0
transform 1 0 8004 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_83
timestamp 0
transform 1 0 8740 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_97
timestamp 0
transform 1 0 10028 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 0
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 0
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 0
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 0
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 0
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 0
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 0
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 0
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 0
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 0
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 0
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 0
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_293
timestamp 0
transform 1 0 28060 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_303
timestamp 0
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_315
timestamp 0
transform 1 0 30084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 0
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 0
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_348
timestamp 0
transform 1 0 33120 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_360
timestamp 0
transform 1 0 34224 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_372
timestamp 0
transform 1 0 35328 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_384
timestamp 0
transform 1 0 36432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 0
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_39
timestamp 0
transform 1 0 4692 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_45
timestamp 0
transform 1 0 5244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_64
timestamp 0
transform 1 0 6992 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_70
timestamp 0
transform 1 0 7544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 0
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_97
timestamp 0
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_101
timestamp 0
transform 1 0 10396 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_122
timestamp 0
transform 1 0 12328 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 0
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 0
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_155
timestamp 0
transform 1 0 15364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp 0
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 0
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_233
timestamp 0
transform 1 0 22540 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_239
timestamp 0
transform 1 0 23092 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_282
timestamp 0
transform 1 0 27048 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 0
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 0
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 0
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 0
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 0
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 0
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_377
timestamp 0
transform 1 0 35788 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_385
timestamp 0
transform 1 0 36524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_7
timestamp 0
transform 1 0 1748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_11
timestamp 0
transform 1 0 2116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_42
timestamp 0
transform 1 0 4968 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 0
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 0
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 0
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 0
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_180
timestamp 0
transform 1 0 17664 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 0
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 0
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 0
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_301
timestamp 0
transform 1 0 28796 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_323
timestamp 0
transform 1 0 30820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 0
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_357
timestamp 0
transform 1 0 33948 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_369
timestamp 0
transform 1 0 35052 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_381
timestamp 0
transform 1 0 36156 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_387
timestamp 0
transform 1 0 36708 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 0
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_32
timestamp 0
transform 1 0 4048 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_38
timestamp 0
transform 1 0 4600 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_62
timestamp 0
transform 1 0 6808 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_99
timestamp 0
transform 1 0 10212 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 0
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_174
timestamp 0
transform 1 0 17112 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_182
timestamp 0
transform 1 0 17848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_217
timestamp 0
transform 1 0 21068 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_230
timestamp 0
transform 1 0 22264 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_240
timestamp 0
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 0
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 0
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 0
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 0
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_333
timestamp 0
transform 1 0 31740 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_341
timestamp 0
transform 1 0 32476 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 0
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 0
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_377
timestamp 0
transform 1 0 35788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_385
timestamp 0
transform 1 0 36524 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_13
timestamp 0
transform 1 0 2300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_25
timestamp 0
transform 1 0 3404 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_37
timestamp 0
transform 1 0 4508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_41
timestamp 0
transform 1 0 4876 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 0
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_62
timestamp 0
transform 1 0 6808 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_74
timestamp 0
transform 1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_80
timestamp 0
transform 1 0 8464 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_84
timestamp 0
transform 1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_92
timestamp 0
transform 1 0 9568 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 0
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_129
timestamp 0
transform 1 0 12972 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_139
timestamp 0
transform 1 0 13892 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_151
timestamp 0
transform 1 0 14996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_155
timestamp 0
transform 1 0 15364 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 0
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_182
timestamp 0
transform 1 0 17848 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_188
timestamp 0
transform 1 0 18400 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_209
timestamp 0
transform 1 0 20332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 0
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_261
timestamp 0
transform 1 0 25116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 0
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_290
timestamp 0
transform 1 0 27784 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_302
timestamp 0
transform 1 0 28888 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_314
timestamp 0
transform 1 0 29992 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_327
timestamp 0
transform 1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 0
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_370
timestamp 0
transform 1 0 35144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_382
timestamp 0
transform 1 0 36248 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 0
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_73
timestamp 0
transform 1 0 7820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 0
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 0
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_109
timestamp 0
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_117
timestamp 0
transform 1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_165
timestamp 0
transform 1 0 16284 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_186
timestamp 0
transform 1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 0
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_209
timestamp 0
transform 1 0 20332 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 0
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_293
timestamp 0
transform 1 0 28060 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_338
timestamp 0
transform 1 0 32200 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 0
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_377
timestamp 0
transform 1 0 35788 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_385
timestamp 0
transform 1 0 36524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_34
timestamp 0
transform 1 0 4232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_47
timestamp 0
transform 1 0 5428 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_61
timestamp 0
transform 1 0 6716 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_82
timestamp 0
transform 1 0 8648 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_94
timestamp 0
transform 1 0 9752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 0
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_144
timestamp 0
transform 1 0 14352 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_156
timestamp 0
transform 1 0 15456 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 0
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 0
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 0
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 0
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 0
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_337
timestamp 0
transform 1 0 32108 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_363
timestamp 0
transform 1 0 34500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_375
timestamp 0
transform 1 0 35604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_387
timestamp 0
transform 1 0 36708 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_6
timestamp 0
transform 1 0 1656 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_14
timestamp 0
transform 1 0 2392 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 0
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_49
timestamp 0
transform 1 0 5612 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_67
timestamp 0
transform 1 0 7268 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 0
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 0
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 0
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_106
timestamp 0
transform 1 0 10856 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_114
timestamp 0
transform 1 0 11592 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 0
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_170
timestamp 0
transform 1 0 16744 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 0
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 0
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_212
timestamp 0
transform 1 0 20608 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_242
timestamp 0
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 0
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_279
timestamp 0
transform 1 0 26772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 0
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 0
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 0
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_324
timestamp 0
transform 1 0 30912 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 0
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 0
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_377
timestamp 0
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_385
timestamp 0
transform 1 0 36524 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_23
timestamp 0
transform 1 0 3220 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_64
timestamp 0
transform 1 0 6992 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_73
timestamp 0
transform 1 0 7820 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_125
timestamp 0
transform 1 0 12604 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_147
timestamp 0
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 0
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 0
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_178
timestamp 0
transform 1 0 17480 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_249
timestamp 0
transform 1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 0
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 0
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_287
timestamp 0
transform 1 0 27508 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_300
timestamp 0
transform 1 0 28704 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_357
timestamp 0
transform 1 0 33948 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_369
timestamp 0
transform 1 0 35052 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_381
timestamp 0
transform 1 0 36156 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_387
timestamp 0
transform 1 0 36708 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_18
timestamp 0
transform 1 0 2760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 0
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_53
timestamp 0
transform 1 0 5980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_63
timestamp 0
transform 1 0 6900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_93
timestamp 0
transform 1 0 9660 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_99
timestamp 0
transform 1 0 10212 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_120
timestamp 0
transform 1 0 12144 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_128
timestamp 0
transform 1 0 12880 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 0
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 0
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_234
timestamp 0
transform 1 0 22632 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 0
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 0
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_279
timestamp 0
transform 1 0 26772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 0
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 0
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 0
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_342
timestamp 0
transform 1 0 32568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_355
timestamp 0
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 0
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 0
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_377
timestamp 0
transform 1 0 35788 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_385
timestamp 0
transform 1 0 36524 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_23
timestamp 0
transform 1 0 3220 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_35
timestamp 0
transform 1 0 4324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_45
timestamp 0
transform 1 0 5244 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_62
timestamp 0
transform 1 0 6808 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_75
timestamp 0
transform 1 0 8004 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_84
timestamp 0
transform 1 0 8832 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 0
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 0
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_129
timestamp 0
transform 1 0 12972 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_175
timestamp 0
transform 1 0 17204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_185
timestamp 0
transform 1 0 18124 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_196
timestamp 0
transform 1 0 19136 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 0
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 0
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 0
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 0
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_358
timestamp 0
transform 1 0 34040 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_370
timestamp 0
transform 1 0 35144 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_382
timestamp 0
transform 1 0 36248 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_7
timestamp 0
transform 1 0 1748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_34
timestamp 0
transform 1 0 4232 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_42
timestamp 0
transform 1 0 4968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_53
timestamp 0
transform 1 0 5980 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 0
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 0
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_99
timestamp 0
transform 1 0 10212 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_161
timestamp 0
transform 1 0 15916 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 0
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 0
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 0
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_237
timestamp 0
transform 1 0 22908 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_257
timestamp 0
transform 1 0 24748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_278
timestamp 0
transform 1 0 26680 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 0
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_329
timestamp 0
transform 1 0 31372 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_337
timestamp 0
transform 1 0 32108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_358
timestamp 0
transform 1 0 34040 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 0
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_377
timestamp 0
transform 1 0 35788 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_385
timestamp 0
transform 1 0 36524 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 0
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_9
timestamp 0
transform 1 0 1932 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_26
timestamp 0
transform 1 0 3496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_36
timestamp 0
transform 1 0 4416 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_44
timestamp 0
transform 1 0 5152 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_64
timestamp 0
transform 1 0 6992 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_76
timestamp 0
transform 1 0 8096 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_82
timestamp 0
transform 1 0 8648 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 0
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 0
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_135
timestamp 0
transform 1 0 13524 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_147
timestamp 0
transform 1 0 14628 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_189
timestamp 0
transform 1 0 18492 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 0
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 0
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 0
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 0
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_261
timestamp 0
transform 1 0 25116 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 0
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 0
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_293
timestamp 0
transform 1 0 28060 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_314
timestamp 0
transform 1 0 29992 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 0
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_357
timestamp 0
transform 1 0 33948 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_369
timestamp 0
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_381
timestamp 0
transform 1 0 36156 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_387
timestamp 0
transform 1 0 36708 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 0
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_9
timestamp 0
transform 1 0 1932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_22
timestamp 0
transform 1 0 3128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_41
timestamp 0
transform 1 0 4876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_49
timestamp 0
transform 1 0 5612 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_56
timestamp 0
transform 1 0 6256 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_68
timestamp 0
transform 1 0 7360 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 0
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 0
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 0
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 0
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_121
timestamp 0
transform 1 0 12236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_134
timestamp 0
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 0
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_158
timestamp 0
transform 1 0 15640 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_170
timestamp 0
transform 1 0 16744 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_48_197
timestamp 0
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_209
timestamp 0
transform 1 0 20332 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 0
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_273
timestamp 0
transform 1 0 26220 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_281
timestamp 0
transform 1 0 26956 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_293
timestamp 0
transform 1 0 28060 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_309
timestamp 0
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_335
timestamp 0
transform 1 0 31924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_355
timestamp 0
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 0
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 0
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 0
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_385
timestamp 0
transform 1 0 36524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_23
timestamp 0
transform 1 0 3220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_29
timestamp 0
transform 1 0 3772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_35
timestamp 0
transform 1 0 4324 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 0
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 0
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_89
timestamp 0
transform 1 0 9292 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_98
timestamp 0
transform 1 0 10120 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 0
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 0
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 0
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_121
timestamp 0
transform 1 0 12236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_133
timestamp 0
transform 1 0 13340 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 0
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 0
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_178
timestamp 0
transform 1 0 17480 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_186
timestamp 0
transform 1 0 18216 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_198
timestamp 0
transform 1 0 19320 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_211
timestamp 0
transform 1 0 20516 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 0
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 0
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_265
timestamp 0
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 0
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 0
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_337
timestamp 0
transform 1 0 32108 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_358
timestamp 0
transform 1 0 34040 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_370
timestamp 0
transform 1 0 35144 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_382
timestamp 0
transform 1 0 36248 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 0
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_7
timestamp 0
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_43
timestamp 0
transform 1 0 5060 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_64
timestamp 0
transform 1 0 6992 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 0
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 0
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 0
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 0
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 0
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 0
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_155
timestamp 0
transform 1 0 15364 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_179
timestamp 0
transform 1 0 17572 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_191
timestamp 0
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 0
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 0
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 0
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 0
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 0
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_264
timestamp 0
transform 1 0 25392 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_268
timestamp 0
transform 1 0 25760 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_298
timestamp 0
transform 1 0 28520 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 0
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_318
timestamp 0
transform 1 0 30360 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_322
timestamp 0
transform 1 0 30728 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_339
timestamp 0
transform 1 0 32292 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_354
timestamp 0
transform 1 0 33672 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 0
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 0
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_377
timestamp 0
transform 1 0 35788 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_385
timestamp 0
transform 1 0 36524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 0
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_45
timestamp 0
transform 1 0 5244 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 0
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_66
timestamp 0
transform 1 0 7176 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_74
timestamp 0
transform 1 0 7912 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_79
timestamp 0
transform 1 0 8372 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_93
timestamp 0
transform 1 0 9660 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_106
timestamp 0
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_113
timestamp 0
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_134
timestamp 0
transform 1 0 13432 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_157
timestamp 0
transform 1 0 15548 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 0
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 0
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 0
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_191
timestamp 0
transform 1 0 18676 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_203
timestamp 0
transform 1 0 19780 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_215
timestamp 0
transform 1 0 20884 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 0
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 0
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 0
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 0
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 0
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_305
timestamp 0
transform 1 0 29164 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_313
timestamp 0
transform 1 0 29900 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_337
timestamp 0
transform 1 0 32108 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_360
timestamp 0
transform 1 0 34224 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_372
timestamp 0
transform 1 0 35328 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_384
timestamp 0
transform 1 0 36432 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 0
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 0
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 0
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_29
timestamp 0
transform 1 0 3772 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_33
timestamp 0
transform 1 0 4140 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 0
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 0
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 0
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_121
timestamp 0
transform 1 0 12236 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 0
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 0
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_153
timestamp 0
transform 1 0 15180 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_206
timestamp 0
transform 1 0 20056 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_218
timestamp 0
transform 1 0 21160 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_230
timestamp 0
transform 1 0 22264 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_242
timestamp 0
transform 1 0 23368 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 0
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_273
timestamp 0
transform 1 0 26220 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_290
timestamp 0
transform 1 0 27784 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_302
timestamp 0
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_338
timestamp 0
transform 1 0 32200 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 0
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_377
timestamp 0
transform 1 0 35788 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_385
timestamp 0
transform 1 0 36524 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 0
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 0
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 0
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 0
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 0
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 0
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 0
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_69
timestamp 0
transform 1 0 7452 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_75
timestamp 0
transform 1 0 8004 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_99
timestamp 0
transform 1 0 10212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 0
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 0
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_125
timestamp 0
transform 1 0 12604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 0
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 0
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_179
timestamp 0
transform 1 0 17572 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_183
timestamp 0
transform 1 0 17940 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 0
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 0
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_321
timestamp 0
transform 1 0 30636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_337
timestamp 0
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_368
timestamp 0
transform 1 0 34960 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_380
timestamp 0
transform 1 0 36064 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 0
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 0
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 0
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 0
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 0
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 0
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 0
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 0
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 0
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 0
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 0
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_109
timestamp 0
transform 1 0 11132 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_115
timestamp 0
transform 1 0 11684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 0
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_141
timestamp 0
transform 1 0 14076 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_174
timestamp 0
transform 1 0 17112 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_186
timestamp 0
transform 1 0 18216 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 0
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 0
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 0
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_233
timestamp 0
transform 1 0 22540 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 0
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_262
timestamp 0
transform 1 0 25208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_295
timestamp 0
transform 1 0 28244 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_316
timestamp 0
transform 1 0 30176 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 0
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_377
timestamp 0
transform 1 0 35788 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_385
timestamp 0
transform 1 0 36524 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 0
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 0
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 0
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 0
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 0
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 0
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 0
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 0
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 0
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 0
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 0
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 0
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 0
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_125
timestamp 0
transform 1 0 12604 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_148
timestamp 0
transform 1 0 14720 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_160
timestamp 0
transform 1 0 15824 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_178
timestamp 0
transform 1 0 17480 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_204
timestamp 0
transform 1 0 19872 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_208
timestamp 0
transform 1 0 20240 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 0
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_234
timestamp 0
transform 1 0 22632 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_246
timestamp 0
transform 1 0 23736 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_258
timestamp 0
transform 1 0 24840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 0
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_303
timestamp 0
transform 1 0 28980 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_323
timestamp 0
transform 1 0 30820 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 0
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 0
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_386
timestamp 0
transform 1 0 36616 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 0
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 0
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 0
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 0
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 0
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 0
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 0
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 0
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 0
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 0
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 0
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 0
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_121
timestamp 0
transform 1 0 12236 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_125
timestamp 0
transform 1 0 12604 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_135
timestamp 0
transform 1 0 13524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 0
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_141
timestamp 0
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_193
timestamp 0
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_206
timestamp 0
transform 1 0 20056 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_234
timestamp 0
transform 1 0 22632 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_238
timestamp 0
transform 1 0 23000 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 0
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_253
timestamp 0
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_261
timestamp 0
transform 1 0 25116 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_295
timestamp 0
transform 1 0 28244 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 0
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_313
timestamp 0
transform 1 0 29900 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_327
timestamp 0
transform 1 0 31188 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 0
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 0
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_377
timestamp 0
transform 1 0 35788 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_385
timestamp 0
transform 1 0 36524 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 0
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 0
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 0
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 0
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 0
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 0
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 0
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 0
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 0
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 0
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 0
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 0
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_133
timestamp 0
transform 1 0 13340 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_139
timestamp 0
transform 1 0 13892 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_160
timestamp 0
transform 1 0 15824 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_187
timestamp 0
transform 1 0 18308 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_199
timestamp 0
transform 1 0 19412 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 0
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_254
timestamp 0
transform 1 0 24472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 0
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 0
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_372
timestamp 0
transform 1 0 35328 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_384
timestamp 0
transform 1 0 36432 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 0
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 0
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 0
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 0
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 0
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 0
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 0
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 0
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 0
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 0
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 0
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_109
timestamp 0
transform 1 0 11132 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_115
timestamp 0
transform 1 0 11684 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 0
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 0
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_187
timestamp 0
transform 1 0 18308 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 0
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_197
timestamp 0
transform 1 0 19228 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_218
timestamp 0
transform 1 0 21160 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_242
timestamp 0
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 0
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 0
transform 1 0 26220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_277
timestamp 0
transform 1 0 26588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_298
timestamp 0
transform 1 0 28520 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_328
timestamp 0
transform 1 0 31280 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 0
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_379
timestamp 0
transform 1 0 35972 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_387
timestamp 0
transform 1 0 36708 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 0
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 0
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 0
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 0
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 0
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 0
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 0
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 0
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 0
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 0
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 0
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 0
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_113
timestamp 0
transform 1 0 11500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_135
timestamp 0
transform 1 0 13524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_141
timestamp 0
transform 1 0 14076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_162
timestamp 0
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_181
timestamp 0
transform 1 0 17756 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_189
timestamp 0
transform 1 0 18492 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_218
timestamp 0
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_59_225
timestamp 0
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 0
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 0
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_257
timestamp 0
transform 1 0 24748 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_269
timestamp 0
transform 1 0 25852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 0
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_281
timestamp 0
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 0
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_377
timestamp 0
transform 1 0 35788 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_385
timestamp 0
transform 1 0 36524 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 0
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 0
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 0
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 0
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 0
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 0
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 0
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 0
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 0
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 0
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 0
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_109
timestamp 0
transform 1 0 11132 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_137
timestamp 0
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 0
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_173
timestamp 0
transform 1 0 17020 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_206
timestamp 0
transform 1 0 20056 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_218
timestamp 0
transform 1 0 21160 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_230
timestamp 0
transform 1 0 22264 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 0
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 0
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 0
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_344
timestamp 0
transform 1 0 32752 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 0
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_381
timestamp 0
transform 1 0 36156 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_387
timestamp 0
transform 1 0 36708 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 0
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 0
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 0
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 0
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 0
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 0
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 0
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 0
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 0
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 0
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 0
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 0
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 0
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_125
timestamp 0
transform 1 0 12604 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_135
timestamp 0
transform 1 0 13524 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_147
timestamp 0
transform 1 0 14628 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 0
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_181
timestamp 0
transform 1 0 17756 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_185
timestamp 0
transform 1 0 18124 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_195
timestamp 0
transform 1 0 19044 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_207
timestamp 0
transform 1 0 20148 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_265
timestamp 0
transform 1 0 25484 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_281
timestamp 0
transform 1 0 26956 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_374
timestamp 0
transform 1 0 35512 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_386
timestamp 0
transform 1 0 36616 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 0
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 0
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 0
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 0
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 0
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 0
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 0
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 0
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 0
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 0
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 0
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_109
timestamp 0
transform 1 0 11132 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_132
timestamp 0
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_141
timestamp 0
transform 1 0 14076 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_151
timestamp 0
transform 1 0 14996 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_163
timestamp 0
transform 1 0 16100 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 0
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 0
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 0
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 0
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_253
timestamp 0
transform 1 0 24380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_273
timestamp 0
transform 1 0 26220 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_316
timestamp 0
transform 1 0 30176 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 0
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_369
timestamp 0
transform 1 0 35052 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_381
timestamp 0
transform 1 0 36156 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_387
timestamp 0
transform 1 0 36708 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 0
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 0
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 0
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 0
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 0
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 0
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 0
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 0
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 0
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 0
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 0
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 0
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_113
timestamp 0
transform 1 0 11500 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_178
timestamp 0
transform 1 0 17480 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_182
timestamp 0
transform 1 0 17848 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_212
timestamp 0
transform 1 0 20608 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 0
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_369
timestamp 0
transform 1 0 35052 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_381
timestamp 0
transform 1 0 36156 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_387
timestamp 0
transform 1 0 36708 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_19
timestamp 0
transform 1 0 2852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 0
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 0
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 0
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 0
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 0
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 0
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 0
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 0
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 0
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_109
timestamp 0
transform 1 0 11132 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_117
timestamp 0
transform 1 0 11868 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 0
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_141
timestamp 0
transform 1 0 14076 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_147
timestamp 0
transform 1 0 14628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_168
timestamp 0
transform 1 0 16560 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_174
timestamp 0
transform 1 0 17112 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 0
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_226
timestamp 0
transform 1 0 21896 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 0
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_309
timestamp 0
transform 1 0 29532 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_352
timestamp 0
transform 1 0 33488 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 0
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_377
timestamp 0
transform 1 0 35788 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_385
timestamp 0
transform 1 0 36524 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 0
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 0
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_27
timestamp 0
transform 1 0 3588 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_29
timestamp 0
transform 1 0 3772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_41
timestamp 0
transform 1 0 4876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_53
timestamp 0
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 0
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 0
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_81
timestamp 0
transform 1 0 8556 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_85
timestamp 0
transform 1 0 8924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_97
timestamp 0
transform 1 0 10028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_109
timestamp 0
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 0
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_125
timestamp 0
transform 1 0 12604 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_141
timestamp 0
transform 1 0 14076 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_153
timestamp 0
transform 1 0 15180 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_157
timestamp 0
transform 1 0 15548 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 0
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 0
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_181
timestamp 0
transform 1 0 17756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_185
timestamp 0
transform 1 0 18124 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_195
timestamp 0
transform 1 0 19044 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_197
timestamp 0
transform 1 0 19228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_209
timestamp 0
transform 1 0 20332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_221
timestamp 0
transform 1 0 21436 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 0
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_237
timestamp 0
transform 1 0 22908 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_249
timestamp 0
transform 1 0 24012 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_253
timestamp 0
transform 1 0 24380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_261
timestamp 0
transform 1 0 25116 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_265
timestamp 0
transform 1 0 25484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_277
timestamp 0
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_288
timestamp 0
transform 1 0 27600 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_296
timestamp 0
transform 1 0 28336 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_306
timestamp 0
transform 1 0 29256 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_309
timestamp 0
transform 1 0 29532 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_325
timestamp 0
transform 1 0 31004 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_329
timestamp 0
transform 1 0 31372 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 0
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_342
timestamp 0
transform 1 0 32568 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_354
timestamp 0
transform 1 0 33672 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_362
timestamp 0
transform 1 0 34408 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_365
timestamp 0
transform 1 0 34684 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_377
timestamp 0
transform 1 0 35788 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_385
timestamp 0
transform 1 0 36524 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 0
transform -1 0 36800 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 0
transform 1 0 29716 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 25484 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input5
timestamp 0
transform 1 0 1380 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  load_slew14
timestamp 0
transform 1 0 11684 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  load_slew15
timestamp 0
transform -1 0 3404 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  max_cap10
timestamp 0
transform -1 0 32292 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap11
timestamp 0
transform 1 0 32384 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap12
timestamp 0
transform -1 0 26864 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap13
timestamp 0
transform -1 0 31832 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 0
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 0
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 0
transform -1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_66
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 37076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_67
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 37076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_68
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 37076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_69
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 37076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_70
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 37076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_71
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 37076 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_72
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 37076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_73
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 37076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_74
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 37076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_75
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 37076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_76
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 37076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_77
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 37076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_78
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 37076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_79
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 37076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_80
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 37076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_81
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 37076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_82
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 37076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_83
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 37076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_84
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 37076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_85
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 37076 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_86
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 37076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_87
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 37076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_88
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 37076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_89
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 37076 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_90
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 37076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_91
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 37076 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_92
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 37076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_93
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 37076 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_94
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 37076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_95
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 37076 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_96
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 37076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_97
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 0
transform -1 0 37076 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_98
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 0
transform -1 0 37076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_99
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 0
transform -1 0 37076 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_100
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 0
transform -1 0 37076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_101
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 0
transform -1 0 37076 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_102
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 0
transform -1 0 37076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_103
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 0
transform -1 0 37076 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_104
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 0
transform -1 0 37076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_105
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 0
transform -1 0 37076 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_106
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 0
transform -1 0 37076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_107
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 0
transform -1 0 37076 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_108
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 0
transform -1 0 37076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_109
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 0
transform -1 0 37076 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_110
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 0
transform -1 0 37076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_111
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 0
transform -1 0 37076 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_112
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 0
transform -1 0 37076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_113
timestamp 0
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 0
transform -1 0 37076 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_114
timestamp 0
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 0
transform -1 0 37076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_115
timestamp 0
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 0
transform -1 0 37076 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_116
timestamp 0
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 0
transform -1 0 37076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_117
timestamp 0
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 0
transform -1 0 37076 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_118
timestamp 0
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 0
transform -1 0 37076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_119
timestamp 0
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 0
transform -1 0 37076 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_120
timestamp 0
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 0
transform -1 0 37076 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_121
timestamp 0
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 0
transform -1 0 37076 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_122
timestamp 0
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 0
transform -1 0 37076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_123
timestamp 0
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 0
transform -1 0 37076 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_124
timestamp 0
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 0
transform -1 0 37076 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_125
timestamp 0
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 0
transform -1 0 37076 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_126
timestamp 0
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 0
transform -1 0 37076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_127
timestamp 0
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 0
transform -1 0 37076 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_128
timestamp 0
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 0
transform -1 0 37076 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_129
timestamp 0
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 0
transform -1 0 37076 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_130
timestamp 0
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 0
transform -1 0 37076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_131
timestamp 0
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 0
transform -1 0 37076 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer4
timestamp 0
transform -1 0 35420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer5
timestamp 0
transform 1 0 33672 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_8  rebuffer6
timestamp 0
transform -1 0 32936 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer7
timestamp 0
transform -1 0 26864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  rebuffer8
timestamp 0
transform -1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer9
timestamp 0
transform -1 0 29256 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer10
timestamp 0
transform 1 0 31096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  rebuffer12
timestamp 0
transform -1 0 31648 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer13
timestamp 0
transform -1 0 31464 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  rebuffer14
timestamp 0
transform 1 0 30636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  rebuffer15
timestamp 0
transform 1 0 34684 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  rebuffer16
timestamp 0
transform -1 0 36156 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer17
timestamp 0
transform 1 0 33856 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__buf_8  rebuffer18
timestamp 0
transform -1 0 34408 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer19
timestamp 0
transform 1 0 29532 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  rebuffer20
timestamp 0
transform -1 0 29532 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  rebuffer21
timestamp 0
transform -1 0 29440 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  rebuffer22
timestamp 0
transform 1 0 28612 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer23
timestamp 0
transform -1 0 32660 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer25
timestamp 0
transform -1 0 32016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer26
timestamp 0
transform -1 0 35328 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  rebuffer27
timestamp 0
transform -1 0 35696 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  rebuffer28
timestamp 0
transform 1 0 30912 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer474
timestamp 0
transform -1 0 32752 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer475
timestamp 0
transform -1 0 32752 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer476
timestamp 0
transform 1 0 31004 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer477
timestamp 0
transform -1 0 30912 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer478
timestamp 0
transform 1 0 33580 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer479
timestamp 0
transform -1 0 31924 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer480
timestamp 0
transform 1 0 31372 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer481
timestamp 0
transform -1 0 33580 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer483
timestamp 0
transform 1 0 30636 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer484
timestamp 0
transform 1 0 29256 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer485
timestamp 0
transform -1 0 26864 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer486
timestamp 0
transform 1 0 28612 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer487
timestamp 0
transform -1 0 29256 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer488
timestamp 0
transform 1 0 30176 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer489
timestamp 0
transform -1 0 30176 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer490
timestamp 0
transform 1 0 29532 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer492
timestamp 0
transform -1 0 35052 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  rebuffer493
timestamp 0
transform -1 0 35420 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  rebuffer625
timestamp 0
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  rebuffer628
timestamp 0
transform -1 0 33120 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  rebuffer629
timestamp 0
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer713
timestamp 0
transform -1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  rebuffer715
timestamp 0
transform -1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  rebuffer717
timestamp 0
transform -1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer720
timestamp 0
transform 1 0 29992 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  rebuffer721
timestamp 0
transform -1 0 31280 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  rebuffer723
timestamp 0
transform -1 0 30912 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer794
timestamp 0
transform -1 0 29900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer795
timestamp 0
transform 1 0 30820 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  rebuffer798
timestamp 0
transform 1 0 34224 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer800
timestamp 0
transform 1 0 33580 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  rebuffer802
timestamp 0
transform 1 0 34040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer804
timestamp 0
transform 1 0 31004 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  rebuffer805
timestamp 0
transform -1 0 35512 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer830
timestamp 0
transform -1 0 33304 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer832
timestamp 0
transform -1 0 33304 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  split1
timestamp 0
transform 1 0 35696 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  split3
timestamp 0
transform -1 0 33856 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  split11
timestamp 0
transform 1 0 32384 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  Systolic4x4_serial_io_16
timestamp 0
transform 1 0 36524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 0
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 0
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_144
timestamp 0
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_145
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_146
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_147
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_148
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_149
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_150
timestamp 0
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_151
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_152
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_153
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_154
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_155
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_156
timestamp 0
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_157
timestamp 0
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_158
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_159
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_160
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_161
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_162
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_163
timestamp 0
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_164
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_165
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_166
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_167
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_168
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_169
timestamp 0
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_170
timestamp 0
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_171
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_172
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_173
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_174
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_175
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_176
timestamp 0
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_177
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_178
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_179
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_180
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_181
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_182
timestamp 0
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_183
timestamp 0
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_184
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_185
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_186
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_187
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_188
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_189
timestamp 0
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_190
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_191
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_192
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_193
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_194
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_195
timestamp 0
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_196
timestamp 0
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_197
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_198
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_199
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_200
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_201
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_202
timestamp 0
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_203
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_204
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_205
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_206
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_207
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_208
timestamp 0
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_209
timestamp 0
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_210
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_211
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_212
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_213
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_214
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_215
timestamp 0
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_216
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_217
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_218
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_219
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_220
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_221
timestamp 0
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_222
timestamp 0
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_223
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_224
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_225
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_226
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_227
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_228
timestamp 0
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_229
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_230
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_231
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_232
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_233
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_234
timestamp 0
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_235
timestamp 0
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_236
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_237
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_238
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_239
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_240
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_241
timestamp 0
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_242
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_243
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_244
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_245
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_246
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_247
timestamp 0
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_248
timestamp 0
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_249
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_250
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_251
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_252
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_253
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_254
timestamp 0
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_255
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_256
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_257
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_258
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_259
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_260
timestamp 0
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_261
timestamp 0
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_262
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_263
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_264
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_265
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_266
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_267
timestamp 0
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_268
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_269
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_270
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_271
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_272
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_273
timestamp 0
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_274
timestamp 0
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_275
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_276
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_277
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_278
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_279
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_280
timestamp 0
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_281
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_282
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_283
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_284
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_285
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_286
timestamp 0
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_287
timestamp 0
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_288
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_289
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_290
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_291
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_292
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_293
timestamp 0
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_294
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_295
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_296
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_297
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_298
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_299
timestamp 0
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_300
timestamp 0
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_301
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_302
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_303
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_304
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_305
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_306
timestamp 0
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_307
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_308
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_309
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_310
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_311
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_312
timestamp 0
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_313
timestamp 0
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_314
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_315
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_316
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_317
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_318
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_319
timestamp 0
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_320
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_321
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_322
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_323
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_324
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_325
timestamp 0
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_326
timestamp 0
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_327
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_328
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_329
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_330
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_331
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_332
timestamp 0
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_333
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_334
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_335
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_336
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_337
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_338
timestamp 0
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_339
timestamp 0
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_340
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_341
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_342
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_343
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_344
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_345
timestamp 0
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_346
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_347
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_348
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_349
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_350
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_351
timestamp 0
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_352
timestamp 0
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_353
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_354
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_355
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_356
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_357
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_358
timestamp 0
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_359
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_360
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_361
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_362
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_363
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_364
timestamp 0
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_365
timestamp 0
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_366
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_367
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_368
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_369
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_370
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_371
timestamp 0
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_372
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_373
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_374
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_375
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_376
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_377
timestamp 0
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_378
timestamp 0
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_379
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_380
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_381
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_382
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_383
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_384
timestamp 0
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_385
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_386
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_387
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_388
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_389
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_390
timestamp 0
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_391
timestamp 0
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_392
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_393
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_394
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_395
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_396
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_397
timestamp 0
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_398
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_399
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_400
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_401
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_402
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_403
timestamp 0
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_404
timestamp 0
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_405
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_406
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_407
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_408
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_409
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_410
timestamp 0
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_411
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_412
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_413
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_414
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_415
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_416
timestamp 0
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_417
timestamp 0
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_418
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_419
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_420
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_421
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_422
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_423
timestamp 0
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_424
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_425
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_426
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_427
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_428
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_429
timestamp 0
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_430
timestamp 0
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_431
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_432
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_433
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_434
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_435
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_436
timestamp 0
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_437
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_438
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_439
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_440
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_441
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_442
timestamp 0
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_443
timestamp 0
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_444
timestamp 0
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_445
timestamp 0
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_446
timestamp 0
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_447
timestamp 0
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_448
timestamp 0
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_449
timestamp 0
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_450
timestamp 0
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_451
timestamp 0
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_452
timestamp 0
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_453
timestamp 0
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_454
timestamp 0
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_455
timestamp 0
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_456
timestamp 0
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_457
timestamp 0
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_458
timestamp 0
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_459
timestamp 0
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_460
timestamp 0
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_461
timestamp 0
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_462
timestamp 0
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_463
timestamp 0
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_464
timestamp 0
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_465
timestamp 0
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_466
timestamp 0
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_467
timestamp 0
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_468
timestamp 0
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_469
timestamp 0
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_470
timestamp 0
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_471
timestamp 0
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_472
timestamp 0
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_473
timestamp 0
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_474
timestamp 0
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_475
timestamp 0
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_476
timestamp 0
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_477
timestamp 0
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_478
timestamp 0
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_479
timestamp 0
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_480
timestamp 0
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_481
timestamp 0
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_482
timestamp 0
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_483
timestamp 0
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_484
timestamp 0
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_485
timestamp 0
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_486
timestamp 0
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_487
timestamp 0
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_488
timestamp 0
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_489
timestamp 0
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_490
timestamp 0
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_491
timestamp 0
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_492
timestamp 0
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_493
timestamp 0
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_494
timestamp 0
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_495
timestamp 0
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_496
timestamp 0
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_497
timestamp 0
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_498
timestamp 0
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_499
timestamp 0
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_500
timestamp 0
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_501
timestamp 0
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_502
timestamp 0
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_503
timestamp 0
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_504
timestamp 0
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_505
timestamp 0
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_506
timestamp 0
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_507
timestamp 0
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_508
timestamp 0
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_509
timestamp 0
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_510
timestamp 0
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_511
timestamp 0
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_512
timestamp 0
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_513
timestamp 0
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_514
timestamp 0
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_515
timestamp 0
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_516
timestamp 0
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_517
timestamp 0
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_518
timestamp 0
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_519
timestamp 0
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_520
timestamp 0
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_521
timestamp 0
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_522
timestamp 0
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_523
timestamp 0
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_524
timestamp 0
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_525
timestamp 0
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_526
timestamp 0
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_527
timestamp 0
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_528
timestamp 0
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_529
timestamp 0
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_530
timestamp 0
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_531
timestamp 0
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_532
timestamp 0
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_533
timestamp 0
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_534
timestamp 0
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_535
timestamp 0
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_536
timestamp 0
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_537
timestamp 0
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_538
timestamp 0
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_539
timestamp 0
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_540
timestamp 0
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_541
timestamp 0
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_542
timestamp 0
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_543
timestamp 0
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_544
timestamp 0
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_545
timestamp 0
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_546
timestamp 0
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_547
timestamp 0
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_548
timestamp 0
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_549
timestamp 0
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_550
timestamp 0
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_551
timestamp 0
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_552
timestamp 0
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_553
timestamp 0
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_554
timestamp 0
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_555
timestamp 0
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_556
timestamp 0
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_557
timestamp 0
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_558
timestamp 0
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_559
timestamp 0
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_560
timestamp 0
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_561
timestamp 0
transform 1 0 3680 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_562
timestamp 0
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_563
timestamp 0
transform 1 0 8832 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_564
timestamp 0
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_565
timestamp 0
transform 1 0 13984 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_566
timestamp 0
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_567
timestamp 0
transform 1 0 19136 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_568
timestamp 0
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_569
timestamp 0
transform 1 0 24288 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_570
timestamp 0
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_571
timestamp 0
transform 1 0 29440 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_572
timestamp 0
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_573
timestamp 0
transform 1 0 34592 0 -1 38080
box -38 -48 130 592
<< labels >>
rlabel metal1 s 19090 38080 19090 38080 4 VGND
rlabel metal1 s 19090 37536 19090 37536 4 VPWR
rlabel metal2 s 36662 16439 36662 16439 4 A_in_frame_sync
rlabel metal1 s 22218 12240 22218 12240 4 A_in_serial_clk
rlabel metal2 s 23230 1588 23230 1588 4 A_in_serial_data
rlabel metal2 s 29762 38743 29762 38743 4 B_in_frame_sync
rlabel metal1 s 28566 30158 28566 30158 4 B_in_serial_clk
rlabel metal2 s 25254 38743 25254 38743 4 B_in_serial_data
rlabel metal1 s 1380 14042 1380 14042 4 C_out_frame_sync
rlabel metal3 s 1050 17748 1050 17748 4 C_out_serial_clk
rlabel metal1 s 31648 6834 31648 6834 4 _0000_
rlabel metal1 s 30360 31858 30360 31858 4 _0001_
rlabel metal1 s 5198 16490 5198 16490 4 _0002_
rlabel metal1 s 2070 25228 2070 25228 4 _0003_
rlabel metal2 s 1886 24616 1886 24616 4 _0004_
rlabel metal1 s 1840 26554 1840 26554 4 _0005_
rlabel metal2 s 2155 27642 2155 27642 4 _0006_
rlabel metal1 s 1886 28730 1886 28730 4 _0007_
rlabel metal1 s 3726 29716 3726 29716 4 _0008_
rlabel metal2 s 3818 29988 3818 29988 4 _0009_
rlabel metal2 s 5566 29410 5566 29410 4 _0010_
rlabel metal2 s 6394 30498 6394 30498 4 _0011_
rlabel metal1 s 6164 26758 6164 26758 4 _0012_
rlabel metal2 s 7130 24548 7130 24548 4 _0013_
rlabel metal1 s 4547 26554 4547 26554 4 _0014_
rlabel metal2 s 4370 25058 4370 25058 4 _0015_
rlabel metal2 s 5290 23324 5290 23324 4 _0016_
rlabel metal2 s 1695 22202 1695 22202 4 _0017_
rlabel metal2 s 3450 22814 3450 22814 4 _0018_
rlabel metal2 s 3450 21284 3450 21284 4 _0019_
rlabel metal2 s 6118 21148 6118 21148 4 _0020_
rlabel metal2 s 6670 20638 6670 20638 4 _0021_
rlabel metal2 s 9706 19788 9706 19788 4 _0022_
rlabel metal1 s 7544 18802 7544 18802 4 _0023_
rlabel metal1 s 10626 20026 10626 20026 4 _0024_
rlabel metal2 s 10350 21148 10350 21148 4 _0025_
rlabel metal1 s 10708 22202 10708 22202 4 _0026_
rlabel metal2 s 10074 22882 10074 22882 4 _0027_
rlabel metal1 s 7774 22746 7774 22746 4 _0028_
rlabel metal2 s 9246 26146 9246 26146 4 _0029_
rlabel metal1 s 10764 25466 10764 25466 4 _0030_
rlabel metal2 s 10902 27098 10902 27098 4 _0031_
rlabel metal1 s 9292 27642 9292 27642 4 _0032_
rlabel metal1 s 7866 28730 7866 28730 4 _0033_
rlabel metal2 s 8326 30328 8326 30328 4 _0034_
rlabel metal2 s 8970 31076 8970 31076 4 _0035_
rlabel metal2 s 9982 29852 9982 29852 4 _0036_
rlabel metal1 s 30360 5882 30360 5882 4 _0037_
rlabel metal1 s 30498 3570 30498 3570 4 _0038_
rlabel metal1 s 29578 4522 29578 4522 4 _0039_
rlabel metal2 s 30498 3502 30498 3502 4 _0040_
rlabel metal2 s 32430 3230 32430 3230 4 _0041_
rlabel metal1 s 35236 4182 35236 4182 4 _0042_
rlabel metal1 s 34270 6392 34270 6392 4 _0043_
rlabel metal2 s 32614 6528 32614 6528 4 _0044_
rlabel metal2 s 28474 7582 28474 7582 4 _0045_
rlabel metal1 s 29808 8534 29808 8534 4 _0046_
rlabel metal1 s 29532 10234 29532 10234 4 _0047_
rlabel metal2 s 30409 10778 30409 10778 4 _0048_
rlabel metal1 s 31408 11322 31408 11322 4 _0049_
rlabel metal1 s 33911 9146 33911 9146 4 _0050_
rlabel metal1 s 34914 10234 34914 10234 4 _0051_
rlabel metal1 s 32982 10744 32982 10744 4 _0052_
rlabel metal1 s 27232 5270 27232 5270 4 _0053_
rlabel metal1 s 26765 5882 26765 5882 4 _0054_
rlabel metal1 s 26673 6970 26673 6970 4 _0055_
rlabel metal2 s 28014 8024 28014 8024 4 _0056_
rlabel metal1 s 28060 9010 28060 9010 4 _0057_
rlabel metal1 s 27048 9622 27048 9622 4 _0058_
rlabel metal1 s 27692 12614 27692 12614 4 _0059_
rlabel metal1 s 27376 11322 27376 11322 4 _0060_
rlabel metal1 s 28428 11662 28428 11662 4 _0061_
rlabel metal1 s 30176 12886 30176 12886 4 _0062_
rlabel metal1 s 31234 12750 31234 12750 4 _0063_
rlabel metal2 s 32154 13056 32154 13056 4 _0064_
rlabel metal2 s 33902 13464 33902 13464 4 _0065_
rlabel metal1 s 34500 12138 34500 12138 4 _0066_
rlabel metal1 s 34261 13158 34261 13158 4 _0067_
rlabel metal2 s 34730 14688 34730 14688 4 _0068_
rlabel metal1 s 32982 13974 32982 13974 4 _0069_
rlabel metal2 s 32062 15028 32062 15028 4 _0070_
rlabel metal2 s 31418 14926 31418 14926 4 _0071_
rlabel metal2 s 32246 15708 32246 15708 4 _0072_
rlabel metal2 s 28934 15844 28934 15844 4 _0073_
rlabel metal2 s 27830 16796 27830 16796 4 _0074_
rlabel metal1 s 27508 15062 27508 15062 4 _0075_
rlabel metal1 s 26772 14042 26772 14042 4 _0076_
rlabel metal1 s 25392 13974 25392 13974 4 _0077_
rlabel metal1 s 24564 13362 24564 13362 4 _0078_
rlabel metal1 s 24288 12750 24288 12750 4 _0079_
rlabel metal1 s 23000 11798 23000 11798 4 _0080_
rlabel metal2 s 24702 11492 24702 11492 4 _0081_
rlabel metal2 s 24702 10268 24702 10268 4 _0082_
rlabel metal1 s 25116 9146 25116 9146 4 _0083_
rlabel metal1 s 24840 7786 24840 7786 4 _0084_
rlabel metal2 s 24610 8160 24610 8160 4 _0085_
rlabel metal1 s 24012 7446 24012 7446 4 _0086_
rlabel metal1 s 23414 7956 23414 7956 4 _0087_
rlabel metal1 s 22586 9010 22586 9010 4 _0088_
rlabel metal2 s 23230 10336 23230 10336 4 _0089_
rlabel metal2 s 22218 10608 22218 10608 4 _0090_
rlabel metal1 s 21797 12410 21797 12410 4 _0091_
rlabel metal1 s 21482 13838 21482 13838 4 _0092_
rlabel metal1 s 20470 15096 20470 15096 4 _0093_
rlabel metal1 s 19826 16966 19826 16966 4 _0094_
rlabel metal2 s 21942 16796 21942 16796 4 _0095_
rlabel metal2 s 20930 18224 20930 18224 4 _0096_
rlabel metal1 s 20056 18326 20056 18326 4 _0097_
rlabel metal1 s 20010 19414 20010 19414 4 _0098_
rlabel metal1 s 20424 20366 20424 20366 4 _0099_
rlabel metal2 s 22126 20672 22126 20672 4 _0100_
rlabel metal1 s 24426 20808 24426 20808 4 _0101_
rlabel metal1 s 22954 19482 22954 19482 4 _0102_
rlabel metal1 s 23000 17850 23000 17850 4 _0103_
rlabel metal1 s 25438 18632 25438 18632 4 _0104_
rlabel metal1 s 26312 17578 26312 17578 4 _0105_
rlabel metal1 s 26588 19414 26588 19414 4 _0106_
rlabel metal2 s 25070 19992 25070 19992 4 _0107_
rlabel metal2 s 27738 20128 27738 20128 4 _0108_
rlabel metal2 s 27646 21148 27646 21148 4 _0109_
rlabel metal2 s 31050 21148 31050 21148 4 _0110_
rlabel metal1 s 31188 20502 31188 20502 4 _0111_
rlabel metal2 s 32982 21080 32982 21080 4 _0112_
rlabel metal1 s 33442 20842 33442 20842 4 _0113_
rlabel metal1 s 35098 20502 35098 20502 4 _0114_
rlabel metal2 s 34730 19516 34730 19516 4 _0115_
rlabel metal2 s 35374 18632 35374 18632 4 _0116_
rlabel metal2 s 33350 18326 33350 18326 4 _0117_
rlabel metal1 s 34132 16218 34132 16218 4 _0118_
rlabel metal2 s 32430 16864 32430 16864 4 _0119_
rlabel metal2 s 31786 17714 31786 17714 4 _0120_
rlabel metal1 s 30452 17578 30452 17578 4 _0121_
rlabel metal1 s 30130 18802 30130 18802 4 _0122_
rlabel metal1 s 27830 18632 27830 18632 4 _0123_
rlabel metal1 s 27462 18190 27462 18190 4 _0124_
rlabel metal1 s 26082 17102 26082 17102 4 _0125_
rlabel metal2 s 25714 16354 25714 16354 4 _0126_
rlabel metal2 s 24426 15776 24426 15776 4 _0127_
rlabel metal2 s 22678 16320 22678 16320 4 _0128_
rlabel metal1 s 22540 15130 22540 15130 4 _0129_
rlabel metal1 s 22862 13974 22862 13974 4 _0130_
rlabel metal1 s 21482 12818 21482 12818 4 _0131_
rlabel metal1 s 19458 12750 19458 12750 4 _0132_
rlabel metal2 s 19366 10846 19366 10846 4 _0133_
rlabel metal1 s 19320 10098 19320 10098 4 _0134_
rlabel metal1 s 20240 9622 20240 9622 4 _0135_
rlabel metal2 s 18814 8160 18814 8160 4 _0136_
rlabel metal2 s 18538 6800 18538 6800 4 _0137_
rlabel metal1 s 17158 6358 17158 6358 4 _0138_
rlabel metal1 s 16928 5270 16928 5270 4 _0139_
rlabel metal2 s 15594 5134 15594 5134 4 _0140_
rlabel metal2 s 14398 5440 14398 5440 4 _0141_
rlabel metal1 s 14904 6698 14904 6698 4 _0142_
rlabel metal1 s 14812 7446 14812 7446 4 _0143_
rlabel metal1 s 14444 8874 14444 8874 4 _0144_
rlabel metal1 s 14352 9962 14352 9962 4 _0145_
rlabel metal1 s 14812 10574 14812 10574 4 _0146_
rlabel metal1 s 14996 11662 14996 11662 4 _0147_
rlabel metal1 s 14950 12750 14950 12750 4 _0148_
rlabel metal1 s 14858 13362 14858 13362 4 _0149_
rlabel metal2 s 15594 14620 15594 14620 4 _0150_
rlabel metal2 s 14398 15776 14398 15776 4 _0151_
rlabel metal1 s 15180 16626 15180 16626 4 _0152_
rlabel metal1 s 14950 17578 14950 17578 4 _0153_
rlabel metal2 s 14950 18462 14950 18462 4 _0154_
rlabel metal2 s 15042 19040 15042 19040 4 _0155_
rlabel metal1 s 14904 20366 14904 20366 4 _0156_
rlabel metal1 s 16652 19414 16652 19414 4 _0157_
rlabel metal1 s 17342 20502 17342 20502 4 _0158_
rlabel metal1 s 17894 19278 17894 19278 4 _0159_
rlabel metal1 s 17655 18394 17655 18394 4 _0160_
rlabel metal1 s 18308 17306 18308 17306 4 _0161_
rlabel metal1 s 17480 17102 17480 17102 4 _0162_
rlabel metal2 s 18814 15776 18814 15776 4 _0163_
rlabel metal2 s 17618 14484 17618 14484 4 _0164_
rlabel metal2 s 18446 14144 18446 14144 4 _0165_
rlabel metal1 s 17296 11798 17296 11798 4 _0166_
rlabel metal1 s 18124 10710 18124 10710 4 _0167_
rlabel metal1 s 18124 9622 18124 9622 4 _0168_
rlabel metal1 s 17296 10098 17296 10098 4 _0169_
rlabel metal1 s 17756 8874 17756 8874 4 _0170_
rlabel metal2 s 21206 8670 21206 8670 4 _0171_
rlabel metal2 s 22218 7344 22218 7344 4 _0172_
rlabel metal1 s 21068 6358 21068 6358 4 _0173_
rlabel metal2 s 19550 6222 19550 6222 4 _0174_
rlabel metal2 s 20838 4896 20838 4896 4 _0175_
rlabel metal2 s 23322 5678 23322 5678 4 _0176_
rlabel metal1 s 23046 5610 23046 5610 4 _0177_
rlabel metal2 s 24426 4896 24426 4896 4 _0178_
rlabel metal2 s 24426 5984 24426 5984 4 _0179_
rlabel metal1 s 28060 35054 28060 35054 4 _0180_
rlabel metal2 s 27738 37230 27738 37230 4 _0181_
rlabel metal1 s 27600 35734 27600 35734 4 _0182_
rlabel metal2 s 28566 33558 28566 33558 4 _0183_
rlabel metal1 s 27784 32334 27784 32334 4 _0184_
rlabel metal1 s 29900 35734 29900 35734 4 _0185_
rlabel metal1 s 29808 33422 29808 33422 4 _0186_
rlabel metal2 s 30314 31518 30314 31518 4 _0187_
rlabel metal1 s 30406 36210 30406 36210 4 _0188_
rlabel metal1 s 31786 37162 31786 37162 4 _0189_
rlabel metal2 s 33534 36516 33534 36516 4 _0190_
rlabel metal1 s 33810 35598 33810 35598 4 _0191_
rlabel metal1 s 34040 34510 34040 34510 4 _0192_
rlabel metal2 s 34454 33728 34454 33728 4 _0193_
rlabel metal1 s 33948 32334 33948 32334 4 _0194_
rlabel metal1 s 32384 31450 32384 31450 4 _0195_
rlabel metal1 s 34132 8534 34132 8534 4 _0196_
rlabel metal1 s 24840 34986 24840 34986 4 _0197_
rlabel metal1 s 24886 34034 24886 34034 4 _0198_
rlabel metal1 s 25070 33082 25070 33082 4 _0199_
rlabel metal1 s 27186 31858 27186 31858 4 _0200_
rlabel metal1 s 27140 30906 27140 30906 4 _0201_
rlabel metal1 s 27462 29716 27462 29716 4 _0202_
rlabel metal2 s 27278 28900 27278 28900 4 _0203_
rlabel metal1 s 29946 28730 29946 28730 4 _0204_
rlabel metal1 s 29624 28118 29624 28118 4 _0205_
rlabel metal1 s 31234 28594 31234 28594 4 _0206_
rlabel metal1 s 31004 30158 31004 30158 4 _0207_
rlabel metal1 s 34224 30294 34224 30294 4 _0208_
rlabel metal2 s 32522 29342 32522 29342 4 _0209_
rlabel metal2 s 32706 28288 32706 28288 4 _0210_
rlabel metal2 s 33258 27370 33258 27370 4 _0211_
rlabel metal1 s 32706 26214 32706 26214 4 _0212_
rlabel metal2 s 33350 24956 33350 24956 4 _0213_
rlabel metal1 s 33718 23834 33718 23834 4 _0214_
rlabel metal1 s 33120 23018 33120 23018 4 _0215_
rlabel metal2 s 32430 23154 32430 23154 4 _0216_
rlabel metal1 s 31280 24310 31280 24310 4 _0217_
rlabel metal1 s 30360 24242 30360 24242 4 _0218_
rlabel metal2 s 29394 24480 29394 24480 4 _0219_
rlabel metal1 s 27738 25806 27738 25806 4 _0220_
rlabel metal1 s 26772 23834 26772 23834 4 _0221_
rlabel metal1 s 25300 23834 25300 23834 4 _0222_
rlabel metal1 s 24886 24242 24886 24242 4 _0223_
rlabel metal2 s 23966 24242 23966 24242 4 _0224_
rlabel metal1 s 22218 25194 22218 25194 4 _0225_
rlabel metal2 s 20838 24718 20838 24718 4 _0226_
rlabel metal2 s 22126 27098 22126 27098 4 _0227_
rlabel metal1 s 21574 26486 21574 26486 4 _0228_
rlabel metal2 s 22862 26724 22862 26724 4 _0229_
rlabel metal2 s 25346 27166 25346 27166 4 _0230_
rlabel metal2 s 25898 27132 25898 27132 4 _0231_
rlabel metal1 s 25070 25738 25070 25738 4 _0232_
rlabel metal1 s 28336 27030 28336 27030 4 _0233_
rlabel metal2 s 28474 26860 28474 26860 4 _0234_
rlabel metal2 s 30682 27438 30682 27438 4 _0235_
rlabel metal2 s 32154 27336 32154 27336 4 _0236_
rlabel metal1 s 30084 25942 30084 25942 4 _0237_
rlabel metal2 s 30222 23392 30222 23392 4 _0238_
rlabel metal1 s 29440 22066 29440 22066 4 _0239_
rlabel metal2 s 27915 22202 27915 22202 4 _0240_
rlabel metal2 s 27278 22848 27278 22848 4 _0241_
rlabel metal1 s 25530 22984 25530 22984 4 _0242_
rlabel metal1 s 24879 22202 24879 22202 4 _0243_
rlabel metal1 s 24150 21998 24150 21998 4 _0244_
rlabel metal2 s 22218 22814 22218 22814 4 _0245_
rlabel metal1 s 21107 22202 21107 22202 4 _0246_
rlabel metal2 s 20010 22848 20010 22848 4 _0247_
rlabel metal2 s 18078 22848 18078 22848 4 _0248_
rlabel metal1 s 19642 24106 19642 24106 4 _0249_
rlabel metal1 s 19596 24718 19596 24718 4 _0250_
rlabel metal2 s 17986 26350 17986 26350 4 _0251_
rlabel metal2 s 17250 26044 17250 26044 4 _0252_
rlabel metal2 s 17434 26146 17434 26146 4 _0253_
rlabel metal1 s 15456 24922 15456 24922 4 _0254_
rlabel metal1 s 15134 23834 15134 23834 4 _0255_
rlabel metal2 s 17802 23970 17802 23970 4 _0256_
rlabel metal1 s 16783 22202 16783 22202 4 _0257_
rlabel metal2 s 15594 22610 15594 22610 4 _0258_
rlabel metal1 s 14490 22202 14490 22202 4 _0259_
rlabel metal1 s 13294 22542 13294 22542 4 _0260_
rlabel metal2 s 12466 23324 12466 23324 4 _0261_
rlabel metal1 s 12788 24242 12788 24242 4 _0262_
rlabel metal1 s 13103 25466 13103 25466 4 _0263_
rlabel metal1 s 13616 25806 13616 25806 4 _0264_
rlabel metal1 s 14720 27098 14720 27098 4 _0265_
rlabel metal1 s 12742 26554 12742 26554 4 _0266_
rlabel metal2 s 12006 28254 12006 28254 4 _0267_
rlabel metal2 s 11822 29410 11822 29410 4 _0268_
rlabel metal2 s 12650 30362 12650 30362 4 _0269_
rlabel metal1 s 15272 29818 15272 29818 4 _0270_
rlabel metal1 s 14536 28730 14536 28730 4 _0271_
rlabel metal1 s 17342 29274 17342 29274 4 _0272_
rlabel metal2 s 16330 27778 16330 27778 4 _0273_
rlabel metal1 s 18216 27642 18216 27642 4 _0274_
rlabel metal2 s 18814 28764 18814 28764 4 _0275_
rlabel metal2 s 19543 27642 19543 27642 4 _0276_
rlabel metal1 s 19642 29274 19642 29274 4 _0277_
rlabel metal2 s 20746 28764 20746 28764 4 _0278_
rlabel metal1 s 23184 28730 23184 28730 4 _0279_
rlabel metal1 s 23782 28730 23782 28730 4 _0280_
rlabel metal2 s 25162 29376 25162 29376 4 _0281_
rlabel metal2 s 25898 29308 25898 29308 4 _0282_
rlabel metal1 s 25300 30770 25300 30770 4 _0283_
rlabel metal1 s 24380 31382 24380 31382 4 _0284_
rlabel metal1 s 22540 31382 22540 31382 4 _0285_
rlabel metal1 s 23046 33082 23046 33082 4 _0286_
rlabel metal2 s 22126 34136 22126 34136 4 _0287_
rlabel metal2 s 21114 33116 21114 33116 4 _0288_
rlabel metal2 s 21022 32028 21022 32028 4 _0289_
rlabel metal1 s 20286 30906 20286 30906 4 _0290_
rlabel metal1 s 18814 30906 18814 30906 4 _0291_
rlabel metal1 s 17756 30362 17756 30362 4 _0292_
rlabel metal1 s 15916 30634 15916 30634 4 _0293_
rlabel metal2 s 15594 32028 15594 32028 4 _0294_
rlabel metal2 s 14490 31518 14490 31518 4 _0295_
rlabel metal1 s 13294 31450 13294 31450 4 _0296_
rlabel metal2 s 12098 32300 12098 32300 4 _0297_
rlabel metal1 s 11822 33592 11822 33592 4 _0298_
rlabel metal2 s 12098 34204 12098 34204 4 _0299_
rlabel metal2 s 13386 35224 13386 35224 4 _0300_
rlabel metal2 s 11730 36380 11730 36380 4 _0301_
rlabel metal2 s 13478 37468 13478 37468 4 _0302_
rlabel metal1 s 14306 36346 14306 36346 4 _0303_
rlabel metal2 s 16238 37468 16238 37468 4 _0304_
rlabel metal1 s 16629 36618 16629 36618 4 _0305_
rlabel metal2 s 15502 35224 15502 35224 4 _0306_
rlabel metal1 s 16629 34510 16629 34510 4 _0307_
rlabel metal2 s 14306 33864 14306 33864 4 _0308_
rlabel metal2 s 15962 33762 15962 33762 4 _0309_
rlabel metal2 s 18538 33116 18538 33116 4 _0310_
rlabel metal2 s 19550 32606 19550 32606 4 _0311_
rlabel metal2 s 19734 33762 19734 33762 4 _0312_
rlabel metal1 s 19136 34510 19136 34510 4 _0313_
rlabel metal2 s 17618 35292 17618 35292 4 _0314_
rlabel metal2 s 17526 36380 17526 36380 4 _0315_
rlabel metal2 s 17526 37468 17526 37468 4 _0316_
rlabel metal1 s 20102 36686 20102 36686 4 _0317_
rlabel metal2 s 21482 36890 21482 36890 4 _0318_
rlabel metal1 s 20608 36210 20608 36210 4 _0319_
rlabel metal1 s 23506 36686 23506 36686 4 _0320_
rlabel metal1 s 25208 35734 25208 35734 4 _0321_
rlabel metal2 s 22402 37468 22402 37468 4 _0322_
rlabel metal1 s 25990 36890 25990 36890 4 _0323_
rlabel metal1 s 26680 36890 26680 36890 4 _0324_
rlabel metal1 s 30176 5338 30176 5338 4 _0325_
rlabel metal2 s 1886 13906 1886 13906 4 _0326_
rlabel metal2 s 4462 14110 4462 14110 4 _0327_
rlabel metal2 s 1702 15708 1702 15708 4 _0328_
rlabel metal1 s 1886 16762 1886 16762 4 _0329_
rlabel metal2 s 4370 17374 4370 17374 4 _0330_
rlabel metal1 s 5888 18802 5888 18802 4 _0331_
rlabel metal1 s 5106 19278 5106 19278 4 _0332_
rlabel metal1 s 1794 20366 1794 20366 4 _0333_
rlabel metal2 s 2346 19482 2346 19482 4 _0334_
rlabel metal1 s 1794 18190 1794 18190 4 _0335_
rlabel metal1 s 30123 30906 30123 30906 4 _0336_
rlabel metal2 s 5290 14620 5290 14620 4 _0337_
rlabel metal1 s 6338 13702 6338 13702 4 _0338_
rlabel metal2 s 7222 15708 7222 15708 4 _0339_
rlabel metal1 s 8970 13974 8970 13974 4 _0340_
rlabel metal1 s 9982 14314 9982 14314 4 _0341_
rlabel metal2 s 10902 15708 10902 15708 4 _0342_
rlabel metal2 s 10902 16796 10902 16796 4 _0343_
rlabel metal1 s 10074 17850 10074 17850 4 _0344_
rlabel metal1 s 8188 16762 8188 16762 4 _0345_
rlabel metal2 s 6578 17442 6578 17442 4 _0346_
rlabel metal1 s 31970 35802 31970 35802 4 _0347_
rlabel metal1 s 31234 33966 31234 33966 4 _0348_
rlabel metal2 s 27094 36142 27094 36142 4 _0349_
rlabel metal2 s 27278 36108 27278 36108 4 _0350_
rlabel metal2 s 28106 37638 28106 37638 4 _0351_
rlabel metal2 s 28934 33694 28934 33694 4 _0352_
rlabel metal2 s 29026 33116 29026 33116 4 _0353_
rlabel metal1 s 28934 33422 28934 33422 4 _0354_
rlabel metal1 s 28244 33490 28244 33490 4 _0355_
rlabel metal1 s 31418 35530 31418 35530 4 _0356_
rlabel metal1 s 30636 35258 30636 35258 4 _0357_
rlabel metal2 s 30314 33728 30314 33728 4 _0358_
rlabel metal2 s 30130 31994 30130 31994 4 _0359_
rlabel metal2 s 32246 36856 32246 36856 4 _0360_
rlabel metal1 s 32706 36550 32706 36550 4 _0361_
rlabel metal1 s 32430 34578 32430 34578 4 _0362_
rlabel metal2 s 33350 36346 33350 36346 4 _0363_
rlabel metal1 s 33534 36176 33534 36176 4 _0364_
rlabel metal2 s 33626 35462 33626 35462 4 _0365_
rlabel metal1 s 33902 33490 33902 33490 4 _0366_
rlabel metal1 s 33764 33626 33764 33626 4 _0367_
rlabel metal1 s 34960 34034 34960 34034 4 _0368_
rlabel metal2 s 34638 33201 34638 33201 4 _0369_
rlabel metal1 s 34116 33558 34116 33558 4 _0370_
rlabel metal1 s 34592 31382 34592 31382 4 _0371_
rlabel metal1 s 34546 33082 34546 33082 4 _0372_
rlabel metal1 s 34822 32266 34822 32266 4 _0373_
rlabel metal1 s 31970 31348 31970 31348 4 _0374_
rlabel metal1 s 26082 36346 26082 36346 4 _0375_
rlabel metal2 s 29578 5372 29578 5372 4 _0376_
rlabel metal2 s 3542 15300 3542 15300 4 _0377_
rlabel metal1 s 4002 14416 4002 14416 4 _0378_
rlabel metal2 s 3826 17238 3826 17238 4 _0379_
rlabel metal2 s 3450 15878 3450 15878 4 _0380_
rlabel metal2 s 4554 17306 4554 17306 4 _0381_
rlabel metal1 s 4324 17646 4324 17646 4 _0382_
rlabel metal1 s 4094 19346 4094 19346 4 _0383_
rlabel metal1 s 4508 19346 4508 19346 4 _0384_
rlabel metal2 s 2622 19006 2622 19006 4 _0385_
rlabel metal1 s 2158 19482 2158 19482 4 _0386_
rlabel metal1 s 5566 14926 5566 14926 4 _0387_
rlabel metal1 s 5428 14994 5428 14994 4 _0388_
rlabel metal2 s 7682 15572 7682 15572 4 _0389_
rlabel metal2 s 7774 15538 7774 15538 4 _0390_
rlabel metal1 s 9614 14450 9614 14450 4 _0391_
rlabel metal2 s 9246 14620 9246 14620 4 _0392_
rlabel metal1 s 10764 17646 10764 17646 4 _0393_
rlabel metal2 s 11086 15538 11086 15538 4 _0394_
rlabel metal1 s 9936 17170 9936 17170 4 _0395_
rlabel metal1 s 10258 17680 10258 17680 4 _0396_
rlabel metal1 s 7728 17102 7728 17102 4 _0397_
rlabel metal1 s 9062 16762 9062 16762 4 _0398_
rlabel metal1 s 8556 23698 8556 23698 4 _0399_
rlabel metal2 s 9982 30906 9982 30906 4 _0400_
rlabel metal2 s 10534 29716 10534 29716 4 _0401_
rlabel metal1 s 4416 16626 4416 16626 4 _0402_
rlabel metal1 s 35328 8602 35328 8602 4 _0403_
rlabel metal2 s 30774 32572 30774 32572 4 _0404_
rlabel metal2 s 10074 25466 10074 25466 4 _0405_
rlabel metal2 s 10166 24650 10166 24650 4 _0406_
rlabel metal2 s 10258 27166 10258 27166 4 _0407_
rlabel metal1 s 6210 26350 6210 26350 4 _0408_
rlabel metal1 s 6256 25466 6256 25466 4 _0409_
rlabel metal1 s 6394 26418 6394 26418 4 _0410_
rlabel metal1 s 5934 21862 5934 21862 4 _0411_
rlabel metal1 s 10166 25194 10166 25194 4 _0412_
rlabel metal1 s 8188 25330 8188 25330 4 _0413_
rlabel metal1 s 6716 25398 6716 25398 4 _0414_
rlabel metal1 s 33442 4590 33442 4590 4 _0415_
rlabel metal2 s 35098 5440 35098 5440 4 _0416_
rlabel metal1 s 34316 6698 34316 6698 4 _0417_
rlabel metal1 s 32706 6290 32706 6290 4 _0418_
rlabel metal1 s 31280 6834 31280 6834 4 _0419_
rlabel metal2 s 34914 5151 34914 5151 4 _0420_
rlabel metal1 s 29854 34578 29854 34578 4 _0421_
rlabel metal1 s 30498 34544 30498 34544 4 _0422_
rlabel metal1 s 30268 32198 30268 32198 4 _0423_
rlabel metal1 s 29762 32368 29762 32368 4 _0424_
rlabel metal2 s 29578 36448 29578 36448 4 _0425_
rlabel metal2 s 31878 33966 31878 33966 4 _0426_
rlabel metal2 s 2254 25772 2254 25772 4 _0427_
rlabel metal1 s 4094 28492 4094 28492 4 _0428_
rlabel metal1 s 4508 16694 4508 16694 4 _0429_
rlabel metal2 s 4094 16388 4094 16388 4 _0430_
rlabel metal1 s 4784 16558 4784 16558 4 _0431_
rlabel metal1 s 2484 27982 2484 27982 4 _0432_
rlabel metal1 s 4416 27642 4416 27642 4 _0433_
rlabel metal1 s 4102 29206 4102 29206 4 _0434_
rlabel metal2 s 7498 21114 7498 21114 4 _0435_
rlabel metal1 s 4188 21998 4188 21998 4 _0436_
rlabel metal1 s 2392 28390 2392 28390 4 _0437_
rlabel metal1 s 4600 28662 4600 28662 4 _0438_
rlabel metal1 s 4416 29614 4416 29614 4 _0439_
rlabel metal1 s 4232 29478 4232 29478 4 _0440_
rlabel metal1 s 5474 27302 5474 27302 4 _0441_
rlabel metal2 s 5842 29716 5842 29716 4 _0442_
rlabel metal1 s 6302 30158 6302 30158 4 _0443_
rlabel metal1 s 5796 28186 5796 28186 4 _0444_
rlabel metal2 s 6026 27336 6026 27336 4 _0445_
rlabel metal1 s 5750 27438 5750 27438 4 _0446_
rlabel metal3 s 7130 26741 7130 26741 4 _0447_
rlabel metal1 s 7314 22066 7314 22066 4 _0448_
rlabel metal1 s 6131 27098 6131 27098 4 _0449_
rlabel metal1 s 7452 24174 7452 24174 4 _0450_
rlabel metal1 s 5198 24820 5198 24820 4 _0451_
rlabel metal2 s 4830 25874 4830 25874 4 _0452_
rlabel metal1 s 5750 26826 5750 26826 4 _0453_
rlabel metal1 s 5198 23528 5198 23528 4 _0454_
rlabel metal2 s 6578 24140 6578 24140 4 _0455_
rlabel metal1 s 6256 21862 6256 21862 4 _0456_
rlabel metal1 s 4968 23290 4968 23290 4 _0457_
rlabel metal2 s 2714 22814 2714 22814 4 _0458_
rlabel metal1 s 2208 22610 2208 22610 4 _0459_
rlabel metal1 s 3910 22202 3910 22202 4 _0460_
rlabel metal2 s 4370 21879 4370 21879 4 _0461_
rlabel metal2 s 4094 21165 4094 21165 4 _0462_
rlabel metal2 s 6302 22440 6302 22440 4 _0463_
rlabel metal1 s 7774 21998 7774 21998 4 _0464_
rlabel metal1 s 7820 20910 7820 20910 4 _0465_
rlabel metal2 s 6946 21250 6946 21250 4 _0466_
rlabel metal1 s 6532 21522 6532 21522 4 _0467_
rlabel metal2 s 8142 20230 8142 20230 4 _0468_
rlabel metal1 s 8510 20570 8510 20570 4 _0469_
rlabel metal1 s 9108 20910 9108 20910 4 _0470_
rlabel metal1 s 9108 20434 9108 20434 4 _0471_
rlabel metal2 s 9798 20332 9798 20332 4 _0472_
rlabel metal1 s 9292 21454 9292 21454 4 _0473_
rlabel metal1 s 10488 21658 10488 21658 4 _0474_
rlabel metal2 s 9982 21284 9982 21284 4 _0475_
rlabel metal1 s 10304 23290 10304 23290 4 _0476_
rlabel metal2 s 10534 23222 10534 23222 4 _0477_
rlabel metal1 s 10258 22576 10258 22576 4 _0478_
rlabel metal1 s 9200 23290 9200 23290 4 _0479_
rlabel metal1 s 9246 22542 9246 22542 4 _0480_
rlabel metal2 s 8694 23120 8694 23120 4 _0481_
rlabel metal1 s 9752 25806 9752 25806 4 _0482_
rlabel metal2 s 8970 26554 8970 26554 4 _0483_
rlabel metal1 s 9292 26282 9292 26282 4 _0484_
rlabel metal1 s 10580 25466 10580 25466 4 _0485_
rlabel metal2 s 10166 26180 10166 26180 4 _0486_
rlabel metal1 s 10396 26554 10396 26554 4 _0487_
rlabel metal1 s 11178 26996 11178 26996 4 _0488_
rlabel metal1 s 10350 26860 10350 26860 4 _0489_
rlabel metal1 s 10028 27438 10028 27438 4 _0490_
rlabel metal1 s 9522 27098 9522 27098 4 _0491_
rlabel metal1 s 9200 27030 9200 27030 4 _0492_
rlabel metal2 s 8326 29172 8326 29172 4 _0493_
rlabel metal2 s 8142 30022 8142 30022 4 _0494_
rlabel metal2 s 7866 30022 7866 30022 4 _0495_
rlabel metal2 s 8602 30566 8602 30566 4 _0496_
rlabel metal1 s 9614 30634 9614 30634 4 _0497_
rlabel metal1 s 10626 30124 10626 30124 4 _0498_
rlabel metal2 s 10810 29716 10810 29716 4 _0499_
rlabel metal1 s 30268 6834 30268 6834 4 _0500_
rlabel metal1 s 33994 3570 33994 3570 4 _0501_
rlabel metal1 s 30498 5134 30498 5134 4 _0502_
rlabel metal1 s 30958 5270 30958 5270 4 _0503_
rlabel metal1 s 31418 5168 31418 5168 4 _0504_
rlabel metal2 s 31326 4318 31326 4318 4 _0505_
rlabel metal1 s 32154 3706 32154 3706 4 _0506_
rlabel metal1 s 33350 3536 33350 3536 4 _0507_
rlabel metal1 s 32154 3536 32154 3536 4 _0508_
rlabel metal2 s 35550 4522 35550 4522 4 _0509_
rlabel metal1 s 35420 4794 35420 4794 4 _0510_
rlabel metal2 s 33626 6120 33626 6120 4 _0511_
rlabel metal1 s 34086 6358 34086 6358 4 _0512_
rlabel metal1 s 33120 8330 33120 8330 4 _0513_
rlabel metal2 s 29670 9588 29670 9588 4 _0514_
rlabel metal2 s 31418 8670 31418 8670 4 _0515_
rlabel metal1 s 31648 10642 31648 10642 4 _0516_
rlabel metal1 s 30314 10064 30314 10064 4 _0517_
rlabel metal1 s 30314 10574 30314 10574 4 _0518_
rlabel metal2 s 31786 10948 31786 10948 4 _0519_
rlabel metal1 s 31234 11696 31234 11696 4 _0520_
rlabel metal1 s 33994 9520 33994 9520 4 _0521_
rlabel metal1 s 34454 9384 34454 9384 4 _0522_
rlabel metal1 s 32384 9146 32384 9146 4 _0523_
rlabel metal2 s 34730 10642 34730 10642 4 _0524_
rlabel metal1 s 34500 9486 34500 9486 4 _0525_
rlabel metal2 s 35466 10710 35466 10710 4 _0526_
rlabel metal1 s 34362 11084 34362 11084 4 _0527_
rlabel metal3 s 912 29308 912 29308 4 clk
rlabel metal1 s 23000 10030 23000 10030 4 clknet_0_A_in_serial_clk
rlabel metal2 s 25806 26081 25806 26081 4 clknet_0_B_in_serial_clk
rlabel metal1 s 7728 18326 7728 18326 4 clknet_0_clk
rlabel metal2 s 1426 21488 1426 21488 4 clknet_2_0__leaf_clk
rlabel metal2 s 6394 19856 6394 19856 4 clknet_2_1__leaf_clk
rlabel metal1 s 1426 26826 1426 26826 4 clknet_2_2__leaf_clk
rlabel metal2 s 10350 24752 10350 24752 4 clknet_2_3__leaf_clk
rlabel metal2 s 19090 6800 19090 6800 4 clknet_4_0_0_A_in_serial_clk
rlabel metal1 s 15870 21998 15870 21998 4 clknet_4_0_0_B_in_serial_clk
rlabel metal1 s 33534 6222 33534 6222 4 clknet_4_10_0_A_in_serial_clk
rlabel metal1 s 29486 23086 29486 23086 4 clknet_4_10_0_B_in_serial_clk
rlabel metal1 s 30958 12274 30958 12274 4 clknet_4_11_0_A_in_serial_clk
rlabel metal1 s 28888 26894 28888 26894 4 clknet_4_11_0_B_in_serial_clk
rlabel metal2 s 26266 14212 26266 14212 4 clknet_4_12_0_A_in_serial_clk
rlabel metal2 s 24426 30464 24426 30464 4 clknet_4_12_0_B_in_serial_clk
rlabel metal1 s 26404 17714 26404 17714 4 clknet_4_13_0_A_in_serial_clk
rlabel metal2 s 24426 33728 24426 33728 4 clknet_4_13_0_B_in_serial_clk
rlabel metal2 s 34454 14144 34454 14144 4 clknet_4_14_0_A_in_serial_clk
rlabel metal1 s 31142 31314 31142 31314 4 clknet_4_14_0_B_in_serial_clk
rlabel metal1 s 34132 20434 34132 20434 4 clknet_4_15_0_A_in_serial_clk
rlabel metal2 s 29854 36448 29854 36448 4 clknet_4_15_0_B_in_serial_clk
rlabel metal2 s 13754 11152 13754 11152 4 clknet_4_1_0_A_in_serial_clk
rlabel metal2 s 16422 26690 16422 26690 4 clknet_4_1_0_B_in_serial_clk
rlabel metal1 s 23598 5270 23598 5270 4 clknet_4_2_0_A_in_serial_clk
rlabel metal1 s 20700 22066 20700 22066 4 clknet_4_2_0_B_in_serial_clk
rlabel metal2 s 23598 9826 23598 9826 4 clknet_4_3_0_A_in_serial_clk
rlabel metal1 s 19182 28594 19182 28594 4 clknet_4_3_0_B_in_serial_clk
rlabel metal1 s 17802 16626 17802 16626 4 clknet_4_4_0_A_in_serial_clk
rlabel metal1 s 11730 31790 11730 31790 4 clknet_4_4_0_B_in_serial_clk
rlabel metal2 s 16882 17408 16882 17408 4 clknet_4_5_0_A_in_serial_clk
rlabel metal1 s 11500 36006 11500 36006 4 clknet_4_5_0_B_in_serial_clk
rlabel metal2 s 21850 15266 21850 15266 4 clknet_4_6_0_A_in_serial_clk
rlabel metal1 s 19826 32266 19826 32266 4 clknet_4_6_0_B_in_serial_clk
rlabel metal1 s 21850 20298 21850 20298 4 clknet_4_7_0_A_in_serial_clk
rlabel metal2 s 20562 36380 20562 36380 4 clknet_4_7_0_B_in_serial_clk
rlabel metal1 s 25576 5678 25576 5678 4 clknet_4_8_0_A_in_serial_clk
rlabel metal1 s 24058 24242 24058 24242 4 clknet_4_8_0_B_in_serial_clk
rlabel metal2 s 27002 9248 27002 9248 4 clknet_4_9_0_A_in_serial_clk
rlabel metal1 s 24426 25976 24426 25976 4 clknet_4_9_0_B_in_serial_clk
rlabel metal1 s 32338 6222 32338 6222 4 deser_A.bit_idx\[0\]
rlabel metal1 s 33442 4182 33442 4182 4 deser_A.bit_idx\[1\]
rlabel metal1 s 30544 4046 30544 4046 4 deser_A.bit_idx\[2\]
rlabel metal1 s 32108 4590 32108 4590 4 deser_A.bit_idx\[3\]
rlabel metal1 s 35098 4692 35098 4692 4 deser_A.bit_idx\[4\]
rlabel metal2 s 33442 5440 33442 5440 4 deser_A.bit_idx\[5\]
rlabel metal1 s 33166 5780 33166 5780 4 deser_A.bit_idx\[6\]
rlabel metal1 s 34546 6834 34546 6834 4 deser_A.bit_idx\[7\]
rlabel metal1 s 31786 8500 31786 8500 4 deser_A.kept_bit_idx\[0\]
rlabel metal1 s 30866 8874 30866 8874 4 deser_A.kept_bit_idx\[1\]
rlabel metal1 s 30268 9962 30268 9962 4 deser_A.kept_bit_idx\[2\]
rlabel metal2 s 31878 10132 31878 10132 4 deser_A.kept_bit_idx\[3\]
rlabel metal1 s 32246 10031 32246 10031 4 deser_A.kept_bit_idx\[4\]
rlabel metal1 s 32614 9010 32614 9010 4 deser_A.kept_bit_idx\[5\]
rlabel metal1 s 35190 9554 35190 9554 4 deser_A.kept_bit_idx\[6\]
rlabel metal2 s 34454 10268 34454 10268 4 deser_A.kept_bit_idx\[7\]
rlabel metal1 s 35512 8466 35512 8466 4 deser_A.kept_receiving
rlabel metal2 s 29946 5678 29946 5678 4 deser_A.kept_shift_reg\[0\]
rlabel metal2 s 15870 15946 15870 15946 4 deser_A.kept_shift_reg\[100\]
rlabel metal1 s 16238 16966 16238 16966 4 deser_A.kept_shift_reg\[101\]
rlabel metal1 s 16468 18394 16468 18394 4 deser_A.kept_shift_reg\[102\]
rlabel metal1 s 15824 18802 15824 18802 4 deser_A.kept_shift_reg\[103\]
rlabel metal2 s 15594 19482 15594 19482 4 deser_A.kept_shift_reg\[104\]
rlabel metal1 s 17434 19414 17434 19414 4 deser_A.kept_shift_reg\[105\]
rlabel metal1 s 18170 20366 18170 20366 4 deser_A.kept_shift_reg\[106\]
rlabel metal2 s 18446 20230 18446 20230 4 deser_A.kept_shift_reg\[107\]
rlabel metal1 s 18538 18938 18538 18938 4 deser_A.kept_shift_reg\[108\]
rlabel metal2 s 19090 18088 19090 18088 4 deser_A.kept_shift_reg\[109\]
rlabel metal1 s 29072 13226 29072 13226 4 deser_A.kept_shift_reg\[10\]
rlabel metal1 s 18906 17102 18906 17102 4 deser_A.kept_shift_reg\[110\]
rlabel metal1 s 18262 15538 18262 15538 4 deser_A.kept_shift_reg\[111\]
rlabel metal1 s 18216 14790 18216 14790 4 deser_A.kept_shift_reg\[112\]
rlabel metal2 s 18078 14144 18078 14144 4 deser_A.kept_shift_reg\[113\]
rlabel metal1 s 19090 13872 19090 13872 4 deser_A.kept_shift_reg\[114\]
rlabel metal1 s 18170 11764 18170 11764 4 deser_A.kept_shift_reg\[115\]
rlabel metal1 s 17204 10642 17204 10642 4 deser_A.kept_shift_reg\[116\]
rlabel metal2 s 17894 10608 17894 10608 4 deser_A.kept_shift_reg\[117\]
rlabel metal1 s 18676 8942 18676 8942 4 deser_A.kept_shift_reg\[118\]
rlabel metal1 s 19136 9010 19136 9010 4 deser_A.kept_shift_reg\[119\]
rlabel metal1 s 29624 12410 29624 12410 4 deser_A.kept_shift_reg\[11\]
rlabel metal2 s 20562 7548 20562 7548 4 deser_A.kept_shift_reg\[120\]
rlabel metal1 s 22379 6766 22379 6766 4 deser_A.kept_shift_reg\[121\]
rlabel metal1 s 21436 5882 21436 5882 4 deser_A.kept_shift_reg\[122\]
rlabel metal1 s 21666 4590 21666 4590 4 deser_A.kept_shift_reg\[123\]
rlabel metal2 s 22126 5253 22126 5253 4 deser_A.kept_shift_reg\[124\]
rlabel metal2 s 22310 5984 22310 5984 4 deser_A.kept_shift_reg\[125\]
rlabel metal1 s 24104 4998 24104 4998 4 deser_A.kept_shift_reg\[126\]
rlabel metal2 s 25162 5916 25162 5916 4 deser_A.kept_shift_reg\[127\]
rlabel metal1 s 32315 12750 32315 12750 4 deser_A.kept_shift_reg\[12\]
rlabel metal2 s 32430 13668 32430 13668 4 deser_A.kept_shift_reg\[13\]
rlabel metal1 s 35466 12342 35466 12342 4 deser_A.kept_shift_reg\[14\]
rlabel metal1 s 35282 12614 35282 12614 4 deser_A.kept_shift_reg\[15\]
rlabel metal2 s 35466 14620 35466 14620 4 deser_A.kept_shift_reg\[16\]
rlabel metal2 s 34362 14348 34362 14348 4 deser_A.kept_shift_reg\[17\]
rlabel metal2 s 33534 15062 33534 15062 4 deser_A.kept_shift_reg\[18\]
rlabel metal2 s 32154 15028 32154 15028 4 deser_A.kept_shift_reg\[19\]
rlabel metal2 s 28566 6018 28566 6018 4 deser_A.kept_shift_reg\[1\]
rlabel metal1 s 32016 15470 32016 15470 4 deser_A.kept_shift_reg\[20\]
rlabel metal1 s 29072 15402 29072 15402 4 deser_A.kept_shift_reg\[21\]
rlabel metal1 s 29440 16762 29440 16762 4 deser_A.kept_shift_reg\[22\]
rlabel metal2 s 28842 16184 28842 16184 4 deser_A.kept_shift_reg\[23\]
rlabel metal1 s 28060 14586 28060 14586 4 deser_A.kept_shift_reg\[24\]
rlabel metal1 s 26358 13838 26358 13838 4 deser_A.kept_shift_reg\[25\]
rlabel metal2 s 26174 13804 26174 13804 4 deser_A.kept_shift_reg\[26\]
rlabel metal2 s 24978 13124 24978 13124 4 deser_A.kept_shift_reg\[27\]
rlabel metal1 s 24932 11866 24932 11866 4 deser_A.kept_shift_reg\[28\]
rlabel metal2 s 25070 11594 25070 11594 4 deser_A.kept_shift_reg\[29\]
rlabel metal2 s 27462 6018 27462 6018 4 deser_A.kept_shift_reg\[2\]
rlabel metal2 s 25162 10438 25162 10438 4 deser_A.kept_shift_reg\[30\]
rlabel metal2 s 26174 10166 26174 10166 4 deser_A.kept_shift_reg\[31\]
rlabel metal1 s 25852 6834 25852 6834 4 deser_A.kept_shift_reg\[32\]
rlabel metal1 s 25852 7514 25852 7514 4 deser_A.kept_shift_reg\[33\]
rlabel metal1 s 23644 8398 23644 8398 4 deser_A.kept_shift_reg\[34\]
rlabel metal2 s 23782 8126 23782 8126 4 deser_A.kept_shift_reg\[35\]
rlabel metal2 s 23690 9894 23690 9894 4 deser_A.kept_shift_reg\[36\]
rlabel metal1 s 22402 11118 22402 11118 4 deser_A.kept_shift_reg\[37\]
rlabel metal2 s 22586 10676 22586 10676 4 deser_A.kept_shift_reg\[38\]
rlabel metal2 s 22954 11628 22954 11628 4 deser_A.kept_shift_reg\[39\]
rlabel metal1 s 27922 5746 27922 5746 4 deser_A.kept_shift_reg\[3\]
rlabel metal1 s 21942 13906 21942 13906 4 deser_A.kept_shift_reg\[40\]
rlabel metal2 s 21482 15198 21482 15198 4 deser_A.kept_shift_reg\[41\]
rlabel metal1 s 20746 17238 20746 17238 4 deser_A.kept_shift_reg\[42\]
rlabel metal1 s 21114 17170 21114 17170 4 deser_A.kept_shift_reg\[43\]
rlabel metal2 s 22402 18326 22402 18326 4 deser_A.kept_shift_reg\[44\]
rlabel metal1 s 21620 18598 21620 18598 4 deser_A.kept_shift_reg\[45\]
rlabel metal1 s 20976 19346 20976 19346 4 deser_A.kept_shift_reg\[46\]
rlabel metal1 s 21206 20366 21206 20366 4 deser_A.kept_shift_reg\[47\]
rlabel metal2 s 22862 20740 22862 20740 4 deser_A.kept_shift_reg\[48\]
rlabel metal2 s 23690 20774 23690 20774 4 deser_A.kept_shift_reg\[49\]
rlabel metal1 s 27692 7514 27692 7514 4 deser_A.kept_shift_reg\[4\]
rlabel metal1 s 24472 20026 24472 20026 4 deser_A.kept_shift_reg\[50\]
rlabel metal1 s 23920 18190 23920 18190 4 deser_A.kept_shift_reg\[51\]
rlabel metal2 s 24150 18462 24150 18462 4 deser_A.kept_shift_reg\[52\]
rlabel metal1 s 25530 17850 25530 17850 4 deser_A.kept_shift_reg\[53\]
rlabel metal2 s 26174 18989 26174 18989 4 deser_A.kept_shift_reg\[54\]
rlabel metal2 s 26542 20230 26542 20230 4 deser_A.kept_shift_reg\[55\]
rlabel metal1 s 27738 20230 27738 20230 4 deser_A.kept_shift_reg\[56\]
rlabel metal1 s 28750 20774 28750 20774 4 deser_A.kept_shift_reg\[57\]
rlabel metal2 s 29578 21318 29578 21318 4 deser_A.kept_shift_reg\[58\]
rlabel metal1 s 30682 21454 30682 21454 4 deser_A.kept_shift_reg\[59\]
rlabel metal2 s 28750 9350 28750 9350 4 deser_A.kept_shift_reg\[5\]
rlabel metal2 s 31602 21284 31602 21284 4 deser_A.kept_shift_reg\[60\]
rlabel metal2 s 32798 21012 32798 21012 4 deser_A.kept_shift_reg\[61\]
rlabel metal2 s 34454 20604 34454 20604 4 deser_A.kept_shift_reg\[62\]
rlabel metal1 s 35006 19890 35006 19890 4 deser_A.kept_shift_reg\[63\]
rlabel metal1 s 35190 18734 35190 18734 4 deser_A.kept_shift_reg\[64\]
rlabel metal1 s 34362 18598 34362 18598 4 deser_A.kept_shift_reg\[65\]
rlabel metal1 s 33948 17510 33948 17510 4 deser_A.kept_shift_reg\[66\]
rlabel metal2 s 33534 16490 33534 16490 4 deser_A.kept_shift_reg\[67\]
rlabel metal2 s 31970 16949 31970 16949 4 deser_A.kept_shift_reg\[68\]
rlabel metal2 s 31970 18088 31970 18088 4 deser_A.kept_shift_reg\[69\]
rlabel metal1 s 28704 9690 28704 9690 4 deser_A.kept_shift_reg\[6\]
rlabel metal1 s 31510 19278 31510 19278 4 deser_A.kept_shift_reg\[70\]
rlabel metal2 s 30314 19380 30314 19380 4 deser_A.kept_shift_reg\[71\]
rlabel metal1 s 29486 18394 29486 18394 4 deser_A.kept_shift_reg\[72\]
rlabel metal1 s 26864 17306 26864 17306 4 deser_A.kept_shift_reg\[73\]
rlabel metal1 s 26312 16422 26312 16422 4 deser_A.kept_shift_reg\[74\]
rlabel metal1 s 25852 16014 25852 16014 4 deser_A.kept_shift_reg\[75\]
rlabel metal1 s 24610 16422 24610 16422 4 deser_A.kept_shift_reg\[76\]
rlabel metal1 s 23460 15674 23460 15674 4 deser_A.kept_shift_reg\[77\]
rlabel metal2 s 23966 14722 23966 14722 4 deser_A.kept_shift_reg\[78\]
rlabel metal1 s 23092 13498 23092 13498 4 deser_A.kept_shift_reg\[79\]
rlabel metal1 s 26634 12070 26634 12070 4 deser_A.kept_shift_reg\[7\]
rlabel metal2 s 20700 12308 20700 12308 4 deser_A.kept_shift_reg\[80\]
rlabel metal1 s 20240 11526 20240 11526 4 deser_A.kept_shift_reg\[81\]
rlabel metal1 s 20102 10030 20102 10030 4 deser_A.kept_shift_reg\[82\]
rlabel metal2 s 18446 10370 18446 10370 4 deser_A.kept_shift_reg\[83\]
rlabel metal1 s 18395 8398 18395 8398 4 deser_A.kept_shift_reg\[84\]
rlabel metal1 s 18860 7174 18860 7174 4 deser_A.kept_shift_reg\[85\]
rlabel metal1 s 18262 6290 18262 6290 4 deser_A.kept_shift_reg\[86\]
rlabel metal2 s 18354 5372 18354 5372 4 deser_A.kept_shift_reg\[87\]
rlabel metal1 s 16928 4794 16928 4794 4 deser_A.kept_shift_reg\[88\]
rlabel metal1 s 16146 5712 16146 5712 4 deser_A.kept_shift_reg\[89\]
rlabel metal1 s 26726 11220 26726 11220 4 deser_A.kept_shift_reg\[8\]
rlabel metal1 s 15502 6086 15502 6086 4 deser_A.kept_shift_reg\[90\]
rlabel metal1 s 15916 7378 15916 7378 4 deser_A.kept_shift_reg\[91\]
rlabel metal1 s 15548 8602 15548 8602 4 deser_A.kept_shift_reg\[92\]
rlabel metal1 s 15456 9690 15456 9690 4 deser_A.kept_shift_reg\[93\]
rlabel metal1 s 15732 10778 15732 10778 4 deser_A.kept_shift_reg\[94\]
rlabel metal1 s 15916 11866 15916 11866 4 deser_A.kept_shift_reg\[95\]
rlabel metal1 s 16008 12614 16008 12614 4 deser_A.kept_shift_reg\[96\]
rlabel metal1 s 15962 13362 15962 13362 4 deser_A.kept_shift_reg\[97\]
rlabel metal2 s 15778 14756 15778 14756 4 deser_A.kept_shift_reg\[98\]
rlabel metal2 s 15686 15674 15686 15674 4 deser_A.kept_shift_reg\[99\]
rlabel metal1 s 27508 11866 27508 11866 4 deser_A.kept_shift_reg\[9\]
rlabel metal2 s 34086 8398 34086 8398 4 deser_A.receiving
rlabel metal1 s 26542 35598 26542 35598 4 deser_B.bit_idx\[0\]
rlabel metal1 s 28014 37230 28014 37230 4 deser_B.bit_idx\[1\]
rlabel metal1 s 28888 36346 28888 36346 4 deser_B.bit_idx\[2\]
rlabel metal2 s 28198 34714 28198 34714 4 deser_B.bit_idx\[3\]
rlabel metal1 s 29072 33422 29072 33422 4 deser_B.bit_idx\[4\]
rlabel metal2 s 31878 35037 31878 35037 4 deser_B.bit_idx\[5\]
rlabel metal2 s 31602 34000 31602 34000 4 deser_B.bit_idx\[6\]
rlabel metal1 s 28934 31450 28934 31450 4 deser_B.bit_idx\[7\]
rlabel metal1 s 32062 36074 32062 36074 4 deser_B.kept_bit_idx\[0\]
rlabel metal1 s 33028 36822 33028 36822 4 deser_B.kept_bit_idx\[1\]
rlabel metal2 s 32982 37400 32982 37400 4 deser_B.kept_bit_idx\[2\]
rlabel metal2 s 35650 35258 35650 35258 4 deser_B.kept_bit_idx\[3\]
rlabel metal2 s 33258 34510 33258 34510 4 deser_B.kept_bit_idx\[4\]
rlabel metal1 s 33350 34170 33350 34170 4 deser_B.kept_bit_idx\[5\]
rlabel metal1 s 35144 32198 35144 32198 4 deser_B.kept_bit_idx\[6\]
rlabel metal1 s 34500 31926 34500 31926 4 deser_B.kept_bit_idx\[7\]
rlabel metal1 s 31234 30906 31234 30906 4 deser_B.kept_receiving
rlabel metal2 s 26636 36754 26636 36754 4 deser_B.kept_shift_reg\[0\]
rlabel metal1 s 14904 31858 14904 31858 4 deser_B.kept_shift_reg\[100\]
rlabel metal1 s 13340 31994 13340 31994 4 deser_B.kept_shift_reg\[101\]
rlabel metal1 s 13202 33626 13202 33626 4 deser_B.kept_shift_reg\[102\]
rlabel metal1 s 12742 34646 12742 34646 4 deser_B.kept_shift_reg\[103\]
rlabel metal2 s 11914 35462 11914 35462 4 deser_B.kept_shift_reg\[104\]
rlabel metal1 s 12834 36346 12834 36346 4 deser_B.kept_shift_reg\[105\]
rlabel metal2 s 12558 37366 12558 37366 4 deser_B.kept_shift_reg\[106\]
rlabel metal1 s 13018 36550 13018 36550 4 deser_B.kept_shift_reg\[107\]
rlabel metal1 s 15410 37434 15410 37434 4 deser_B.kept_shift_reg\[108\]
rlabel metal1 s 16468 36890 16468 36890 4 deser_B.kept_shift_reg\[109\]
rlabel metal2 s 30130 29070 30130 29070 4 deser_B.kept_shift_reg\[10\]
rlabel metal2 s 17158 36283 17158 36283 4 deser_B.kept_shift_reg\[110\]
rlabel metal1 s 16974 34578 16974 34578 4 deser_B.kept_shift_reg\[111\]
rlabel metal1 s 17848 33898 17848 33898 4 deser_B.kept_shift_reg\[112\]
rlabel metal1 s 17756 33830 17756 33830 4 deser_B.kept_shift_reg\[113\]
rlabel metal1 s 17526 33490 17526 33490 4 deser_B.kept_shift_reg\[114\]
rlabel metal2 s 18078 32980 18078 32980 4 deser_B.kept_shift_reg\[115\]
rlabel metal1 s 20378 33490 20378 33490 4 deser_B.kept_shift_reg\[116\]
rlabel metal2 s 20562 34816 20562 34816 4 deser_B.kept_shift_reg\[117\]
rlabel metal2 s 19090 35462 19090 35462 4 deser_B.kept_shift_reg\[118\]
rlabel metal1 s 18906 36346 18906 36346 4 deser_B.kept_shift_reg\[119\]
rlabel metal2 s 31970 29580 31970 29580 4 deser_B.kept_shift_reg\[11\]
rlabel metal1 s 18814 37434 18814 37434 4 deser_B.kept_shift_reg\[120\]
rlabel metal1 s 18768 36890 18768 36890 4 deser_B.kept_shift_reg\[121\]
rlabel metal2 s 20102 36822 20102 36822 4 deser_B.kept_shift_reg\[122\]
rlabel metal1 s 21390 36346 21390 36346 4 deser_B.kept_shift_reg\[123\]
rlabel metal1 s 21620 36550 21620 36550 4 deser_B.kept_shift_reg\[124\]
rlabel metal2 s 24150 36244 24150 36244 4 deser_B.kept_shift_reg\[125\]
rlabel metal2 s 23874 37604 23874 37604 4 deser_B.kept_shift_reg\[126\]
rlabel metal1 s 24058 37434 24058 37434 4 deser_B.kept_shift_reg\[127\]
rlabel metal2 s 32430 30566 32430 30566 4 deser_B.kept_shift_reg\[12\]
rlabel metal1 s 34316 29274 34316 29274 4 deser_B.kept_shift_reg\[13\]
rlabel metal2 s 33442 29036 33442 29036 4 deser_B.kept_shift_reg\[14\]
rlabel metal2 s 33994 28084 33994 28084 4 deser_B.kept_shift_reg\[15\]
rlabel metal1 s 33810 26010 33810 26010 4 deser_B.kept_shift_reg\[16\]
rlabel metal1 s 33764 25330 33764 25330 4 deser_B.kept_shift_reg\[17\]
rlabel metal2 s 34546 24786 34546 24786 4 deser_B.kept_shift_reg\[18\]
rlabel metal2 s 34454 23460 34454 23460 4 deser_B.kept_shift_reg\[19\]
rlabel metal2 s 25990 35700 25990 35700 4 deser_B.kept_shift_reg\[1\]
rlabel metal2 s 33902 23222 33902 23222 4 deser_B.kept_shift_reg\[20\]
rlabel metal2 s 31786 24922 31786 24922 4 deser_B.kept_shift_reg\[21\]
rlabel metal1 s 31280 24378 31280 24378 4 deser_B.kept_shift_reg\[22\]
rlabel metal1 s 29716 24582 29716 24582 4 deser_B.kept_shift_reg\[23\]
rlabel metal1 s 28658 24922 28658 24922 4 deser_B.kept_shift_reg\[24\]
rlabel metal1 s 28152 24378 28152 24378 4 deser_B.kept_shift_reg\[25\]
rlabel metal2 s 27462 24446 27462 24446 4 deser_B.kept_shift_reg\[26\]
rlabel metal1 s 26036 24378 26036 24378 4 deser_B.kept_shift_reg\[27\]
rlabel metal1 s 24334 24582 24334 24582 4 deser_B.kept_shift_reg\[28\]
rlabel metal1 s 23506 24718 23506 24718 4 deser_B.kept_shift_reg\[29\]
rlabel metal1 s 25484 34714 25484 34714 4 deser_B.kept_shift_reg\[2\]
rlabel metal1 s 22954 25296 22954 25296 4 deser_B.kept_shift_reg\[30\]
rlabel metal2 s 22494 27200 22494 27200 4 deser_B.kept_shift_reg\[31\]
rlabel metal2 s 22218 26860 22218 26860 4 deser_B.kept_shift_reg\[32\]
rlabel metal2 s 22310 26588 22310 26588 4 deser_B.kept_shift_reg\[33\]
rlabel metal1 s 23598 26758 23598 26758 4 deser_B.kept_shift_reg\[34\]
rlabel metal1 s 23782 27540 23782 27540 4 deser_B.kept_shift_reg\[35\]
rlabel metal1 s 25346 25840 25346 25840 4 deser_B.kept_shift_reg\[36\]
rlabel metal1 s 25829 25874 25829 25874 4 deser_B.kept_shift_reg\[37\]
rlabel metal2 s 27738 26928 27738 26928 4 deser_B.kept_shift_reg\[38\]
rlabel metal1 s 29624 26894 29624 26894 4 deser_B.kept_shift_reg\[39\]
rlabel metal1 s 26266 33626 26266 33626 4 deser_B.kept_shift_reg\[3\]
rlabel metal1 s 30728 27982 30728 27982 4 deser_B.kept_shift_reg\[40\]
rlabel metal1 s 30452 26010 30452 26010 4 deser_B.kept_shift_reg\[41\]
rlabel metal1 s 30774 23630 30774 23630 4 deser_B.kept_shift_reg\[42\]
rlabel metal2 s 30774 23222 30774 23222 4 deser_B.kept_shift_reg\[43\]
rlabel metal2 s 29394 22576 29394 22576 4 deser_B.kept_shift_reg\[44\]
rlabel metal1 s 28244 23086 28244 23086 4 deser_B.kept_shift_reg\[45\]
rlabel metal1 s 26956 22950 26956 22950 4 deser_B.kept_shift_reg\[46\]
rlabel metal1 s 26082 22202 26082 22202 4 deser_B.kept_shift_reg\[47\]
rlabel metal1 s 26082 22474 26082 22474 4 deser_B.kept_shift_reg\[48\]
rlabel metal1 s 23644 22746 23644 22746 4 deser_B.kept_shift_reg\[49\]
rlabel metal1 s 27416 31722 27416 31722 4 deser_B.kept_shift_reg\[4\]
rlabel metal2 s 22494 22644 22494 22644 4 deser_B.kept_shift_reg\[50\]
rlabel metal1 s 21850 23120 21850 23120 4 deser_B.kept_shift_reg\[51\]
rlabel metal1 s 20056 22542 20056 22542 4 deser_B.kept_shift_reg\[52\]
rlabel metal1 s 19320 23834 19320 23834 4 deser_B.kept_shift_reg\[53\]
rlabel metal1 s 20378 24650 20378 24650 4 deser_B.kept_shift_reg\[54\]
rlabel metal1 s 20240 25670 20240 25670 4 deser_B.kept_shift_reg\[55\]
rlabel metal2 s 18814 26180 18814 26180 4 deser_B.kept_shift_reg\[56\]
rlabel metal1 s 17434 26894 17434 26894 4 deser_B.kept_shift_reg\[57\]
rlabel metal1 s 16836 25466 16836 25466 4 deser_B.kept_shift_reg\[58\]
rlabel metal1 s 16192 24378 16192 24378 4 deser_B.kept_shift_reg\[59\]
rlabel metal2 s 27922 31178 27922 31178 4 deser_B.kept_shift_reg\[5\]
rlabel metal1 s 16698 23766 16698 23766 4 deser_B.kept_shift_reg\[60\]
rlabel metal1 s 17710 22066 17710 22066 4 deser_B.kept_shift_reg\[61\]
rlabel metal1 s 16468 21930 16468 21930 4 deser_B.kept_shift_reg\[62\]
rlabel metal1 s 15962 22066 15962 22066 4 deser_B.kept_shift_reg\[63\]
rlabel metal1 s 14536 22406 14536 22406 4 deser_B.kept_shift_reg\[64\]
rlabel metal2 s 13938 23494 13938 23494 4 deser_B.kept_shift_reg\[65\]
rlabel metal2 s 13938 24582 13938 24582 4 deser_B.kept_shift_reg\[66\]
rlabel metal2 s 14030 25024 14030 25024 4 deser_B.kept_shift_reg\[67\]
rlabel metal1 s 14536 26010 14536 26010 4 deser_B.kept_shift_reg\[68\]
rlabel metal2 s 14122 26860 14122 26860 4 deser_B.kept_shift_reg\[69\]
rlabel metal2 s 27646 30192 27646 30192 4 deser_B.kept_shift_reg\[6\]
rlabel metal2 s 13386 27200 13386 27200 4 deser_B.kept_shift_reg\[70\]
rlabel metal2 s 13478 27132 13478 27132 4 deser_B.kept_shift_reg\[71\]
rlabel metal1 s 13110 29274 13110 29274 4 deser_B.kept_shift_reg\[72\]
rlabel metal2 s 13202 30022 13202 30022 4 deser_B.kept_shift_reg\[73\]
rlabel metal2 s 13754 29818 13754 29818 4 deser_B.kept_shift_reg\[74\]
rlabel metal2 s 15686 29376 15686 29376 4 deser_B.kept_shift_reg\[75\]
rlabel metal2 s 15778 28968 15778 28968 4 deser_B.kept_shift_reg\[76\]
rlabel metal1 s 16698 28186 16698 28186 4 deser_B.kept_shift_reg\[77\]
rlabel metal1 s 16744 27506 16744 27506 4 deser_B.kept_shift_reg\[78\]
rlabel metal2 s 17342 28934 17342 28934 4 deser_B.kept_shift_reg\[79\]
rlabel metal1 s 27922 29478 27922 29478 4 deser_B.kept_shift_reg\[7\]
rlabel metal2 s 19918 28798 19918 28798 4 deser_B.kept_shift_reg\[80\]
rlabel metal1 s 20148 29274 20148 29274 4 deser_B.kept_shift_reg\[81\]
rlabel metal1 s 20746 29138 20746 29138 4 deser_B.kept_shift_reg\[82\]
rlabel metal2 s 22678 29002 22678 29002 4 deser_B.kept_shift_reg\[83\]
rlabel metal2 s 22586 29308 22586 29308 4 deser_B.kept_shift_reg\[84\]
rlabel metal1 s 24242 29274 24242 29274 4 deser_B.kept_shift_reg\[85\]
rlabel metal2 s 25070 29920 25070 29920 4 deser_B.kept_shift_reg\[86\]
rlabel metal2 s 26358 30634 26358 30634 4 deser_B.kept_shift_reg\[87\]
rlabel metal2 s 25806 31586 25806 31586 4 deser_B.kept_shift_reg\[88\]
rlabel metal1 s 24242 31450 24242 31450 4 deser_B.kept_shift_reg\[89\]
rlabel metal2 s 29026 28730 29026 28730 4 deser_B.kept_shift_reg\[8\]
rlabel metal1 s 23966 32878 23966 32878 4 deser_B.kept_shift_reg\[90\]
rlabel metal1 s 23414 34170 23414 34170 4 deser_B.kept_shift_reg\[91\]
rlabel metal1 s 22402 33626 22402 33626 4 deser_B.kept_shift_reg\[92\]
rlabel metal1 s 22264 32538 22264 32538 4 deser_B.kept_shift_reg\[93\]
rlabel metal2 s 22126 31042 22126 31042 4 deser_B.kept_shift_reg\[94\]
rlabel metal2 s 19642 30906 19642 30906 4 deser_B.kept_shift_reg\[95\]
rlabel metal1 s 19412 30770 19412 30770 4 deser_B.kept_shift_reg\[96\]
rlabel metal1 s 17802 30566 17802 30566 4 deser_B.kept_shift_reg\[97\]
rlabel metal2 s 17066 32198 17066 32198 4 deser_B.kept_shift_reg\[98\]
rlabel metal1 s 16560 32334 16560 32334 4 deser_B.kept_shift_reg\[99\]
rlabel metal1 s 29440 28594 29440 28594 4 deser_B.kept_shift_reg\[9\]
rlabel metal1 s 33120 31654 33120 31654 4 deser_B.receiving
rlabel metal3 s 0 25168 800 25288 4 done
port 13 nsew
rlabel metal2 s 36018 8398 36018 8398 4 net1
rlabel metal1 s 24012 28594 24012 28594 4 net10
rlabel metal1 s 26082 24752 26082 24752 4 net11
rlabel metal1 s 23506 6834 23506 6834 4 net12
rlabel metal2 s 30682 8398 30682 8398 4 net13
rlabel metal1 s 24794 6365 24794 6365 4 net14
rlabel metal2 s 22586 24514 22586 24514 4 net15
rlabel metal3 s 36754 6171 36754 6171 4 net16
rlabel metal2 s 26082 8687 26082 8687 4 net17
rlabel metal2 s 31970 16677 31970 16677 4 net18
rlabel metal2 s 19826 34238 19826 34238 4 net19
rlabel metal1 s 25024 5678 25024 5678 4 net2
rlabel metal1 s 33672 5678 33672 5678 4 net20
rlabel metal1 s 32430 3468 32430 3468 4 net21
rlabel metal1 s 22862 10676 22862 10676 4 net22
rlabel metal2 s 26266 10846 26266 10846 4 net23
rlabel metal1 s 29532 9486 29532 9486 4 net24
rlabel metal1 s 28796 13362 28796 13362 4 net25
rlabel metal1 s 32384 7174 32384 7174 4 net26
rlabel metal1 s 20516 37298 20516 37298 4 net27
rlabel metal1 s 31740 10098 31740 10098 4 net28
rlabel metal1 s 30636 10030 30636 10030 4 net29
rlabel metal1 s 32154 35530 32154 35530 4 net3
rlabel metal1 s 31280 10710 31280 10710 4 net30
rlabel metal2 s 33626 34238 33626 34238 4 net31
rlabel metal1 s 35834 34952 35834 34952 4 net32
rlabel metal1 s 33856 35190 33856 35190 4 net33
rlabel metal1 s 32798 34136 32798 34136 4 net34
rlabel metal2 s 29210 33456 29210 33456 4 net35
rlabel metal1 s 18538 33966 18538 33966 4 net36
rlabel metal2 s 32154 35632 32154 35632 4 net37
rlabel metal1 s 29532 37162 29532 37162 4 net38
rlabel metal2 s 32338 9792 32338 9792 4 net39
rlabel metal1 s 25530 36890 25530 36890 4 net4
rlabel metal1 s 21390 21012 21390 21012 4 net40
rlabel metal1 s 31372 7446 31372 7446 4 net41
rlabel metal2 s 34454 33252 34454 33252 4 net42
rlabel metal1 s 34822 32878 34822 32878 4 net43
rlabel metal1 s 31924 9622 31924 9622 4 net44
rlabel metal1 s 34776 33558 34776 33558 4 net45
rlabel metal1 s 25162 29716 25162 29716 4 net47
rlabel metal1 s 32292 4250 32292 4250 4 net490
rlabel metal2 s 32330 5338 32330 5338 4 net491
rlabel metal2 s 31142 5440 31142 5440 4 net492
rlabel metal2 s 30406 4352 30406 4352 4 net493
rlabel metal1 s 31878 4692 31878 4692 4 net494
rlabel metal2 s 30866 4930 30866 4930 4 net495
rlabel metal1 s 31924 4250 31924 4250 4 net496
rlabel metal1 s 32752 3502 32752 3502 4 net497
rlabel metal2 s 31878 37485 31878 37485 4 net499
rlabel metal1 s 2951 21930 2951 21930 4 net5
rlabel metal1 s 27048 36822 27048 36822 4 net500
rlabel metal1 s 27868 35802 27868 35802 4 net501
rlabel metal2 s 28566 36448 28566 36448 4 net502
rlabel metal2 s 28014 36652 28014 36652 4 net503
rlabel metal1 s 29624 34714 29624 34714 4 net504
rlabel metal1 s 28704 34510 28704 34510 4 net505
rlabel metal1 s 29578 32878 29578 32878 4 net506
rlabel metal1 s 34040 5746 34040 5746 4 net508
rlabel metal1 s 35098 6766 35098 6766 4 net509
rlabel metal2 s 2162 24480 2162 24480 4 net6
rlabel metal2 s 30590 25330 30590 25330 4 net640
rlabel metal2 s 24150 23902 24150 23902 4 net641
rlabel metal2 s 23506 23494 23506 23494 4 net642
rlabel metal2 s 23966 22848 23966 22848 4 net643
rlabel metal2 s 32614 32198 32614 32198 4 net644
rlabel metal2 s 32430 33082 32430 33082 4 net645
rlabel metal1 s 22908 24038 22908 24038 4 net646
rlabel metal1 s 18584 20298 18584 20298 4 net647
rlabel metal2 s 1702 14178 1702 14178 4 net7
rlabel metal1 s 25392 6766 25392 6766 4 net728
rlabel metal1 s 26910 8466 26910 8466 4 net729
rlabel metal1 s 20700 19346 20700 19346 4 net730
rlabel metal1 s 20838 14314 20838 14314 4 net731
rlabel metal2 s 17158 17782 17158 17782 4 net732
rlabel metal1 s 20470 10642 20470 10642 4 net733
rlabel metal1 s 21390 18122 21390 18122 4 net734
rlabel metal1 s 23690 5610 23690 5610 4 net735
rlabel metal2 s 30314 8466 30314 8466 4 net736
rlabel metal2 s 29670 33694 29670 33694 4 net737
rlabel metal1 s 31234 9554 31234 9554 4 net739
rlabel metal2 s 32798 15572 32798 15572 4 net740
rlabel metal1 s 34914 12206 34914 12206 4 net769
rlabel metal1 s 1748 17850 1748 17850 4 net8
rlabel metal1 s 32706 18156 32706 18156 4 net808
rlabel metal1 s 29256 8874 29256 8874 4 net809
rlabel metal2 s 29854 9724 29854 9724 4 net810
rlabel metal2 s 31786 35394 31786 35394 4 net811
rlabel metal1 s 35098 7446 35098 7446 4 net814
rlabel metal2 s 34822 35598 34822 35598 4 net816
rlabel metal2 s 34362 7548 34362 7548 4 net818
rlabel metal1 s 32384 31314 32384 31314 4 net820
rlabel metal1 s 32982 32470 32982 32470 4 net821
rlabel metal1 s 18814 36686 18814 36686 4 net845
rlabel metal3 s 32798 35547 32798 35547 4 net846
rlabel metal1 s 18906 37740 18906 37740 4 net847
rlabel metal2 s 32798 35853 32798 35853 4 net848
rlabel metal1 s 1518 24922 1518 24922 4 net9
rlabel metal3 s 0 36728 800 36848 4 rst_n
port 14 nsew
rlabel metal1 s 2438 14246 2438 14246 4 ser_C.bit_idx\[0\]
rlabel metal1 s 3220 14314 3220 14314 4 ser_C.bit_idx\[1\]
rlabel metal2 s 4094 15742 4094 15742 4 ser_C.bit_idx\[2\]
rlabel metal1 s 3542 17238 3542 17238 4 ser_C.bit_idx\[3\]
rlabel metal1 s 4508 17578 4508 17578 4 ser_C.bit_idx\[4\]
rlabel metal2 s 5290 17136 5290 17136 4 ser_C.bit_idx\[5\]
rlabel metal1 s 4186 18088 4186 18088 4 ser_C.bit_idx\[6\]
rlabel metal1 s 3542 19754 3542 19754 4 ser_C.bit_idx\[7\]
rlabel metal1 s 3956 19142 3956 19142 4 ser_C.bit_idx\[8\]
rlabel metal2 s 3174 18428 3174 18428 4 ser_C.bit_idx\[9\]
rlabel metal2 s 6762 14722 6762 14722 4 ser_C.kept_bit_idx\[0\]
rlabel metal1 s 5750 13872 5750 13872 4 ser_C.kept_bit_idx\[1\]
rlabel metal1 s 8372 14994 8372 14994 4 ser_C.kept_bit_idx\[2\]
rlabel metal1 s 10534 14926 10534 14926 4 ser_C.kept_bit_idx\[3\]
rlabel metal2 s 10810 14756 10810 14756 4 ser_C.kept_bit_idx\[4\]
rlabel metal2 s 10626 15164 10626 15164 4 ser_C.kept_bit_idx\[5\]
rlabel metal2 s 11086 17136 11086 17136 4 ser_C.kept_bit_idx\[6\]
rlabel metal1 s 11316 17646 11316 17646 4 ser_C.kept_bit_idx\[7\]
rlabel metal2 s 9522 16830 9522 16830 4 ser_C.kept_bit_idx\[8\]
rlabel metal2 s 7498 17340 7498 17340 4 ser_C.kept_bit_idx\[9\]
rlabel metal3 s 0 23808 800 23928 4 start
port 15 nsew
rlabel metal1 s 2346 25364 2346 25364 4 systolic_inst.ce_local
rlabel metal2 s 3174 26588 3174 26588 4 systolic_inst.cycle_cnt\[0\]
rlabel metal2 s 5750 25534 5750 25534 4 systolic_inst.cycle_cnt\[10\]
rlabel metal2 s 6394 24276 6394 24276 4 systolic_inst.cycle_cnt\[11\]
rlabel metal1 s 5658 22032 5658 22032 4 systolic_inst.cycle_cnt\[12\]
rlabel metal1 s 4508 22066 4508 22066 4 systolic_inst.cycle_cnt\[13\]
rlabel metal1 s 4416 21318 4416 21318 4 systolic_inst.cycle_cnt\[14\]
rlabel metal1 s 5382 21896 5382 21896 4 systolic_inst.cycle_cnt\[15\]
rlabel metal2 s 9338 21386 9338 21386 4 systolic_inst.cycle_cnt\[16\]
rlabel metal1 s 8004 20026 8004 20026 4 systolic_inst.cycle_cnt\[17\]
rlabel metal2 s 8786 19652 8786 19652 4 systolic_inst.cycle_cnt\[18\]
rlabel metal1 s 9522 20910 9522 20910 4 systolic_inst.cycle_cnt\[19\]
rlabel metal1 s 2714 28084 2714 28084 4 systolic_inst.cycle_cnt\[1\]
rlabel metal2 s 10810 21284 10810 21284 4 systolic_inst.cycle_cnt\[20\]
rlabel metal1 s 11408 22066 11408 22066 4 systolic_inst.cycle_cnt\[21\]
rlabel metal2 s 10902 22780 10902 22780 4 systolic_inst.cycle_cnt\[22\]
rlabel metal2 s 8786 23494 8786 23494 4 systolic_inst.cycle_cnt\[23\]
rlabel metal2 s 9706 26180 9706 26180 4 systolic_inst.cycle_cnt\[24\]
rlabel metal1 s 11638 25874 11638 25874 4 systolic_inst.cycle_cnt\[25\]
rlabel metal1 s 10810 26996 10810 26996 4 systolic_inst.cycle_cnt\[26\]
rlabel metal1 s 10718 26758 10718 26758 4 systolic_inst.cycle_cnt\[27\]
rlabel metal1 s 9292 29002 9292 29002 4 systolic_inst.cycle_cnt\[28\]
rlabel metal1 s 9430 30362 9430 30362 4 systolic_inst.cycle_cnt\[29\]
rlabel metal1 s 3910 29240 3910 29240 4 systolic_inst.cycle_cnt\[2\]
rlabel metal1 s 9522 30294 9522 30294 4 systolic_inst.cycle_cnt\[30\]
rlabel metal2 s 10626 29308 10626 29308 4 systolic_inst.cycle_cnt\[31\]
rlabel metal1 s 3864 28934 3864 28934 4 systolic_inst.cycle_cnt\[3\]
rlabel metal1 s 4608 28390 4608 28390 4 systolic_inst.cycle_cnt\[4\]
rlabel metal1 s 6072 29138 6072 29138 4 systolic_inst.cycle_cnt\[5\]
rlabel metal1 s 6946 30124 6946 30124 4 systolic_inst.cycle_cnt\[6\]
rlabel metal2 s 5750 28288 5750 28288 4 systolic_inst.cycle_cnt\[7\]
rlabel metal1 s 7222 25228 7222 25228 4 systolic_inst.cycle_cnt\[8\]
rlabel metal2 s 5934 26724 5934 26724 4 systolic_inst.cycle_cnt\[9\]
flabel metal3 s 37408 16328 38208 16448 0 FreeSans 600 0 0 0 A_in_frame_sync
port 1 nsew
flabel metal2 s 10322 0 10378 800 0 FreeSans 280 90 0 0 A_in_serial_clk
port 2 nsew
flabel metal2 s 23202 0 23258 800 0 FreeSans 280 90 0 0 A_in_serial_data
port 3 nsew
flabel metal2 s 29642 39552 29698 40352 0 FreeSans 280 90 0 0 B_in_frame_sync
port 4 nsew
flabel metal2 s 30930 39552 30986 40352 0 FreeSans 280 90 0 0 B_in_serial_clk
port 5 nsew
flabel metal2 s 25134 39552 25190 40352 0 FreeSans 280 90 0 0 B_in_serial_data
port 6 nsew
flabel metal3 s 0 14288 800 14408 0 FreeSans 600 0 0 0 C_out_frame_sync
port 7 nsew
flabel metal3 s 0 17688 800 17808 0 FreeSans 600 0 0 0 C_out_serial_clk
port 8 nsew
flabel metal3 s 37408 6128 38208 6248 0 FreeSans 600 0 0 0 C_out_serial_data
port 9 nsew
flabel metal5 s 1056 36642 37124 36962 0 FreeSans 3200 0 0 0 VGND
port 10 nsew
flabel metal5 s 1056 6006 37124 6326 0 FreeSans 3200 0 0 0 VGND
port 10 nsew
flabel metal4 s 35588 2128 35908 38128 0 FreeSans 2400 90 0 0 VGND
port 10 nsew
flabel metal4 s 4868 2128 5188 38128 0 FreeSans 2400 90 0 0 VGND
port 10 nsew
flabel metal5 s 1056 35982 37124 36302 0 FreeSans 3200 0 0 0 VPWR
port 11 nsew
flabel metal5 s 1056 5346 37124 5666 0 FreeSans 3200 0 0 0 VPWR
port 11 nsew
flabel metal4 s 34928 2128 35248 38128 0 FreeSans 2400 90 0 0 VPWR
port 11 nsew
flabel metal4 s 4208 2128 4528 38128 0 FreeSans 2400 90 0 0 VPWR
port 11 nsew
flabel metal3 s 0 29248 800 29368 0 FreeSans 600 0 0 0 clk
port 12 nsew
flabel metal3 s 400 25228 400 25228 0 FreeSans 600 0 0 0 done
flabel metal3 s 400 36788 400 36788 0 FreeSans 600 0 0 0 rst_n
flabel metal3 s 400 23868 400 23868 0 FreeSans 600 0 0 0 start
<< properties >>
string FIXED_BBOX 0 0 38208 40352
<< end >>
