* NGSPICE file created from Systolic4x4_serial_io.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

.subckt Systolic4x4_serial_io A_in_frame_sync A_in_serial_clk A_in_serial_data B_in_frame_sync
+ B_in_serial_clk B_in_serial_data C_out_frame_sync C_out_serial_clk C_out_serial_data
+ VGND VPWR clk done rst_n start
XFILLER_228_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_199_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18869_ _05977_ _05978_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__nand2_1
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20900_ _07774_ _07775_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__or2_1
X_21880_ _08677_ _08678_ _08670_ _08673_ VGND VGND VPWR VPWR _08679_ sky130_fd_sc_hd__a211o_1
XFILLER_55_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20831_ systolic_inst.A_outs\[4\]\[4\] systolic_inst.A_shift\[8\]\[4\] net121 VGND
+ VGND VPWR VPWR _01654_ sky130_fd_sc_hd__mux2_1
XFILLER_242_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20762_ _07660_ _07666_ _07667_ net60 VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__a31o_1
X_23550_ _10130_ _10132_ _10171_ VGND VGND VPWR VPWR _10173_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22501_ _09226_ _09227_ _09225_ VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__a21bo_1
XFILLER_196_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23481_ _10073_ _10075_ _10074_ VGND VGND VPWR VPWR _10105_ sky130_fd_sc_hd__o21ba_1
XFILLER_211_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20693_ _07603_ _07605_ _07601_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__a21bo_1
XFILLER_51_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22432_ _09170_ _09171_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__nor2_1
XFILLER_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25220_ net110 ser_C.shift_reg\[438\] VGND VGND VPWR VPWR _11080_ sky130_fd_sc_hd__and2_1
XFILLER_91_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22363_ _09096_ _09104_ VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__nand2_1
XFILLER_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25151_ C_out\[402\] net101 net73 ser_C.shift_reg\[402\] _11045_ VGND VGND VPWR VPWR
+ _02652_ sky130_fd_sc_hd__a221o_1
XFILLER_148_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24102_ _10560_ systolic_inst.B_shift\[19\]\[6\] net71 VGND VGND VPWR VPWR _02088_
+ sky130_fd_sc_hd__mux2_1
X_21314_ net63 _08168_ _08169_ systolic_inst.acc_wires\[4\]\[9\] net108 VGND VGND
+ VPWR VPWR _01691_ sky130_fd_sc_hd__a32o_1
X_25082_ net112 ser_C.shift_reg\[369\] VGND VGND VPWR VPWR _11011_ sky130_fd_sc_hd__and2_1
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22294_ _09029_ _09037_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24033_ systolic_inst.B_shift\[8\]\[4\] B_in\[36\] _00008_ VGND VGND VPWR VPWR _10534_
+ sky130_fd_sc_hd__mux2_1
X_28910_ clknet_leaf_281_clk _02708_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[458\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21245_ _08074_ _08093_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__xor2_1
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28841_ clknet_leaf_333_clk _02639_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[389\]
+ sky130_fd_sc_hd__dfrtp_1
X_21176_ _08000_ _08010_ _08008_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__a21o_1
XFILLER_172_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20127_ net60 _07103_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__nor2_1
XFILLER_132_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28772_ clknet_leaf_295_clk _02570_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[320\]
+ sky130_fd_sc_hd__dfrtp_1
X_25984_ systolic_inst.acc_wires\[14\]\[12\] ser_C.parallel_data\[460\] net26 VGND
+ VGND VPWR VPWR _03286_ sky130_fd_sc_hd__mux2_1
XFILLER_218_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27723_ clknet_leaf_190_clk _01521_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_20058_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[6\]\[7\]
+ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__nand2_1
X_24935_ C_out\[294\] net102 net76 ser_C.shift_reg\[294\] _10937_ VGND VGND VPWR VPWR
+ _02544_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27654_ clknet_leaf_303_clk _01452_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_24866_ net110 ser_C.shift_reg\[261\] VGND VGND VPWR VPWR _10903_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26605_ clknet_leaf_16_B_in_serial_clk _00408_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_23817_ _11258_ systolic_inst.acc_wires\[0\]\[18\] net64 _10415_ VGND VGND VPWR VPWR
+ _01948_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27585_ clknet_leaf_216_clk _01383_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_27_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24797_ C_out\[225\] net99 net79 ser_C.shift_reg\[225\] _10868_ VGND VGND VPWR VPWR
+ _02475_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29324_ clknet_leaf_304_clk _03122_ net138 VGND VGND VPWR VPWR C_out\[296\] sky130_fd_sc_hd__dfrtp_1
XFILLER_199_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14550_ _11721_ _11722_ _11723_ VGND VGND VPWR VPWR _11725_ sky130_fd_sc_hd__and3_1
X_26536_ clknet_leaf_21_A_in_serial_clk _00339_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_23748_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[0\]\[8\]
+ _10353_ _10355_ VGND VGND VPWR VPWR _10356_ sky130_fd_sc_hd__a211o_1
XFILLER_148_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13501_ deser_A.shift_reg\[65\] deser_A.shift_reg\[66\] net129 VGND VGND VPWR VPWR
+ _00338_ sky130_fd_sc_hd__mux2_1
XFILLER_199_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29255_ clknet_leaf_197_clk _03053_ net147 VGND VGND VPWR VPWR C_out\[227\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26467_ clknet_leaf_346_clk deser_A.serial_toggle_sync1 net132 VGND VGND VPWR VPWR
+ deser_A.serial_toggle_sync2 sky130_fd_sc_hd__dfrtp_2
X_14481_ _11593_ _11630_ _11629_ VGND VGND VPWR VPWR _11662_ sky130_fd_sc_hd__a21bo_1
XFILLER_202_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23679_ _10274_ _10276_ VGND VGND VPWR VPWR _10298_ sky130_fd_sc_hd__nor2_1
XFILLER_109_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28206_ clknet_leaf_94_clk _02004_ VGND VGND VPWR VPWR systolic_inst.B_shift\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_23_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _03602_ _03601_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__nand2b_1
XFILLER_70_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25418_ _11178_ systolic_inst.A_shift\[0\]\[0\] net71 VGND VGND VPWR VPWR _02786_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13432_ _11316_ VGND VGND VPWR VPWR _11317_ sky130_fd_sc_hd__inv_2
X_29186_ clknet_leaf_133_clk _02984_ net142 VGND VGND VPWR VPWR C_out\[158\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26398_ clknet_leaf_31_clk _00205_ net137 VGND VGND VPWR VPWR A_in\[66\] sky130_fd_sc_hd__dfrtp_1
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28137_ clknet_leaf_126_clk _01935_ net144 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16151_ _03526_ _03534_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__xnor2_1
X_25349_ ser_C.parallel_data\[501\] net98 net78 ser_C.shift_reg\[501\] _11144_ VGND
+ VGND VPWR VPWR _02751_ sky130_fd_sc_hd__a221o_1
X_13363_ A_in\[72\] deser_A.word_buffer\[72\] net94 VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__mux2_1
XFILLER_220_1169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15102_ _12216_ _12217_ VGND VGND VPWR VPWR _12219_ sky130_fd_sc_hd__xor2_1
X_28068_ clknet_leaf_120_clk _01866_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_16082_ _13031_ _13033_ _13076_ VGND VGND VPWR VPWR _13078_ sky130_fd_sc_hd__and3_1
X_13294_ A_in\[3\] deser_A.word_buffer\[3\] net94 VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__mux2_1
XFILLER_142_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19910_ _06906_ _06907_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__nand2_1
XFILLER_142_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27019_ clknet_leaf_23_B_in_serial_clk _00817_ net137 VGND VGND VPWR VPWR deser_B.shift_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_15033_ _12112_ _12114_ _12113_ VGND VGND VPWR VPWR _12152_ sky130_fd_sc_hd__o21ba_1
XFILLER_108_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19841_ _06839_ _06840_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__nand2_1
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19772_ _06741_ _06773_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__and2b_1
XFILLER_7_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16984_ _04294_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15935_ systolic_inst.acc_wires\[13\]\[26\] systolic_inst.acc_wires\[13\]\[27\] systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12957_ sky130_fd_sc_hd__o21a_1
X_18723_ _05835_ _05847_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__xor2_1
XFILLER_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18654_ _05779_ _05780_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__nand2_1
XFILLER_236_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15866_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[17\]
+ VGND VGND VPWR VPWR _12899_ sky130_fd_sc_hd__xor2_2
XFILLER_188_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_B_in_serial_clk clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_23_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
Xwire29 net30 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_8
XFILLER_40_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14817_ systolic_inst.A_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[5\] VGND VGND
+ VPWR VPWR _11942_ sky130_fd_sc_hd__nand2_1
XFILLER_64_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17605_ _11712_ _04848_ _04849_ systolic_inst.acc_wires\[10\]\[4\] net107 VGND VGND
+ VPWR VPWR _01302_ sky130_fd_sc_hd__a32o_1
XFILLER_236_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18585_ _05639_ _05674_ _05676_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_194_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _12833_ _12834_ _12832_ VGND VGND VPWR VPWR _12840_ sky130_fd_sc_hd__a21bo_1
X_17536_ _04785_ _04786_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__and2b_1
X_14748_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[9\]\[0\] net115 VGND
+ VGND VPWR VPWR _01018_ sky130_fd_sc_hd__mux2_1
XFILLER_75_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_190_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17467_ _04720_ _04719_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__nand2b_1
XFILLER_225_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14679_ _11826_ _11827_ VGND VGND VPWR VPWR _11835_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_211_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19206_ _06269_ _06270_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__xor2_1
X_16418_ _03784_ _03785_ net67 VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17398_ _04653_ _04652_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__nand2b_1
XFILLER_203_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19137_ _06201_ _06202_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__nand2_1
X_16349_ _03659_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19068_ _06129_ _06135_ _06136_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__and3_1
XFILLER_118_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18019_ _05208_ _05209_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_209_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21030_ _07902_ _07901_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_147_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22981_ systolic_inst.A_outs\[1\]\[5\] systolic_inst.B_outs\[1\]\[6\] systolic_inst.A_outs\[1\]\[6\]
+ systolic_inst.B_outs\[1\]\[7\] VGND VGND VPWR VPWR _09658_ sky130_fd_sc_hd__and4b_1
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24720_ net113 ser_C.shift_reg\[188\] VGND VGND VPWR VPWR _10830_ sky130_fd_sc_hd__and2_1
X_21932_ _08720_ _08722_ VGND VGND VPWR VPWR _08723_ sky130_fd_sc_hd__or2_1
XFILLER_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24651_ C_out\[152\] net104 _10643_ ser_C.shift_reg\[152\] _10795_ VGND VGND VPWR
+ VPWR _02402_ sky130_fd_sc_hd__a221o_1
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21863_ _08663_ _08664_ VGND VGND VPWR VPWR _08665_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_156_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23602_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[5\] _10222_ VGND
+ VGND VPWR VPWR _10223_ sky130_fd_sc_hd__a21o_1
XFILLER_230_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20814_ net106 systolic_inst.acc_wires\[5\]\[29\] net68 _07713_ VGND VGND VPWR VPWR
+ _01647_ sky130_fd_sc_hd__a22o_1
X_27370_ clknet_leaf_339_clk _01168_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24582_ net114 ser_C.shift_reg\[119\] VGND VGND VPWR VPWR _10761_ sky130_fd_sc_hd__and2_1
X_21794_ _08597_ _08598_ VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__nand2_1
XFILLER_196_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26321_ clknet_leaf_0_A_in_serial_clk _00129_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_23533_ systolic_inst.A_outs\[0\]\[4\] systolic_inst.B_outs\[0\]\[6\] _10155_ VGND
+ VGND VPWR VPWR _10156_ sky130_fd_sc_hd__and3_1
XFILLER_54_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20745_ net106 systolic_inst.acc_wires\[5\]\[18\] net68 _07655_ VGND VGND VPWR VPWR
+ _01636_ sky130_fd_sc_hd__a22o_1
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29040_ clknet_leaf_122_clk _02838_ net152 VGND VGND VPWR VPWR C_out\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_196_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26252_ clknet_leaf_10_A_in_serial_clk _00060_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_23464_ _10044_ _10047_ _10088_ VGND VGND VPWR VPWR _10089_ sky130_fd_sc_hd__a21o_1
XFILLER_149_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20676_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[5\]\[8\]
+ _07593_ _07595_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__a211o_1
XFILLER_195_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25203_ C_out\[428\] net101 net73 ser_C.shift_reg\[428\] _11071_ VGND VGND VPWR VPWR
+ _02678_ sky130_fd_sc_hd__a221o_1
XFILLER_104_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22415_ systolic_inst.A_outs\[2\]\[6\] _11265_ VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__nor2_1
X_26183_ ser_C.bit_idx\[4\] _11303_ _11247_ ser_C.bit_idx\[3\] VGND VGND VPWR VPWR
+ _11251_ sky130_fd_sc_hd__a22oi_1
XFILLER_183_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23395_ _09986_ _09988_ _10020_ VGND VGND VPWR VPWR _10022_ sky130_fd_sc_hd__and3_1
XFILLER_137_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25134_ net110 ser_C.shift_reg\[395\] VGND VGND VPWR VPWR _11037_ sky130_fd_sc_hd__and2_1
XFILLER_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22346_ _09086_ _09087_ VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__xor2_1
XFILLER_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22277_ _08991_ _08993_ _08990_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__o21ba_1
XFILLER_136_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25065_ C_out\[359\] net97 net77 ser_C.shift_reg\[359\] _11002_ VGND VGND VPWR VPWR
+ _02609_ sky130_fd_sc_hd__a221o_1
XFILLER_88_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24016_ systolic_inst.B_shift\[7\]\[7\] _11332_ net83 systolic_inst.B_shift\[11\]\[7\]
+ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__a22o_1
X_21228_ _08063_ _08064_ _08066_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__o21ba_1
XFILLER_105_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21159_ _07992_ _08027_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__nor2_1
X_28824_ clknet_leaf_239_clk _02622_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[372\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_1260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28755_ clknet_leaf_220_clk _02553_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[303\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13981_ deser_B.shift_reg\[15\] deser_B.shift_reg\[16\] net125 VGND VGND VPWR VPWR
+ _00807_ sky130_fd_sc_hd__mux2_1
X_25967_ systolic_inst.acc_wires\[13\]\[27\] ser_C.parallel_data\[443\] net19 VGND
+ VGND VPWR VPWR _03269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27706_ clknet_leaf_190_clk _01504_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_15720_ _11272_ systolic_inst.A_outs\[13\]\[7\] _12720_ _12746_ VGND VGND VPWR VPWR
+ _12772_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_66_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24918_ net110 ser_C.shift_reg\[287\] VGND VGND VPWR VPWR _10929_ sky130_fd_sc_hd__and2_1
XFILLER_218_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28686_ clknet_leaf_192_clk _02484_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[234\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25898_ systolic_inst.acc_wires\[11\]\[22\] C_out\[374\] net41 VGND VGND VPWR VPWR
+ _03200_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_215_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _12644_ _12705_ VGND VGND VPWR VPWR _12706_ sky130_fd_sc_hd__xnor2_1
X_27637_ clknet_leaf_315_clk _01435_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24849_ C_out\[251\] net98 net78 ser_C.shift_reg\[251\] _10894_ VGND VGND VPWR VPWR
+ _02501_ sky130_fd_sc_hd__a221o_1
XFILLER_209_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14602_ _11767_ _11768_ VGND VGND VPWR VPWR _11769_ sky130_fd_sc_hd__nand2_1
XFILLER_233_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18370_ _05520_ _05522_ _05528_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_17_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15582_ _12637_ _12610_ VGND VGND VPWR VPWR _12639_ sky130_fd_sc_hd__and2b_1
X_27568_ clknet_leaf_298_clk _01366_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29307_ clknet_leaf_313_clk _03105_ net141 VGND VGND VPWR VPWR C_out\[279\] sky130_fd_sc_hd__dfrtp_1
X_17321_ systolic_inst.A_outs\[10\]\[1\] systolic_inst.B_outs\[10\]\[6\] _04578_ VGND
+ VGND VPWR VPWR _04579_ sky130_fd_sc_hd__and3_1
XFILLER_159_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14533_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[15\]\[0\]
+ _11708_ _11709_ VGND VGND VPWR VPWR _11710_ sky130_fd_sc_hd__and4_1
XFILLER_14_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26519_ clknet_leaf_10_A_in_serial_clk _00322_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27499_ clknet_leaf_225_clk _01297_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29238_ clknet_leaf_179_clk _03036_ net148 VGND VGND VPWR VPWR C_out\[210\] sky130_fd_sc_hd__dfrtp_1
XFILLER_187_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17252_ systolic_inst.A_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[5\] VGND VGND
+ VPWR VPWR _04512_ sky130_fd_sc_hd__nand2_1
XFILLER_159_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14464_ _11580_ _11584_ _11613_ _11615_ VGND VGND VPWR VPWR _11646_ sky130_fd_sc_hd__o31a_1
X_16203_ _03547_ _03551_ _03585_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__or3_1
XFILLER_31_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13415_ A_in\[124\] deser_A.word_buffer\[124\] net92 VGND VGND VPWR VPWR _00263_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29169_ clknet_leaf_43_clk _02967_ net142 VGND VGND VPWR VPWR C_out\[141\] sky130_fd_sc_hd__dfrtp_1
XFILLER_70_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17183_ systolic_inst.A_outs\[10\]\[5\] systolic_inst.A_outs\[9\]\[5\] net120 VGND
+ VGND VPWR VPWR _01271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14395_ _11552_ _11577_ VGND VGND VPWR VPWR _11579_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_42_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16134_ _03518_ _03515_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__and2b_1
XFILLER_6_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13346_ A_in\[55\] deser_A.word_buffer\[55\] net92 VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__mux2_1
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16065_ _13029_ _13059_ VGND VGND VPWR VPWR _13061_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_19_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13277_ deser_A.word_buffer\[115\] deser_A.serial_word\[115\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__mux2_1
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15016_ _12061_ _12067_ _12099_ _12097_ VGND VGND VPWR VPWR _12136_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_55_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_204_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19824_ _06822_ _06823_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__or2_1
XFILLER_150_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19755_ systolic_inst.A_outs\[6\]\[2\] systolic_inst.B_outs\[6\]\[5\] VGND VGND VPWR
+ VPWR _06757_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_196_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16967_ net119 _04270_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_196_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18706_ net117 _05829_ _05830_ _05831_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__a31o_1
X_15918_ _12943_ _12942_ systolic_inst.acc_wires\[13\]\[24\] net108 VGND VGND VPWR
+ VPWR _01130_ sky130_fd_sc_hd__a2bb2o_1
X_19686_ _06685_ _06688_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__xnor2_1
X_16898_ _04214_ _04213_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_192_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15849_ _12881_ _12884_ VGND VGND VPWR VPWR _12885_ sky130_fd_sc_hd__nand2_1
XFILLER_52_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18637_ _05695_ _05763_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__nor2_1
XFILLER_64_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18568_ _05696_ _05693_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__and2b_1
XFILLER_224_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17519_ systolic_inst.B_outs\[10\]\[6\] systolic_inst.A_outs\[10\]\[7\] VGND VGND
+ VPWR VPWR _04771_ sky130_fd_sc_hd__nand2_1
X_18499_ _05629_ _05626_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__and2b_1
XFILLER_240_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20530_ _07323_ _07461_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__nand2_1
XFILLER_138_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20461_ _07394_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__or2_1
XFILLER_193_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22200_ _08894_ _08921_ _08920_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__a21oi_1
X_23180_ _09835_ _09836_ VGND VGND VPWR VPWR _09837_ sky130_fd_sc_hd__nand2_1
XFILLER_238_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20392_ systolic_inst.B_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[5\]
+ systolic_inst.B_outs\[5\]\[3\] VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_149_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22131_ _08860_ _08877_ _08879_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_149_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22062_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[29\]
+ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_145_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21013_ systolic_inst.A_outs\[4\]\[3\] _07884_ _07885_ VGND VGND VPWR VPWR _07886_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26870_ clknet_leaf_14_A_in_serial_clk _00668_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25821_ systolic_inst.acc_wires\[9\]\[9\] C_out\[297\] net15 VGND VGND VPWR VPWR
+ _03123_ sky130_fd_sc_hd__mux2_1
XFILLER_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28540_ clknet_leaf_159_clk _02338_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_228_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25752_ systolic_inst.acc_wires\[7\]\[4\] C_out\[228\] net40 VGND VGND VPWR VPWR
+ _03054_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22964_ _09588_ _09606_ _09605_ VGND VGND VPWR VPWR _09642_ sky130_fd_sc_hd__o21a_1
XFILLER_74_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24703_ C_out\[178\] net99 net79 ser_C.shift_reg\[178\] _10821_ VGND VGND VPWR VPWR
+ _02428_ sky130_fd_sc_hd__a221o_1
X_28471_ clknet_leaf_102_clk _02269_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_21915_ _08701_ _08704_ _08706_ _08707_ VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__o211ai_2
X_25683_ systolic_inst.acc_wires\[4\]\[31\] C_out\[159\] net31 VGND VGND VPWR VPWR
+ _02985_ sky130_fd_sc_hd__mux2_1
XFILLER_82_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22895_ _09573_ _09574_ VGND VGND VPWR VPWR _09575_ sky130_fd_sc_hd__and2_1
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27422_ clknet_leaf_248_clk _01220_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24634_ net7 ser_C.shift_reg\[145\] VGND VGND VPWR VPWR _10787_ sky130_fd_sc_hd__and2_1
XFILLER_203_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21846_ _08585_ _08648_ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27353_ clknet_leaf_233_clk _01151_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_24565_ C_out\[109\] net100 net80 ser_C.shift_reg\[109\] _10752_ VGND VGND VPWR VPWR
+ _02359_ sky130_fd_sc_hd__a221o_1
XFILLER_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21777_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[7\] _08554_ _08519_
+ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__a31o_1
XFILLER_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26304_ clknet_leaf_23_A_in_serial_clk _00112_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_208_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23516_ _10138_ _10139_ VGND VGND VPWR VPWR _10140_ sky130_fd_sc_hd__and2b_1
XFILLER_212_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20728_ _07639_ _07640_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__and2_1
X_27284_ clknet_leaf_320_clk _01082_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_24496_ net113 ser_C.shift_reg\[76\] VGND VGND VPWR VPWR _10718_ sky130_fd_sc_hd__and2_1
XFILLER_156_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29023_ clknet_leaf_93_clk _02821_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_221_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26235_ clknet_leaf_15_A_in_serial_clk _00043_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23447_ _10064_ _10070_ VGND VGND VPWR VPWR _10072_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20659_ _07575_ _07576_ _07574_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__a21bo_1
XFILLER_17_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ deser_A.word_buffer\[38\] deser_A.serial_word\[38\] net127 VGND VGND VPWR
+ VPWR _00048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26166_ deser_B.serial_word\[121\] deser_B.shift_reg\[121\] net56 VGND VGND VPWR
+ VPWR _03468_ sky130_fd_sc_hd__mux2_1
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14180_ _11364_ _11369_ VGND VGND VPWR VPWR _11370_ sky130_fd_sc_hd__and2b_1
X_23378_ _10003_ _10004_ _09975_ VGND VGND VPWR VPWR _10005_ sky130_fd_sc_hd__or3b_1
XFILLER_109_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13131_ _11284_ VGND VGND VPWR VPWR _11285_ sky130_fd_sc_hd__inv_2
XFILLER_139_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25117_ C_out\[385\] net101 net73 ser_C.shift_reg\[385\] _11028_ VGND VGND VPWR VPWR
+ _02635_ sky130_fd_sc_hd__a221o_1
X_22329_ _09062_ _09070_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__or2_1
XFILLER_139_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26097_ deser_B.serial_word\[52\] deser_B.shift_reg\[52\] net56 VGND VGND VPWR VPWR
+ _03399_ sky130_fd_sc_hd__mux2_1
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_240_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25048_ net112 ser_C.shift_reg\[352\] VGND VGND VPWR VPWR _10994_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_240_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_240_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17870_ _05059_ _05064_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__xor2_1
XFILLER_239_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28807_ clknet_leaf_245_clk _02605_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[355\]
+ sky130_fd_sc_hd__dfrtp_1
X_16821_ _04102_ _04104_ _04103_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__o21ba_1
XFILLER_232_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26999_ clknet_leaf_16_B_in_serial_clk _00797_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19540_ systolic_inst.acc_wires\[7\]\[16\] systolic_inst.acc_wires\[7\]\[17\] systolic_inst.acc_wires\[7\]\[18\]
+ systolic_inst.acc_wires\[7\]\[19\] systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_89_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16752_ _04071_ _04072_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__and2_1
X_28738_ clknet_leaf_301_clk _02536_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[286\]
+ sky130_fd_sc_hd__dfrtp_1
X_13964_ deser_A.serial_word\[125\] deser_A.shift_reg\[125\] _00002_ VGND VGND VPWR
+ VPWR _00790_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15703_ _12754_ _12755_ VGND VGND VPWR VPWR _12756_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_238_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_238_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28669_ clknet_leaf_187_clk _02467_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[217\]
+ sky130_fd_sc_hd__dfrtp_1
X_19471_ _06515_ _06517_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16683_ _04003_ _04004_ _03975_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__a21oi_1
XFILLER_234_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13895_ deser_A.serial_word\[56\] deser_A.shift_reg\[56\] net58 VGND VGND VPWR VPWR
+ _00721_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15634_ systolic_inst.A_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[5\] systolic_inst.B_outs\[13\]\[6\]
+ systolic_inst.B_outs\[13\]\[7\] VGND VGND VPWR VPWR _12689_ sky130_fd_sc_hd__and4b_1
X_18422_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[1\]
+ systolic_inst.B_outs\[8\]\[0\] VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__a22o_1
XFILLER_179_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_234_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18353_ _05467_ _05468_ _05493_ _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__a211o_1
XFILLER_203_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15565_ systolic_inst.A_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[6\]
+ systolic_inst.B_outs\[13\]\[7\] VGND VGND VPWR VPWR _12622_ sky130_fd_sc_hd__and4b_1
XFILLER_72_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _04530_ _04553_ _04552_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__a21boi_1
XFILLER_30_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _11643_ _11671_ _11672_ VGND VGND VPWR VPWR _11696_ sky130_fd_sc_hd__a21bo_1
XFILLER_202_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18284_ _05455_ _05453_ systolic_inst.acc_wires\[9\]\[13\] net107 VGND VGND VPWR
+ VPWR _01375_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_226_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15496_ _12520_ _12553_ VGND VGND VPWR VPWR _12555_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17235_ _04489_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__nor2_1
X_14447_ _11628_ _11627_ VGND VGND VPWR VPWR _11629_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17166_ systolic_inst.acc_wires\[11\]\[28\] systolic_inst.acc_wires\[11\]\[29\] systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__o21ai_1
XFILLER_190_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14378_ systolic_inst.A_outs\[15\]\[3\] systolic_inst.A_outs\[15\]\[4\] systolic_inst.B_outs\[15\]\[6\]
+ systolic_inst.B_outs\[15\]\[7\] VGND VGND VPWR VPWR _11562_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_185_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16117_ _13060_ _13061_ _13074_ _13073_ _13041_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__o32a_1
XFILLER_6_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13329_ A_in\[38\] deser_A.word_buffer\[38\] net94 VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__mux2_1
XFILLER_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17097_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[19\]
+ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16048_ _13034_ _13042_ VGND VGND VPWR VPWR _13045_ sky130_fd_sc_hd__and2_1
XFILLER_83_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19807_ _06807_ _06806_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_140_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17999_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[7\] VGND VGND VPWR
+ VPWR _05191_ sky130_fd_sc_hd__nand2_4
XFILLER_211_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19738_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[6\] _06738_
+ _06740_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__a22o_1
XFILLER_38_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_239_Right_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19669_ _06654_ _06672_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21700_ _08468_ _08470_ _08506_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__and3_1
XFILLER_240_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22680_ systolic_inst.A_outs\[1\]\[7\] systolic_inst.A_outs\[0\]\[7\] net121 VGND
+ VGND VPWR VPWR _01849_ sky130_fd_sc_hd__mux2_1
XFILLER_53_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21631_ systolic_inst.B_outs\[3\]\[7\] _08405_ _08406_ VGND VGND VPWR VPWR _08440_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24350_ net7 ser_C.shift_reg\[3\] VGND VGND VPWR VPWR _10645_ sky130_fd_sc_hd__and2_1
X_21562_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[3\] _08357_ _08356_
+ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__a31o_1
XFILLER_193_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23301_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\]
+ systolic_inst.A_outs\[0\]\[2\] VGND VGND VPWR VPWR _09931_ sky130_fd_sc_hd__nand4_1
X_20513_ _07407_ _07409_ _07445_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__nand3_1
XFILLER_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21493_ _08306_ _08307_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__nand2_1
X_24281_ systolic_inst.B_shift\[27\]\[4\] B_in\[92\] _00008_ VGND VGND VPWR VPWR _10614_
+ sky130_fd_sc_hd__mux2_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26020_ systolic_inst.acc_wires\[15\]\[16\] ser_C.parallel_data\[496\] net23 VGND
+ VGND VPWR VPWR _03322_ sky130_fd_sc_hd__mux2_1
X_23232_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[24\]
+ VGND VGND VPWR VPWR _09881_ sky130_fd_sc_hd__and2_1
XFILLER_181_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20444_ _07363_ _07379_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__or2_1
XFILLER_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23163_ _09820_ _09821_ VGND VGND VPWR VPWR _09822_ sky130_fd_sc_hd__and2_1
X_20375_ _07310_ _07311_ _07259_ _07261_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__o211a_1
Xclkload360 clknet_leaf_12_A_in_serial_clk VGND VGND VPWR VPWR clkload360/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload371 clknet_leaf_2_B_in_serial_clk VGND VGND VPWR VPWR clkload371/Y sky130_fd_sc_hd__bufinv_16
XFILLER_162_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload382 clknet_leaf_25_B_in_serial_clk VGND VGND VPWR VPWR clkload382/Y sky130_fd_sc_hd__clkinv_2
Xclkload393 clknet_leaf_14_B_in_serial_clk VGND VGND VPWR VPWR clkload393/Y sky130_fd_sc_hd__clkinv_2
X_22114_ _08853_ _08862_ _08863_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__nand3_1
XFILLER_122_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload90 clknet_leaf_316_clk VGND VGND VPWR VPWR clkload90/Y sky130_fd_sc_hd__bufinv_16
X_27971_ clknet_leaf_175_clk _01769_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_23094_ _09756_ _09757_ _09755_ VGND VGND VPWR VPWR _09763_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_168_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22045_ _08816_ _08817_ _08818_ VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__or3_1
XFILLER_47_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26922_ clknet_leaf_4_A_in_serial_clk _00720_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26853_ clknet_leaf_70_clk _00655_ net135 VGND VGND VPWR VPWR B_in\[125\] sky130_fd_sc_hd__dfrtp_1
X_29641_ clknet_leaf_30_B_in_serial_clk _03436_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25804_ systolic_inst.acc_wires\[8\]\[24\] C_out\[280\] net28 VGND VGND VPWR VPWR
+ _03106_ sky130_fd_sc_hd__mux2_1
X_29572_ clknet_leaf_21_B_in_serial_clk _03367_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26784_ clknet_leaf_61_clk _00586_ net143 VGND VGND VPWR VPWR B_in\[56\] sky130_fd_sc_hd__dfrtp_1
X_23996_ _10523_ systolic_inst.B_shift\[5\]\[1\] _11332_ VGND VGND VPWR VPWR _02019_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28523_ clknet_leaf_154_clk _02321_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25735_ systolic_inst.acc_wires\[6\]\[19\] C_out\[211\] net46 VGND VGND VPWR VPWR
+ _03037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22947_ systolic_inst.B_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\] VGND VGND VPWR
+ VPWR _09625_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_206_Right_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28454_ clknet_leaf_127_clk _02252_ net144 VGND VGND VPWR VPWR ser_C.shift_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13680_ deser_B.word_buffer\[116\] deser_B.serial_word\[116\] net124 VGND VGND VPWR
+ VPWR _00517_ sky130_fd_sc_hd__mux2_1
X_25666_ systolic_inst.acc_wires\[4\]\[14\] C_out\[142\] net30 VGND VGND VPWR VPWR
+ _02968_ sky130_fd_sc_hd__mux2_1
X_22878_ systolic_inst.B_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[5\] systolic_inst.A_outs\[1\]\[6\]
+ systolic_inst.B_outs\[1\]\[3\] VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__a22oi_1
XFILLER_232_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27405_ clknet_leaf_229_clk _01203_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_54_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24617_ C_out\[135\] net103 net75 ser_C.shift_reg\[135\] _10778_ VGND VGND VPWR VPWR
+ _02385_ sky130_fd_sc_hd__a221o_1
X_21829_ _08631_ _08632_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__nor2_1
XFILLER_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28385_ clknet_leaf_32_clk _02183_ VGND VGND VPWR VPWR systolic_inst.A_shift\[18\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25597_ systolic_inst.acc_wires\[2\]\[9\] C_out\[73\] net34 VGND VGND VPWR VPWR _02899_
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27336_ clknet_leaf_285_clk _01134_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_15350_ _12429_ _12432_ VGND VGND VPWR VPWR _12434_ sky130_fd_sc_hd__or2_1
XFILLER_12_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24548_ net113 ser_C.shift_reg\[102\] VGND VGND VPWR VPWR _10744_ sky130_fd_sc_hd__and2_1
XFILLER_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14301_ systolic_inst.A_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[5\] VGND VGND
+ VPWR VPWR _11487_ sky130_fd_sc_hd__nand2_1
Xwire111 net112 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_12
XFILLER_106_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15281_ _12373_ _12374_ VGND VGND VPWR VPWR _12375_ sky130_fd_sc_hd__and2_1
X_27267_ clknet_leaf_268_clk _01065_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_24479_ C_out\[66\] _11302_ net81 ser_C.shift_reg\[66\] _10709_ VGND VGND VPWR VPWR
+ _02316_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_199_Left_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29006_ clknet_leaf_104_clk _02804_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17020_ _04321_ _04322_ _04320_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__a21bo_1
X_26218_ clknet_leaf_9_A_in_serial_clk _00026_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14232_ _11413_ _11414_ _11418_ VGND VGND VPWR VPWR _11420_ sky130_fd_sc_hd__a21o_1
XFILLER_32_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27198_ clknet_leaf_262_clk _00996_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_165_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_242_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_242_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26149_ deser_B.serial_word\[104\] deser_B.shift_reg\[104\] _00001_ VGND VGND VPWR
+ VPWR _03451_ sky130_fd_sc_hd__mux2_1
X_14163_ _11341_ _11353_ VGND VGND VPWR VPWR _11354_ sky130_fd_sc_hd__nand2_1
XFILLER_109_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_242_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13114_ systolic_inst.A_outs\[0\]\[7\] VGND VGND VPWR VPWR _11270_ sky130_fd_sc_hd__inv_2
XFILLER_113_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14094_ deser_A.receiving net2 net1 VGND VGND VPWR VPWR _11330_ sky130_fd_sc_hd__and3b_1
X_18971_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[25\]
+ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__xor2_2
XFILLER_3_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xload_slew105 net106 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_16
XFILLER_106_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _05110_ _05114_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__and2_1
XFILLER_152_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17853_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[4\] _05049_
+ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__a21bo_1
XFILLER_26_1169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16804_ _04121_ _04123_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__nand2_1
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14996_ _12112_ _12115_ VGND VGND VPWR VPWR _12116_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17784_ _05001_ _05000_ systolic_inst.acc_wires\[10\]\[31\] net105 VGND VGND VPWR
+ VPWR _01329_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_219_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19523_ net105 systolic_inst.acc_wires\[7\]\[17\] net62 _06562_ VGND VGND VPWR VPWR
+ _01507_ sky130_fd_sc_hd__a22o_1
XFILLER_235_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13947_ deser_A.serial_word\[108\] deser_A.shift_reg\[108\] net57 VGND VGND VPWR
+ VPWR _00773_ sky130_fd_sc_hd__mux2_1
X_16735_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[7\]
+ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__o21a_1
XFILLER_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19454_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[7\]\[8\]
+ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16666_ systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[5\] systolic_inst.A_outs\[11\]\[6\]
+ systolic_inst.B_outs\[11\]\[0\] VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__a22oi_1
XFILLER_35_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13878_ deser_A.serial_word\[39\] deser_A.shift_reg\[39\] net58 VGND VGND VPWR VPWR
+ _00704_ sky130_fd_sc_hd__mux2_1
XFILLER_179_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15617_ _12670_ _12671_ VGND VGND VPWR VPWR _12673_ sky130_fd_sc_hd__nand2_1
XFILLER_62_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18405_ systolic_inst.A_outs\[8\]\[2\] systolic_inst.A_shift\[16\]\[2\] net121 VGND
+ VGND VPWR VPWR _01396_ sky130_fd_sc_hd__mux2_1
XFILLER_201_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19385_ _06442_ _06443_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__nor2_1
XFILLER_50_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16597_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _03924_ sky130_fd_sc_hd__and2_1
XFILLER_188_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18336_ _05490_ _05497_ _05498_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__a21oi_1
X_15548_ _12603_ _12604_ VGND VGND VPWR VPWR _12606_ sky130_fd_sc_hd__xor2_1
XFILLER_72_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18267_ _05425_ _05439_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__nand2_1
X_15479_ _12485_ _12513_ _12512_ VGND VGND VPWR VPWR _12538_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17218_ _04477_ _04478_ _04466_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__a21oi_1
X_18198_ _05381_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__inv_2
X_17149_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[27\]
+ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_203_Left_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20160_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[22\]
+ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__nand2_1
XFILLER_116_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20091_ _07055_ _07071_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__nor2_1
XFILLER_131_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23850_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[24\]
+ VGND VGND VPWR VPWR _10443_ sky130_fd_sc_hd__nor2_1
XFILLER_226_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22801_ _09481_ _09482_ VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__and2b_1
XFILLER_242_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23781_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[0\]\[12\]
+ _10381_ VGND VGND VPWR VPWR _10385_ sky130_fd_sc_hd__and3_1
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20993_ _07835_ _07865_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25520_ _11241_ _11242_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_212_Left_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22732_ _09413_ _09415_ _09407_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__a21oi_1
XFILLER_225_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25451_ _11196_ _11197_ systolic_inst.cycle_cnt\[6\] VGND VGND VPWR VPWR _02800_
+ sky130_fd_sc_hd__mux2_1
XFILLER_197_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22663_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[30\]
+ VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__nand2_1
XFILLER_129_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24402_ net114 ser_C.shift_reg\[29\] VGND VGND VPWR VPWR _10671_ sky130_fd_sc_hd__and2_1
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28170_ clknet_leaf_81_clk _01968_ VGND VGND VPWR VPWR systolic_inst.B_shift\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21614_ _08417_ _08423_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__nor2_1
XFILLER_40_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25382_ _11160_ systolic_inst.B_shift\[14\]\[6\] net71 VGND VGND VPWR VPWR _02768_
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22594_ net109 systolic_inst.acc_wires\[2\]\[18\] net65 _09312_ VGND VGND VPWR VPWR
+ _01828_ sky130_fd_sc_hd__a22o_1
XFILLER_194_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27121_ clknet_leaf_0_B_in_serial_clk _00919_ net134 VGND VGND VPWR VPWR deser_B.shift_reg\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_24333_ systolic_inst.A_shift\[10\]\[6\] A_in\[38\] net59 VGND VGND VPWR VPWR _10640_
+ sky130_fd_sc_hd__mux2_1
X_21545_ systolic_inst.A_outs\[3\]\[2\] systolic_inst.B_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\]
+ systolic_inst.A_outs\[3\]\[1\] VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__a22o_1
XFILLER_139_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_141_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_142_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27052_ clknet_leaf_24_B_in_serial_clk _00850_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24264_ systolic_inst.A_shift\[16\]\[7\] net70 net83 systolic_inst.A_shift\[17\]\[7\]
+ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__a22o_1
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21476_ systolic_inst.B_outs\[2\]\[4\] systolic_inst.B_shift\[2\]\[4\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26003_ systolic_inst.acc_wires\[14\]\[31\] ser_C.parallel_data\[479\] net24 VGND
+ VGND VPWR VPWR _03305_ sky130_fd_sc_hd__mux2_1
XFILLER_14_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23215_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[22\]
+ VGND VGND VPWR VPWR _09866_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_221_Left_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20427_ _07361_ _07362_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__or2_1
XFILLER_88_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24195_ systolic_inst.B_shift\[22\]\[2\] net71 _11333_ B_in\[114\] VGND VGND VPWR
+ VPWR _02156_ sky130_fd_sc_hd__a22o_1
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23146_ _09790_ _09806_ VGND VGND VPWR VPWR _09807_ sky130_fd_sc_hd__nor2_1
XFILLER_162_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload190 clknet_leaf_59_clk VGND VGND VPWR VPWR clkload190/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_112_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20358_ systolic_inst.A_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[5\] VGND VGND VPWR
+ VPWR _07296_ sky130_fd_sc_hd__nand2_1
XFILLER_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23077_ net64 _09747_ _09748_ systolic_inst.acc_wires\[1\]\[1\] _11258_ VGND VGND
+ VPWR VPWR _01875_ sky130_fd_sc_hd__a32o_1
X_27954_ clknet_leaf_171_clk _01752_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_20289_ systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[5\]
+ systolic_inst.B_outs\[5\]\[0\] VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22028_ _08786_ _08803_ _08804_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26905_ clknet_leaf_17_A_in_serial_clk _00703_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27885_ clknet_leaf_310_clk _01683_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29624_ clknet_leaf_8_B_in_serial_clk _03419_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_14850_ systolic_inst.A_outs\[14\]\[1\] systolic_inst.B_outs\[14\]\[5\] systolic_inst.B_outs\[14\]\[6\]
+ systolic_inst.A_outs\[14\]\[0\] VGND VGND VPWR VPWR _11974_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_86_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26836_ clknet_leaf_88_clk _00638_ net153 VGND VGND VPWR VPWR B_in\[108\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13801_ B_in\[108\] deser_B.word_buffer\[108\] net88 VGND VGND VPWR VPWR _00638_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_230_Left_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26767_ clknet_leaf_95_clk _00569_ net5 VGND VGND VPWR VPWR B_in\[39\] sky130_fd_sc_hd__dfrtp_1
X_29555_ clknet_leaf_18_B_in_serial_clk _03350_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14781_ _11901_ _11907_ VGND VGND VPWR VPWR _11908_ sky130_fd_sc_hd__or2_1
XFILLER_95_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23979_ systolic_inst.B_shift\[12\]\[1\] B_in\[65\] _00008_ VGND VGND VPWR VPWR _10515_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16520_ _03873_ _03874_ _03872_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__o21ai_1
X_28506_ clknet_leaf_110_clk _02304_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_217_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13732_ B_in\[39\] deser_B.word_buffer\[39\] net90 VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__mux2_1
X_25718_ systolic_inst.acc_wires\[6\]\[2\] C_out\[194\] net47 VGND VGND VPWR VPWR
+ _03020_ sky130_fd_sc_hd__mux2_1
XFILLER_44_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_231_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26698_ clknet_leaf_5_B_in_serial_clk _00501_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_29486_ clknet_leaf_281_clk _03284_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[458\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_231_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16451_ _03811_ _03815_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__or2_1
X_25649_ systolic_inst.acc_wires\[3\]\[29\] C_out\[125\] net49 VGND VGND VPWR VPWR
+ _02951_ sky130_fd_sc_hd__mux2_1
X_13663_ deser_B.word_buffer\[99\] deser_B.serial_word\[99\] net123 VGND VGND VPWR
+ VPWR _00500_ sky130_fd_sc_hd__mux2_1
XFILLER_147_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28437_ clknet_leaf_25_clk _02235_ VGND VGND VPWR VPWR systolic_inst.A_shift\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15402_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.A_outs\[13\]\[1\] systolic_inst.B_outs\[13\]\[3\]
+ systolic_inst.B_outs\[13\]\[4\] VGND VGND VPWR VPWR _12464_ sky130_fd_sc_hd__nand4_1
XFILLER_227_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19170_ systolic_inst.B_outs\[7\]\[7\] _06201_ _06202_ VGND VGND VPWR VPWR _06235_
+ sky130_fd_sc_hd__a21bo_1
X_16382_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[12\]\[3\]
+ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__nand2_1
X_28368_ clknet_leaf_5_clk _02166_ VGND VGND VPWR VPWR systolic_inst.A_shift\[20\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13594_ deser_B.word_buffer\[30\] deser_B.serial_word\[30\] net124 VGND VGND VPWR
+ VPWR _00431_ sky130_fd_sc_hd__mux2_1
XFILLER_160_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18121_ _05257_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__and2b_1
XFILLER_169_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27319_ clknet_leaf_289_clk _01117_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15333_ _12403_ _12405_ _12417_ _12418_ _12411_ VGND VGND VPWR VPWR _12419_ sky130_fd_sc_hd__a311oi_4
XFILLER_8_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28299_ clknet_leaf_123_clk _02097_ VGND VGND VPWR VPWR systolic_inst.B_shift\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_132_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_26_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18052_ _05242_ _05241_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_229_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15264_ _12360_ VGND VGND VPWR VPWR _12361_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_229_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17003_ _04308_ _04309_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__a21o_1
X_14215_ _11360_ _11384_ _11383_ VGND VGND VPWR VPWR _11403_ sky130_fd_sc_hd__a21bo_1
XANTENNA_5 _11176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15195_ _11712_ _12300_ _12301_ systolic_inst.acc_wires\[14\]\[7\] net107 VGND VGND
+ VPWR VPWR _01049_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_39_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14146_ net107 systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _11338_ sky130_fd_sc_hd__and2_1
XFILLER_141_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14077_ deser_B.shift_reg\[111\] deser_B.shift_reg\[112\] deser_B.receiving VGND
+ VGND VPWR VPWR _00903_ sky130_fd_sc_hd__mux2_1
XFILLER_140_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18954_ _06049_ _06050_ _06051_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__or3_1
XFILLER_234_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17905_ _05068_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_199_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_199_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18885_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[8\]\[13\]
+ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__or2_1
XFILLER_121_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17836_ _05029_ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_176_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17767_ net105 systolic_inst.acc_wires\[10\]\[28\] net62 _04987_ VGND VGND VPWR VPWR
+ _01326_ sky130_fd_sc_hd__a22o_1
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14979_ _12099_ VGND VGND VPWR VPWR _12100_ sky130_fd_sc_hd__inv_2
XFILLER_130_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19506_ _06540_ _06544_ _06546_ _06547_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__a211o_1
X_16718_ _04003_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__or2_1
X_17698_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[18\]
+ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__nand2_1
XFILLER_39_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19437_ _06479_ _06483_ _06486_ _06487_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__o211a_1
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16649_ _03970_ _03972_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[3\]
+ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__and4b_1
XFILLER_23_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19368_ _06396_ _06401_ _06427_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_214_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18319_ net66 _05484_ _05485_ systolic_inst.acc_wires\[9\]\[18\] net106 VGND VGND
+ VPWR VPWR _01380_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_123_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19299_ _06359_ _06360_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__nand2_1
XFILLER_241_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21330_ _08160_ _08164_ _08165_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__o21ai_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21261_ net63 _08123_ _08124_ systolic_inst.acc_wires\[4\]\[1\] net108 VGND VGND
+ VPWR VPWR _01683_ sky130_fd_sc_hd__a32o_1
XFILLER_198_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23000_ _09586_ _09645_ _09643_ VGND VGND VPWR VPWR _09677_ sky130_fd_sc_hd__a21oi_1
X_20212_ _07165_ _07168_ _07171_ _07174_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_165_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21192_ systolic_inst.A_outs\[4\]\[6\] _11271_ _07850_ VGND VGND VPWR VPWR _08060_
+ sky130_fd_sc_hd__o21a_1
XFILLER_171_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_165_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20143_ _07115_ _07116_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20074_ net60 _07057_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__nor2_1
X_24951_ C_out\[302\] net103 net76 ser_C.shift_reg\[302\] _10945_ VGND VGND VPWR VPWR
+ _02552_ sky130_fd_sc_hd__a221o_1
XFILLER_213_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23902_ systolic_inst.B_shift\[17\]\[3\] B_in\[75\] _00008_ VGND VGND VPWR VPWR _10484_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27670_ clknet_leaf_146_clk _01468_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24882_ net110 ser_C.shift_reg\[269\] VGND VGND VPWR VPWR _10911_ sky130_fd_sc_hd__and2_1
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26621_ clknet_leaf_22_B_in_serial_clk _00424_ net137 VGND VGND VPWR VPWR deser_B.word_buffer\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23833_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[22\]
+ VGND VGND VPWR VPWR _10428_ sky130_fd_sc_hd__or2_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29340_ clknet_leaf_214_clk _03138_ net149 VGND VGND VPWR VPWR C_out\[312\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26552_ clknet_leaf_26_A_in_serial_clk _00355_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_23764_ _10368_ _10369_ VGND VGND VPWR VPWR _10370_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_159_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20976_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[7\] VGND VGND VPWR
+ VPWR _07850_ sky130_fd_sc_hd__nand2_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25503_ systolic_inst.cycle_cnt\[24\] _11279_ _11228_ systolic_inst.cycle_cnt\[23\]
+ VGND VGND VPWR VPWR _11232_ sky130_fd_sc_hd__a22oi_1
XFILLER_241_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22715_ _09386_ _09388_ _09399_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__a21oi_2
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29271_ clknet_leaf_193_clk _03069_ net146 VGND VGND VPWR VPWR C_out\[243\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26483_ clknet_leaf_12_A_in_serial_clk _00286_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23695_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[0\]\[1\]
+ VGND VGND VPWR VPWR _10311_ sky130_fd_sc_hd__nand2_1
XFILLER_53_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28222_ clknet_leaf_103_clk _02020_ VGND VGND VPWR VPWR systolic_inst.B_shift\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25434_ systolic_inst.cycle_cnt\[1\] systolic_inst.cycle_cnt\[0\] VGND VGND VPWR
+ VPWR _11186_ sky130_fd_sc_hd__nand2_1
XFILLER_224_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22646_ _09354_ _09355_ VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28153_ clknet_leaf_102_clk _01951_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_25365_ ser_C.parallel_data\[509\] net98 net78 ser_C.shift_reg\[509\] _11152_ VGND
+ VGND VPWR VPWR _02759_ sky130_fd_sc_hd__a221o_1
X_22577_ _09296_ _09297_ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_114_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27104_ clknet_leaf_10_B_in_serial_clk _00902_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24316_ _10631_ systolic_inst.A_shift\[10\]\[5\] net71 VGND VGND VPWR VPWR _02231_
+ sky130_fd_sc_hd__mux2_1
X_28084_ clknet_leaf_116_clk _01882_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_21528_ _08338_ _08340_ _08322_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25296_ net111 ser_C.shift_reg\[476\] VGND VGND VPWR VPWR _11118_ sky130_fd_sc_hd__and2_1
XFILLER_215_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27035_ clknet_leaf_13_B_in_serial_clk _00833_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_193_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24247_ systolic_inst.A_shift\[19\]\[7\] A_in\[71\] net59 VGND VGND VPWR VPWR _10609_
+ sky130_fd_sc_hd__mux2_1
X_21459_ net63 _08292_ _08293_ systolic_inst.acc_wires\[4\]\[30\] _11258_ VGND VGND
+ VPWR VPWR _01712_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_A_in_serial_clk clknet_2_2__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_3_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_218_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14000_ deser_B.shift_reg\[34\] deser_B.shift_reg\[35\] deser_B.receiving VGND VGND
+ VPWR VPWR _00826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_224_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput7 net110 VGND VGND VPWR VPWR C_out_frame_sync sky130_fd_sc_hd__buf_1
X_24178_ systolic_inst.A_shift\[25\]\[1\] net70 _10505_ systolic_inst.A_shift\[26\]\[1\]
+ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__a22o_1
XFILLER_150_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23129_ _11713_ _09792_ VGND VGND VPWR VPWR _09793_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_220_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28986_ clknet_leaf_25_clk _02784_ VGND VGND VPWR VPWR systolic_inst.A_shift\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_31_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_95_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27937_ clknet_leaf_171_clk _01735_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_153_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15951_ _12969_ _12970_ VGND VGND VPWR VPWR _12971_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14902_ _11985_ _11988_ _12024_ VGND VGND VPWR VPWR _12025_ sky130_fd_sc_hd__o21ai_1
X_15882_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[20\]
+ VGND VGND VPWR VPWR _12912_ sky130_fd_sc_hd__or2_1
XFILLER_7_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18670_ _05795_ _05796_ _05794_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__a21oi_2
X_27868_ clknet_leaf_317_clk _01666_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29607_ clknet_leaf_24_B_in_serial_clk _03402_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17621_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[10\]\[7\]
+ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__or2_1
XFILLER_236_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26819_ clknet_leaf_67_clk _00621_ net135 VGND VGND VPWR VPWR B_in\[91\] sky130_fd_sc_hd__dfrtp_1
X_14833_ _11928_ _11931_ VGND VGND VPWR VPWR _11958_ sky130_fd_sc_hd__nor2_1
X_27799_ clknet_leaf_45_clk _01597_ net137 VGND VGND VPWR VPWR systolic_inst.B_outs\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_218_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.A_outs\[14\]\[2\] VGND VGND
+ VPWR VPWR _11892_ sky130_fd_sc_hd__nand2_1
X_29538_ clknet_leaf_246_clk _03336_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[510\]
+ sky130_fd_sc_hd__dfrtp_1
X_17552_ _04776_ _04779_ _04801_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__and3_1
XFILLER_229_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13715_ B_in\[22\] deser_B.word_buffer\[22\] net86 VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16503_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[20\]
+ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__xor2_1
X_17483_ _04701_ _04705_ _04733_ _04735_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__o22a_1
XFILLER_189_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29469_ clknet_leaf_286_clk _03267_ net136 VGND VGND VPWR VPWR ser_C.parallel_data\[441\]
+ sky130_fd_sc_hd__dfrtp_1
X_14695_ _11843_ _11845_ _11848_ VGND VGND VPWR VPWR _11849_ sky130_fd_sc_hd__and3_1
XFILLER_72_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19222_ _06282_ _06285_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13646_ deser_B.word_buffer\[82\] deser_B.serial_word\[82\] net124 VGND VGND VPWR
+ VPWR _00483_ sky130_fd_sc_hd__mux2_1
X_16434_ net67 _03799_ _03800_ systolic_inst.acc_wires\[12\]\[10\] net108 VGND VGND
+ VPWR VPWR _01180_ sky130_fd_sc_hd__a32o_1
XFILLER_60_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19153_ _06212_ _06218_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16365_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[12\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_105_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13577_ deser_B.word_buffer\[13\] deser_B.serial_word\[13\] net124 VGND VGND VPWR
+ VPWR _00414_ sky130_fd_sc_hd__mux2_1
XFILLER_34_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15316_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[25\]
+ VGND VGND VPWR VPWR _12405_ sky130_fd_sc_hd__xor2_2
X_18104_ systolic_inst.B_outs\[9\]\[6\] systolic_inst.A_outs\[9\]\[6\] _11263_ systolic_inst.A_outs\[9\]\[5\]
+ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_17__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_17__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_19084_ systolic_inst.A_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\]
+ systolic_inst.A_outs\[7\]\[1\] VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__a22oi_1
XFILLER_118_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16296_ _03674_ _03675_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15247_ net67 _12345_ _12346_ systolic_inst.acc_wires\[14\]\[14\] net107 VGND VGND
+ VPWR VPWR _01056_ sky130_fd_sc_hd__a32o_1
X_18035_ _05191_ _05225_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__xor2_1
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15178_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[14\]\[5\]
+ VGND VGND VPWR VPWR _12287_ sky130_fd_sc_hd__nand2_1
XFILLER_153_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_136_Left_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14129_ systolic_inst.A_outs\[15\]\[5\] systolic_inst.A_outs\[14\]\[5\] net118 VGND
+ VGND VPWR VPWR _00951_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19986_ _06895_ _06980_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__or2_1
XFILLER_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_207_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18937_ _06017_ _06022_ _06027_ _06032_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__or4_1
XFILLER_140_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18868_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[8\]\[11\]
+ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__nand2_1
XFILLER_223_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17819_ _05015_ _05016_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__or2_1
X_18799_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[8\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__a21o_1
XFILLER_242_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20830_ systolic_inst.A_outs\[4\]\[3\] systolic_inst.A_shift\[8\]\[3\] net121 VGND
+ VGND VPWR VPWR _01653_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_145_Left_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20761_ _07660_ _07666_ _07667_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_344_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_344_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22500_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[2\]\[5\]
+ VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_154_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23480_ _11258_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[8\] _10104_
+ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_154_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20692_ _07608_ _07609_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__nand2_1
XFILLER_50_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22431_ _09168_ _09169_ VGND VGND VPWR VPWR _09171_ sky130_fd_sc_hd__and2b_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25150_ net110 ser_C.shift_reg\[403\] VGND VGND VPWR VPWR _11045_ sky130_fd_sc_hd__and2_1
X_22362_ _09101_ _09102_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24101_ systolic_inst.B_shift\[23\]\[6\] B_in\[62\] _00008_ VGND VGND VPWR VPWR _10560_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21313_ _08160_ _08163_ _08166_ VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__a21bo_1
X_25081_ C_out\[367\] net97 net77 ser_C.shift_reg\[367\] _11010_ VGND VGND VPWR VPWR
+ _02617_ sky130_fd_sc_hd__a221o_1
X_22293_ _09034_ _09035_ VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_154_Left_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24032_ _10533_ systolic_inst.B_shift\[4\]\[3\] net72 VGND VGND VPWR VPWR _02045_
+ sky130_fd_sc_hd__mux2_1
X_21244_ net117 _08109_ _08110_ _08088_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__a31o_1
XFILLER_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_1155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28840_ clknet_leaf_328_clk _02638_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[388\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21175_ _08042_ _08043_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__nand2_1
XFILLER_120_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20126_ _07100_ _07101_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__nor2_1
XFILLER_137_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25983_ systolic_inst.acc_wires\[14\]\[11\] ser_C.parallel_data\[459\] net26 VGND
+ VGND VPWR VPWR _03285_ sky130_fd_sc_hd__mux2_1
XFILLER_104_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28771_ clknet_leaf_225_clk _02569_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[319\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_219_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27722_ clknet_leaf_190_clk _01520_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_20057_ net68 _07041_ _07043_ systolic_inst.acc_wires\[6\]\[6\] net106 VGND VGND
+ VPWR VPWR _01560_ sky130_fd_sc_hd__a32o_1
X_24934_ net111 ser_C.shift_reg\[295\] VGND VGND VPWR VPWR _10937_ sky130_fd_sc_hd__and2_1
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24865_ C_out\[259\] net101 net73 ser_C.shift_reg\[259\] _10902_ VGND VGND VPWR VPWR
+ _02509_ sky130_fd_sc_hd__a221o_1
X_27653_ clknet_leaf_313_clk _01451_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_93_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23816_ _10412_ _10414_ VGND VGND VPWR VPWR _10415_ sky130_fd_sc_hd__xor2_1
X_26604_ clknet_leaf_16_B_in_serial_clk _00407_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_27584_ clknet_leaf_216_clk _01382_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24796_ net112 ser_C.shift_reg\[226\] VGND VGND VPWR VPWR _10868_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29323_ clknet_leaf_304_clk _03121_ net138 VGND VGND VPWR VPWR C_out\[295\] sky130_fd_sc_hd__dfrtp_1
X_26535_ clknet_leaf_16_A_in_serial_clk _00338_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_23747_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[0\]\[9\]
+ VGND VGND VPWR VPWR _10355_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_335_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_335_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_53_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20959_ net108 systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[6\] _07833_
+ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__a21bo_1
XFILLER_199_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13500_ deser_A.shift_reg\[64\] deser_A.shift_reg\[65\] net129 VGND VGND VPWR VPWR
+ _00337_ sky130_fd_sc_hd__mux2_1
XFILLER_159_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29254_ clknet_leaf_197_clk _03052_ net147 VGND VGND VPWR VPWR C_out\[226\] sky130_fd_sc_hd__dfrtp_1
X_14480_ _11659_ _11660_ VGND VGND VPWR VPWR _11661_ sky130_fd_sc_hd__nand2_1
X_26466_ clknet_leaf_1_A_in_serial_clk _00273_ net132 VGND VGND VPWR VPWR deser_A.bit_idx\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_23678_ _10295_ _10296_ VGND VGND VPWR VPWR _10297_ sky130_fd_sc_hd__nand2_1
XFILLER_241_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_B_in_serial_clk clknet_2_2__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_10_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28205_ clknet_leaf_94_clk _02003_ VGND VGND VPWR VPWR systolic_inst.B_shift\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25417_ systolic_inst.A_shift\[1\]\[0\] A_in\[0\] net59 VGND VGND VPWR VPWR _11178_
+ sky130_fd_sc_hd__mux2_1
X_13431_ deser_A.bit_idx\[3\] deser_A.bit_idx\[4\] _11312_ VGND VGND VPWR VPWR _11316_
+ sky130_fd_sc_hd__and3_1
X_22629_ _09340_ _09341_ VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__or2_1
X_29185_ clknet_leaf_135_clk _02983_ net142 VGND VGND VPWR VPWR C_out\[157\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26397_ clknet_leaf_27_clk _00204_ net137 VGND VGND VPWR VPWR A_in\[65\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28136_ clknet_leaf_126_clk _01934_ net144 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16150_ _03526_ _03534_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__nand2_1
XFILLER_107_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25348_ net112 ser_C.shift_reg\[502\] VGND VGND VPWR VPWR _11144_ sky130_fd_sc_hd__and2_1
XFILLER_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13362_ A_in\[71\] deser_A.word_buffer\[71\] net94 VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__mux2_1
X_15101_ _12216_ _12217_ VGND VGND VPWR VPWR _12218_ sky130_fd_sc_hd__nand2b_1
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28067_ clknet_leaf_120_clk _01865_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16081_ _13031_ _13033_ _13076_ VGND VGND VPWR VPWR _13077_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13293_ A_in\[2\] deser_A.word_buffer\[2\] net93 VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__mux2_1
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25279_ ser_C.parallel_data\[466\] net102 net74 ser_C.shift_reg\[466\] _11109_ VGND
+ VGND VPWR VPWR _02716_ sky130_fd_sc_hd__a221o_1
XFILLER_182_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27018_ clknet_leaf_22_B_in_serial_clk _00816_ net137 VGND VGND VPWR VPWR deser_B.shift_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_15032_ _12147_ _12150_ VGND VGND VPWR VPWR _12151_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19840_ _06799_ _06801_ _06838_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__nand3_1
XFILLER_29_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19771_ _06742_ _06771_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28969_ clknet_leaf_53_clk _02767_ VGND VGND VPWR VPWR systolic_inst.B_shift\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16983_ _04290_ _04291_ _04292_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_53_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18722_ _05845_ _05846_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__nand2_1
X_15934_ _12949_ _12953_ VGND VGND VPWR VPWR _12956_ sky130_fd_sc_hd__nor2_1
XFILLER_49_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_202_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18653_ _05770_ _05778_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__or2_1
X_15865_ net108 systolic_inst.acc_wires\[13\]\[16\] _12896_ _12898_ VGND VGND VPWR
+ VPWR _01122_ sky130_fd_sc_hd__a22o_1
XFILLER_236_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17604_ _04844_ _04845_ _04846_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__a21o_1
X_14816_ _11920_ _11939_ VGND VGND VPWR VPWR _11941_ sky130_fd_sc_hd__xnor2_1
X_18584_ _05704_ _05712_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_194_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[13\]\[7\]
+ VGND VGND VPWR VPWR _12839_ sky130_fd_sc_hd__or2_1
XFILLER_40_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_194_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _04786_ _04785_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__and2b_1
XFILLER_45_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_326_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_326_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14747_ systolic_inst.A_outs\[14\]\[7\] systolic_inst.A_outs\[13\]\[7\] net116 VGND
+ VGND VPWR VPWR _01017_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_190_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_190_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14678_ systolic_inst.acc_wires\[15\]\[20\] systolic_inst.acc_wires\[15\]\[21\] systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _11834_ sky130_fd_sc_hd__o21a_1
X_17466_ _04679_ _04681_ _04680_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__o21ba_1
XFILLER_220_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19205_ _06231_ _06232_ _06230_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__a21o_1
X_13629_ deser_B.word_buffer\[65\] deser_B.serial_word\[65\] net123 VGND VGND VPWR
+ VPWR _00466_ sky130_fd_sc_hd__mux2_1
X_16417_ _03784_ _03785_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__and2_1
XFILLER_38_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17397_ _04612_ _04614_ _04613_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__o21ba_1
XFILLER_186_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19136_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[6\]
+ systolic_inst.A_outs\[7\]\[7\] VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__nand4_1
XFILLER_203_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16348_ _03725_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__nor2_1
XFILLER_34_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19067_ _06115_ _06133_ _06134_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__or3_1
XFILLER_12_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16279_ _03658_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__nand2_2
XFILLER_161_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_209_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18018_ _05209_ _05208_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19969_ _06962_ _06963_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__xor2_1
XFILLER_99_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22980_ systolic_inst.B_outs\[1\]\[6\] systolic_inst.A_outs\[1\]\[6\] _11277_ systolic_inst.A_outs\[1\]\[5\]
+ VGND VGND VPWR VPWR _09657_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_143_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21931_ _08711_ _08715_ _08721_ VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__a21o_1
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24650_ net7 ser_C.shift_reg\[153\] VGND VGND VPWR VPWR _10795_ sky130_fd_sc_hd__and2_1
XFILLER_242_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21862_ _08583_ _08643_ VGND VGND VPWR VPWR _08664_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23601_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[7\]
+ VGND VGND VPWR VPWR _10222_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20813_ _07710_ _07712_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__xnor2_1
X_24581_ C_out\[117\] net100 net82 ser_C.shift_reg\[117\] _10760_ VGND VGND VPWR VPWR
+ _02367_ sky130_fd_sc_hd__a221o_1
X_21793_ _08563_ _08565_ _08596_ VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_317_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_317_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_151_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26320_ clknet_leaf_0_A_in_serial_clk _00128_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_196_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23532_ systolic_inst.A_outs\[0\]\[6\] _10154_ _10153_ VGND VGND VPWR VPWR _10155_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_180_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20744_ _07652_ _07654_ VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__xor2_1
XFILLER_24_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26251_ clknet_leaf_9_A_in_serial_clk _00059_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23463_ _10086_ _10087_ VGND VGND VPWR VPWR _10088_ sky130_fd_sc_hd__nand2_1
XFILLER_221_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20675_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[5\]\[9\]
+ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__xor2_1
XFILLER_52_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25202_ net110 ser_C.shift_reg\[429\] VGND VGND VPWR VPWR _11071_ sky130_fd_sc_hd__and2_1
X_22414_ systolic_inst.B_outs\[2\]\[6\] systolic_inst.A_outs\[2\]\[7\] VGND VGND VPWR
+ VPWR _09154_ sky130_fd_sc_hd__nand2_1
XFILLER_177_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26182_ ser_C.bit_idx\[3\] ser_C.bit_idx\[4\] _11247_ VGND VGND VPWR VPWR _11250_
+ sky130_fd_sc_hd__and3_1
XFILLER_183_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23394_ _09986_ _09988_ _10020_ VGND VGND VPWR VPWR _10021_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_162_Left_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25133_ C_out\[393\] net101 net73 ser_C.shift_reg\[393\] _11036_ VGND VGND VPWR VPWR
+ _02643_ sky130_fd_sc_hd__a221o_1
X_22345_ _09050_ _09051_ _09086_ _09048_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__a211oi_2
XFILLER_87_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25064_ net112 ser_C.shift_reg\[360\] VGND VGND VPWR VPWR _11002_ sky130_fd_sc_hd__and2_1
XFILLER_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22276_ _08982_ _08988_ _08987_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__a21o_1
XFILLER_163_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24015_ systolic_inst.B_shift\[7\]\[6\] _11332_ net83 systolic_inst.B_shift\[11\]\[6\]
+ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__a22o_1
X_21227_ _08092_ _08093_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__nand2_1
XFILLER_176_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28823_ clknet_leaf_239_clk _02621_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[371\]
+ sky130_fd_sc_hd__dfrtp_1
X_21158_ systolic_inst.A_outs\[4\]\[6\] _07884_ _07923_ _07999_ VGND VGND VPWR VPWR
+ _08027_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20109_ _07085_ _07086_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13980_ deser_B.shift_reg\[14\] deser_B.shift_reg\[15\] net125 VGND VGND VPWR VPWR
+ _00806_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28754_ clknet_leaf_220_clk _02552_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[302\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_171_Left_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21089_ systolic_inst.A_outs\[4\]\[5\] systolic_inst.B_outs\[4\]\[5\] systolic_inst.A_outs\[4\]\[7\]
+ systolic_inst.B_outs\[4\]\[1\] VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__a22o_1
X_25966_ systolic_inst.acc_wires\[13\]\[26\] ser_C.parallel_data\[442\] net19 VGND
+ VGND VPWR VPWR _03268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27705_ clknet_leaf_199_clk _01503_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24917_ C_out\[285\] net103 net75 ser_C.shift_reg\[285\] _10928_ VGND VGND VPWR VPWR
+ _02535_ sky130_fd_sc_hd__a221o_1
XFILLER_101_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28685_ clknet_leaf_194_clk _02483_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[233\]
+ sky130_fd_sc_hd__dfrtp_1
X_25897_ systolic_inst.acc_wires\[11\]\[21\] C_out\[373\] net41 VGND VGND VPWR VPWR
+ _03199_ sky130_fd_sc_hd__mux2_1
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _12703_ _12704_ VGND VGND VPWR VPWR _12705_ sky130_fd_sc_hd__nor2_1
X_27636_ clknet_leaf_315_clk _01434_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_215_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24848_ net113 ser_C.shift_reg\[252\] VGND VGND VPWR VPWR _10894_ sky130_fd_sc_hd__and2_1
XFILLER_46_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14601_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[15\]\[11\]
+ VGND VGND VPWR VPWR _11768_ sky130_fd_sc_hd__nand2_1
XFILLER_61_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15581_ _12610_ _12637_ VGND VGND VPWR VPWR _12638_ sky130_fd_sc_hd__nand2b_1
X_24779_ C_out\[216\] net98 net78 ser_C.shift_reg\[216\] _10859_ VGND VGND VPWR VPWR
+ _02466_ sky130_fd_sc_hd__a221o_1
XFILLER_15_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27567_ clknet_leaf_299_clk _01365_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_308_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_308_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14532_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[15\]\[1\]
+ VGND VGND VPWR VPWR _11709_ sky130_fd_sc_hd__or2_1
XFILLER_18_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29306_ clknet_leaf_326_clk _03104_ net141 VGND VGND VPWR VPWR C_out\[278\] sky130_fd_sc_hd__dfrtp_1
X_17320_ systolic_inst.A_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[7\] VGND VGND
+ VPWR VPWR _04578_ sky130_fd_sc_hd__and2b_1
XFILLER_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26518_ clknet_leaf_10_A_in_serial_clk _00321_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_202_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27498_ clknet_leaf_225_clk _01296_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_230_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29237_ clknet_leaf_182_clk _03035_ net148 VGND VGND VPWR VPWR C_out\[209\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14463_ _11643_ _11644_ VGND VGND VPWR VPWR _11645_ sky130_fd_sc_hd__nor2_1
X_17251_ _04491_ _04510_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26449_ clknet_leaf_9_clk _00256_ net132 VGND VGND VPWR VPWR A_in\[117\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_180_Left_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16202_ _03547_ _03551_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__o21ai_1
X_13414_ A_in\[123\] deser_A.word_buffer\[123\] _00003_ VGND VGND VPWR VPWR _00262_
+ sky130_fd_sc_hd__mux2_1
X_17182_ systolic_inst.A_outs\[10\]\[4\] systolic_inst.A_outs\[9\]\[4\] net120 VGND
+ VGND VPWR VPWR _01270_ sky130_fd_sc_hd__mux2_1
X_29168_ clknet_leaf_39_clk _02966_ net142 VGND VGND VPWR VPWR C_out\[140\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14394_ _11577_ _11552_ VGND VGND VPWR VPWR _11578_ sky130_fd_sc_hd__nand2b_1
XFILLER_167_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16133_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] _03517_ VGND
+ VGND VPWR VPWR _03518_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_42_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28119_ clknet_leaf_126_clk _01917_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13345_ A_in\[54\] deser_A.word_buffer\[54\] net92 VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__mux2_1
X_29099_ clknet_leaf_154_clk _02897_ net150 VGND VGND VPWR VPWR C_out\[71\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16064_ _13029_ _13059_ VGND VGND VPWR VPWR _13060_ sky130_fd_sc_hd__and2_1
XFILLER_192_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13276_ deser_A.word_buffer\[114\] deser_A.serial_word\[114\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__mux2_1
XFILLER_143_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15015_ _12132_ _12133_ VGND VGND VPWR VPWR _12135_ sky130_fd_sc_hd__xor2_1
XFILLER_68_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_204_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19823_ _06783_ _06821_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_204_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19754_ _06752_ _06755_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16966_ _04276_ _04279_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_200_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18705_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[11\] VGND
+ VGND VPWR VPWR _05831_ sky130_fd_sc_hd__and2_1
X_15917_ _12936_ _12938_ _12941_ net61 VGND VGND VPWR VPWR _12943_ sky130_fd_sc_hd__a31o_1
X_19685_ _06688_ _06685_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_5_B_in_serial_clk clknet_2_2__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_5_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_16897_ _04166_ _04182_ _04180_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_192_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_192_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18636_ _05735_ _05736_ _05737_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_192_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _12876_ _12883_ VGND VGND VPWR VPWR _12884_ sky130_fd_sc_hd__nand2_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18567_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] _05695_ VGND
+ VGND VPWR VPWR _05696_ sky130_fd_sc_hd__a21o_1
X_15779_ _12824_ VGND VGND VPWR VPWR _12825_ sky130_fd_sc_hd__inv_2
XFILLER_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17518_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[12\] _04770_ net118
+ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__mux2_1
XFILLER_75_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18498_ _05627_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__or2_1
XFILLER_221_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17449_ _04665_ _04702_ _04703_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__and3_1
XFILLER_220_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20460_ _07322_ _07393_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__and2_1
XFILLER_146_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19119_ _06156_ _06184_ _06185_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__and3_1
XFILLER_146_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20391_ systolic_inst.B_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[4\]
+ systolic_inst.A_outs\[5\]\[5\] VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__and4_1
XFILLER_238_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22130_ systolic_inst.A_outs\[2\]\[4\] _08878_ VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_149_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22061_ net60 _08833_ net106 systolic_inst.acc_wires\[3\]\[28\] VGND VGND VPWR VPWR
+ _01774_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21012_ systolic_inst.A_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[5\] systolic_inst.A_outs\[4\]\[7\]
+ systolic_inst.B_outs\[4\]\[1\] VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__a22o_1
XFILLER_47_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25820_ systolic_inst.acc_wires\[9\]\[8\] C_out\[296\] net15 VGND VGND VPWR VPWR
+ _03122_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25751_ systolic_inst.acc_wires\[7\]\[3\] C_out\[227\] net40 VGND VGND VPWR VPWR
+ _03053_ sky130_fd_sc_hd__mux2_1
XFILLER_68_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22963_ _09624_ _09640_ VGND VGND VPWR VPWR _09641_ sky130_fd_sc_hd__xor2_1
XFILLER_216_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_94_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21914_ _08706_ _08707_ _08701_ _08704_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__a211o_1
X_24702_ net113 ser_C.shift_reg\[179\] VGND VGND VPWR VPWR _10821_ sky130_fd_sc_hd__and2_1
XFILLER_215_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28470_ clknet_leaf_100_clk _02268_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_25682_ systolic_inst.acc_wires\[4\]\[30\] C_out\[158\] net31 VGND VGND VPWR VPWR
+ _02984_ sky130_fd_sc_hd__mux2_1
X_22894_ _09556_ _09572_ VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24633_ C_out\[143\] net104 _10643_ ser_C.shift_reg\[143\] _10786_ VGND VGND VPWR
+ VPWR _02393_ sky130_fd_sc_hd__a221o_1
X_27421_ clknet_leaf_250_clk _01219_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_21845_ _08646_ _08647_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__nor2_1
XFILLER_93_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24564_ net113 ser_C.shift_reg\[110\] VGND VGND VPWR VPWR _10752_ sky130_fd_sc_hd__and2_1
XFILLER_184_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27352_ clknet_leaf_233_clk _01150_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21776_ net122 _08579_ _08580_ _08581_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__a31o_1
XFILLER_180_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23515_ _10136_ _10137_ _10094_ _10096_ VGND VGND VPWR VPWR _10139_ sky130_fd_sc_hd__a211o_1
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26303_ clknet_leaf_24_A_in_serial_clk _00111_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20727_ _07628_ _07634_ _07635_ VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__o21ba_1
X_27283_ clknet_leaf_320_clk _01081_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_24495_ C_out\[74\] _11302_ net81 ser_C.shift_reg\[74\] _10717_ VGND VGND VPWR VPWR
+ _02324_ sky130_fd_sc_hd__a221o_1
XFILLER_196_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29022_ clknet_leaf_93_clk _02820_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_156_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26234_ clknet_leaf_12_A_in_serial_clk _00042_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23446_ _10064_ _10070_ VGND VGND VPWR VPWR _10071_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_134_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20658_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[5\]\[6\]
+ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__or2_1
XFILLER_11_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26165_ deser_B.serial_word\[120\] deser_B.shift_reg\[120\] net56 VGND VGND VPWR
+ VPWR _03467_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23377_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[4\]
+ systolic_inst.A_outs\[0\]\[5\] VGND VGND VPWR VPWR _10004_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_95_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20589_ net109 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[13\] _07518_
+ _07520_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13130_ deser_B.bit_idx\[3\] deser_B.bit_idx\[5\] deser_B.bit_idx\[4\] _11283_ VGND
+ VGND VPWR VPWR _11284_ sky130_fd_sc_hd__and4_1
XFILLER_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25116_ net110 ser_C.shift_reg\[386\] VGND VGND VPWR VPWR _11028_ sky130_fd_sc_hd__and2_1
X_22328_ _09062_ _09070_ VGND VGND VPWR VPWR _09071_ sky130_fd_sc_hd__nand2_1
XFILLER_125_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26096_ deser_B.serial_word\[51\] deser_B.shift_reg\[51\] net56 VGND VGND VPWR VPWR
+ _03398_ sky130_fd_sc_hd__mux2_1
XFILLER_125_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25047_ C_out\[350\] net98 net78 ser_C.shift_reg\[350\] _10993_ VGND VGND VPWR VPWR
+ _02600_ sky130_fd_sc_hd__a221o_1
X_22259_ _08994_ _09002_ VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_240_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_240_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_240_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28806_ clknet_leaf_246_clk _02604_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[354\]
+ sky130_fd_sc_hd__dfrtp_1
X_16820_ _04135_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26998_ clknet_leaf_16_B_in_serial_clk _00796_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28737_ clknet_leaf_301_clk _02535_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[285\]
+ sky130_fd_sc_hd__dfrtp_1
X_16751_ systolic_inst.A_outs\[11\]\[2\] systolic_inst.B_outs\[11\]\[5\] _04035_ _04034_
+ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__a31o_1
X_25949_ systolic_inst.acc_wires\[13\]\[9\] C_out\[425\] net19 VGND VGND VPWR VPWR
+ _03251_ sky130_fd_sc_hd__mux2_1
X_13963_ deser_A.serial_word\[124\] deser_A.shift_reg\[124\] _00002_ VGND VGND VPWR
+ VPWR _00789_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_85_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_47_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15702_ _12687_ _12753_ VGND VGND VPWR VPWR _12755_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_238_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19470_ _06510_ _06516_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__nand2_1
XFILLER_19_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28668_ clknet_leaf_187_clk _02466_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[216\]
+ sky130_fd_sc_hd__dfrtp_1
X_16682_ _03975_ _04003_ _04004_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__and3_1
X_13894_ deser_A.serial_word\[55\] deser_A.shift_reg\[55\] net58 VGND VGND VPWR VPWR
+ _00720_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_238_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18421_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.A_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\]
+ systolic_inst.A_outs\[8\]\[1\] VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__and4_1
X_15633_ systolic_inst.B_outs\[13\]\[5\] systolic_inst.A_outs\[13\]\[6\] VGND VGND
+ VPWR VPWR _12688_ sky130_fd_sc_hd__nand2_1
X_27619_ clknet_leaf_318_clk _01417_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_234_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28599_ clknet_leaf_138_clk _02397_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[147\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18352_ _05491_ _05499_ _05504_ _05509_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__nand4_1
XFILLER_37_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15564_ systolic_inst.A_outs\[13\]\[4\] systolic_inst.B_outs\[13\]\[5\] VGND VGND
+ VPWR VPWR _12621_ sky130_fd_sc_hd__nand2_1
XFILLER_221_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ net118 _04560_ _04561_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__a21oi_1
X_14515_ _11692_ _11694_ VGND VGND VPWR VPWR _11695_ sky130_fd_sc_hd__nor2_1
XFILLER_159_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15495_ systolic_inst.A_outs\[13\]\[1\] systolic_inst.B_outs\[13\]\[6\] _12553_ VGND
+ VGND VPWR VPWR _12554_ sky130_fd_sc_hd__and3_1
X_18283_ _05447_ _05452_ _05454_ net66 VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__o211ai_1
XFILLER_203_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17234_ _04477_ _04493_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__xnor2_1
X_14446_ _11594_ _11596_ _11595_ VGND VGND VPWR VPWR _11628_ sky130_fd_sc_hd__o21ba_1
XFILLER_80_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17165_ net105 systolic_inst.acc_wires\[11\]\[29\] net62 _04448_ VGND VGND VPWR VPWR
+ _01263_ sky130_fd_sc_hd__a22o_1
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14377_ systolic_inst.B_outs\[15\]\[5\] systolic_inst.A_outs\[15\]\[5\] VGND VGND
+ VPWR VPWR _11561_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_185_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16116_ _13094_ _03501_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__xnor2_1
X_13328_ A_in\[37\] deser_A.word_buffer\[37\] net94 VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__mux2_1
XFILLER_155_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17096_ net105 systolic_inst.acc_wires\[11\]\[18\] net62 _04390_ VGND VGND VPWR VPWR
+ _01252_ sky130_fd_sc_hd__a22o_1
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16047_ _13043_ VGND VGND VPWR VPWR _13044_ sky130_fd_sc_hd__inv_2
X_13259_ deser_A.word_buffer\[97\] deser_A.serial_word\[97\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__mux2_1
XFILLER_143_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19806_ _06751_ _06766_ _06765_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__o21a_1
XFILLER_85_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17998_ _05188_ _05189_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__or2_1
XFILLER_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19737_ net106 _06739_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__nor2_1
XFILLER_96_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16949_ _04199_ _04241_ _04240_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__o21a_1
XFILLER_238_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_76_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_226_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19668_ _06654_ _06672_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__nor2_1
XFILLER_93_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18619_ _05744_ _05745_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__xnor2_1
X_19599_ net105 systolic_inst.acc_wires\[7\]\[29\] net62 _06626_ VGND VGND VPWR VPWR
+ _01519_ sky130_fd_sc_hd__a22o_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21630_ _08375_ _08411_ _08409_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__a21o_1
XFILLER_206_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21561_ net122 _08371_ _08372_ _08344_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__a31o_1
XFILLER_240_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23300_ systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[2\]
+ systolic_inst.B_outs\[0\]\[1\] VGND VGND VPWR VPWR _09930_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20512_ _07407_ _07409_ _07445_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__a21o_1
X_24280_ _10613_ systolic_inst.B_shift\[23\]\[3\] net72 VGND VGND VPWR VPWR _02213_
+ sky130_fd_sc_hd__mux2_1
X_21492_ systolic_inst.A_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[2\] VGND VGND VPWR
+ VPWR _08307_ sky130_fd_sc_hd__and2_1
XFILLER_53_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23231_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[24\]
+ VGND VGND VPWR VPWR _09880_ sky130_fd_sc_hd__nor2_1
XFILLER_193_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20443_ _07377_ _07378_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23162_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[1\]\[14\]
+ VGND VGND VPWR VPWR _09821_ sky130_fd_sc_hd__nand2_1
XFILLER_162_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20374_ _07259_ _07261_ _07310_ _07311_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__a211oi_1
Xclkload350 clknet_leaf_25_A_in_serial_clk VGND VGND VPWR VPWR clkload350/X sky130_fd_sc_hd__clkbuf_8
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload361 clknet_leaf_13_A_in_serial_clk VGND VGND VPWR VPWR clkload361/X sky130_fd_sc_hd__clkbuf_8
Xclkload372 clknet_leaf_3_B_in_serial_clk VGND VGND VPWR VPWR clkload372/Y sky130_fd_sc_hd__clkinv_4
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22113_ systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[3\]
+ systolic_inst.B_outs\[2\]\[0\] VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__a22o_1
Xclkload383 clknet_leaf_26_B_in_serial_clk VGND VGND VPWR VPWR clkload383/X sky130_fd_sc_hd__clkbuf_8
Xclkload80 clknet_leaf_21_clk VGND VGND VPWR VPWR clkload80/Y sky130_fd_sc_hd__inv_6
Xclkload394 clknet_leaf_16_B_in_serial_clk VGND VGND VPWR VPWR clkload394/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload91 clknet_leaf_317_clk VGND VGND VPWR VPWR clkload91/Y sky130_fd_sc_hd__inv_6
XFILLER_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27970_ clknet_leaf_165_clk _01768_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_23093_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[1\]\[4\]
+ VGND VGND VPWR VPWR _09762_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_168_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22044_ _08817_ _08818_ _08816_ VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__o21ai_1
X_26921_ clknet_leaf_4_A_in_serial_clk _00719_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29640_ clknet_leaf_29_B_in_serial_clk _03435_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_26852_ clknet_leaf_67_clk _00654_ net134 VGND VGND VPWR VPWR B_in\[124\] sky130_fd_sc_hd__dfrtp_1
XFILLER_125_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25803_ systolic_inst.acc_wires\[8\]\[23\] C_out\[279\] net28 VGND VGND VPWR VPWR
+ _03105_ sky130_fd_sc_hd__mux2_1
XFILLER_102_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29571_ clknet_leaf_21_B_in_serial_clk _03366_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_23995_ systolic_inst.B_shift\[9\]\[1\] B_in\[9\] _00008_ VGND VGND VPWR VPWR _10523_
+ sky130_fd_sc_hd__mux2_1
XFILLER_169_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26783_ clknet_leaf_61_clk _00585_ net143 VGND VGND VPWR VPWR B_in\[55\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_67_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_29_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28522_ clknet_leaf_154_clk _02320_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25734_ systolic_inst.acc_wires\[6\]\[18\] C_out\[210\] net46 VGND VGND VPWR VPWR
+ _03036_ sky130_fd_sc_hd__mux2_1
X_22946_ _09622_ _09623_ VGND VGND VPWR VPWR _09624_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28453_ clknet_leaf_131_clk _02251_ net144 VGND VGND VPWR VPWR ser_C.shift_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22877_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[7\] VGND VGND VPWR
+ VPWR _09557_ sky130_fd_sc_hd__nand2_4
X_25665_ systolic_inst.acc_wires\[4\]\[13\] C_out\[141\] net30 VGND VGND VPWR VPWR
+ _02967_ sky130_fd_sc_hd__mux2_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27404_ clknet_leaf_229_clk _01202_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_21828_ _08629_ _08630_ VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__and2b_1
XFILLER_93_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24616_ net110 ser_C.shift_reg\[136\] VGND VGND VPWR VPWR _10778_ sky130_fd_sc_hd__and2_1
XFILLER_231_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25596_ systolic_inst.acc_wires\[2\]\[8\] C_out\[72\] net34 VGND VGND VPWR VPWR _02898_
+ sky130_fd_sc_hd__mux2_1
X_28384_ clknet_leaf_32_clk _02182_ VGND VGND VPWR VPWR systolic_inst.A_shift\[18\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24547_ C_out\[100\] net99 net79 ser_C.shift_reg\[100\] _10743_ VGND VGND VPWR VPWR
+ _02350_ sky130_fd_sc_hd__a221o_1
X_27335_ clknet_leaf_289_clk _01133_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_240_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21759_ _08556_ _08564_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__nand2_1
XFILLER_145_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14300_ _11447_ _11485_ VGND VGND VPWR VPWR _11486_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15280_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[20\]
+ VGND VGND VPWR VPWR _12374_ sky130_fd_sc_hd__nand2_1
X_24478_ net112 ser_C.shift_reg\[67\] VGND VGND VPWR VPWR _10709_ sky130_fd_sc_hd__and2_1
Xwire112 net114 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_12
XFILLER_200_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27266_ clknet_leaf_268_clk _01064_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29005_ clknet_leaf_105_clk _02803_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14231_ _11413_ _11414_ _11418_ VGND VGND VPWR VPWR _11419_ sky130_fd_sc_hd__nand3_2
X_23429_ _10052_ _10053_ _10010_ _10012_ VGND VGND VPWR VPWR _10055_ sky130_fd_sc_hd__a211oi_2
X_26217_ clknet_leaf_9_A_in_serial_clk _00025_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_27197_ clknet_leaf_262_clk _00995_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_153_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_242_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26148_ deser_B.serial_word\[103\] deser_B.shift_reg\[103\] _00001_ VGND VGND VPWR
+ VPWR _03450_ sky130_fd_sc_hd__mux2_1
X_14162_ _11349_ _11352_ VGND VGND VPWR VPWR _11353_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_242_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_242_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13113_ systolic_inst.A_outs\[0\]\[6\] VGND VGND VPWR VPWR _11269_ sky130_fd_sc_hd__inv_2
XFILLER_153_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26079_ deser_B.serial_word\[34\] deser_B.shift_reg\[34\] net55 VGND VGND VPWR VPWR
+ _03381_ sky130_fd_sc_hd__mux2_1
X_14093_ deser_B.shift_reg\[127\] net4 net126 VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__mux2_1
X_18970_ _06066_ _06065_ systolic_inst.acc_wires\[8\]\[24\] net108 VGND VGND VPWR
+ VPWR _01450_ sky130_fd_sc_hd__a2bb2o_1
Xload_slew106 net107 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_16
XFILLER_112_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17921_ _05110_ _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__nor2_1
XFILLER_106_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17852_ net107 _05047_ _05048_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__or3_1
XFILLER_79_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16803_ _04122_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__inv_2
X_17783_ _04994_ _04998_ _04999_ net60 VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_58_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14995_ _12113_ _12114_ VGND VGND VPWR VPWR _12115_ sky130_fd_sc_hd__nor2_1
X_19522_ _06559_ _06561_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__xnor2_1
X_16734_ _04027_ _04029_ _04028_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__o21bai_1
XFILLER_219_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13946_ deser_A.serial_word\[107\] deser_A.shift_reg\[107\] net57 VGND VGND VPWR
+ VPWR _00772_ sky130_fd_sc_hd__mux2_1
XFILLER_235_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19453_ _06497_ _06500_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__nand2_1
X_16665_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[3\] _03972_ _03970_
+ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__a31o_1
XFILLER_207_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13877_ deser_A.serial_word\[38\] deser_A.shift_reg\[38\] net58 VGND VGND VPWR VPWR
+ _00703_ sky130_fd_sc_hd__mux2_1
XFILLER_201_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18404_ systolic_inst.A_outs\[8\]\[1\] systolic_inst.A_shift\[16\]\[1\] net121 VGND
+ VGND VPWR VPWR _01395_ sky130_fd_sc_hd__mux2_1
X_15616_ _12670_ _12671_ VGND VGND VPWR VPWR _12672_ sky130_fd_sc_hd__or2_2
X_19384_ _06440_ _06441_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__and2b_1
XFILLER_61_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16596_ _03923_ _03921_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[1\]
+ net105 VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18335_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__inv_2
XFILLER_91_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15547_ _12603_ _12604_ VGND VGND VPWR VPWR _12605_ sky130_fd_sc_hd__nor2_1
XFILLER_37_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18266_ _05431_ _05436_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__nor2_1
XFILLER_198_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15478_ _12529_ _12531_ VGND VGND VPWR VPWR _12537_ sky130_fd_sc_hd__nor2_1
XFILLER_175_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17217_ _04466_ _04477_ _04478_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__and3_1
X_14429_ _11554_ _11611_ VGND VGND VPWR VPWR _11612_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18197_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[9\]\[0\]
+ _05379_ _05380_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__and4_1
XFILLER_239_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17148_ net105 systolic_inst.acc_wires\[11\]\[26\] net62 _04434_ VGND VGND VPWR VPWR
+ _01260_ sky130_fd_sc_hd__a22o_1
XFILLER_128_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17079_ _04374_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__and2_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20090_ _07061_ _07066_ _07067_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__nand3_1
XFILLER_83_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
X_22800_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[5\] systolic_inst.A_outs\[1\]\[6\]
+ systolic_inst.B_outs\[1\]\[1\] VGND VGND VPWR VPWR _09482_ sky130_fd_sc_hd__a22o_1
XFILLER_38_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23780_ _10375_ _10376_ _10383_ VGND VGND VPWR VPWR _10384_ sky130_fd_sc_hd__a21o_1
X_20992_ _07835_ _07865_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__nand2b_1
XFILLER_214_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22731_ _09407_ _09413_ _09415_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__and3_1
XFILLER_53_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25450_ _11193_ _11196_ _11197_ systolic_inst.cycle_cnt\[5\] VGND VGND VPWR VPWR
+ _02799_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_172_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22662_ _09359_ _09362_ _09365_ _09368_ VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_172_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24401_ C_out\[27\] _11302_ net82 ser_C.shift_reg\[27\] _10670_ VGND VGND VPWR VPWR
+ _02277_ sky130_fd_sc_hd__a221o_1
XFILLER_181_1330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21613_ _08388_ _08422_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_1412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25381_ systolic_inst.B_shift\[18\]\[6\] B_in\[54\] net59 VGND VGND VPWR VPWR _11160_
+ sky130_fd_sc_hd__mux2_1
XFILLER_240_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22593_ _09309_ _09311_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__xor2_1
XFILLER_16_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27120_ clknet_leaf_0_B_in_serial_clk _00918_ net134 VGND VGND VPWR VPWR deser_B.shift_reg\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24332_ _10639_ systolic_inst.A_shift\[9\]\[5\] net70 VGND VGND VPWR VPWR _02239_
+ sky130_fd_sc_hd__mux2_1
XFILLER_221_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21544_ systolic_inst.A_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[2\] systolic_inst.B_outs\[3\]\[3\]
+ systolic_inst.B_outs\[3\]\[4\] VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__and4_1
XFILLER_55_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27051_ clknet_leaf_24_B_in_serial_clk _00849_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24263_ systolic_inst.A_shift\[16\]\[6\] net70 net83 systolic_inst.A_shift\[17\]\[6\]
+ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__a22o_1
X_21475_ systolic_inst.B_outs\[2\]\[3\] systolic_inst.B_shift\[2\]\[3\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__mux2_1
XFILLER_153_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26002_ systolic_inst.acc_wires\[14\]\[30\] ser_C.parallel_data\[478\] net24 VGND
+ VGND VPWR VPWR _03304_ sky130_fd_sc_hd__mux2_1
XFILLER_101_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23214_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[22\]
+ VGND VGND VPWR VPWR _09865_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_116_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20426_ _07322_ _07360_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__and2_1
XFILLER_135_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24194_ systolic_inst.B_shift\[22\]\[1\] net72 _11333_ B_in\[113\] VGND VGND VPWR
+ VPWR _02155_ sky130_fd_sc_hd__a22o_1
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23145_ _09796_ _09801_ _09802_ VGND VGND VPWR VPWR _09806_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_112_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20357_ systolic_inst.B_outs\[5\]\[3\] systolic_inst.A_outs\[5\]\[4\] VGND VGND VPWR
+ VPWR _07295_ sky130_fd_sc_hd__nand2_1
Xclkload180 clknet_leaf_236_clk VGND VGND VPWR VPWR clkload180/X sky130_fd_sc_hd__clkbuf_8
XFILLER_101_1088 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload191 clknet_leaf_60_clk VGND VGND VPWR VPWR clkload191/Y sky130_fd_sc_hd__bufinv_16
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23076_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[1\]\[0\]
+ _09744_ _09745_ VGND VGND VPWR VPWR _09748_ sky130_fd_sc_hd__a22o_1
X_27953_ clknet_leaf_171_clk _01751_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20288_ _07209_ _07211_ _07210_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__a21bo_1
XFILLER_62_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22027_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[23\]
+ _08787_ _08795_ _08797_ VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__a2111o_1
X_26904_ clknet_leaf_16_A_in_serial_clk _00702_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_222_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27884_ clknet_leaf_310_clk _01682_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29623_ clknet_leaf_8_B_in_serial_clk _03418_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_236_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26835_ clknet_leaf_89_clk _00637_ net5 VGND VGND VPWR VPWR B_in\[107\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ B_in\[107\] deser_B.word_buffer\[107\] net90 VGND VGND VPWR VPWR _00637_
+ sky130_fd_sc_hd__mux2_1
X_29554_ clknet_leaf_18_B_in_serial_clk _03349_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_235_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26766_ clknet_leaf_81_clk _00568_ net153 VGND VGND VPWR VPWR B_in\[38\] sky130_fd_sc_hd__dfrtp_1
X_14780_ _11905_ _11906_ VGND VGND VPWR VPWR _11907_ sky130_fd_sc_hd__nand2_1
X_23978_ _10514_ systolic_inst.B_shift\[8\]\[0\] net72 VGND VGND VPWR VPWR _02010_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28505_ clknet_leaf_108_clk _02303_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_217_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13731_ B_in\[38\] deser_B.word_buffer\[38\] net90 VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__mux2_1
X_25717_ systolic_inst.acc_wires\[6\]\[1\] C_out\[193\] net47 VGND VGND VPWR VPWR
+ _03019_ sky130_fd_sc_hd__mux2_1
XFILLER_17_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22929_ _09570_ _09571_ _09573_ VGND VGND VPWR VPWR _09608_ sky130_fd_sc_hd__o21a_1
X_29485_ clknet_leaf_281_clk _03283_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_231_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26697_ clknet_leaf_5_B_in_serial_clk _00500_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_231_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28436_ clknet_leaf_25_clk _02234_ VGND VGND VPWR VPWR systolic_inst.A_shift\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16450_ _03812_ _03814_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__nor2_1
X_25648_ systolic_inst.acc_wires\[3\]\[28\] C_out\[124\] net49 VGND VGND VPWR VPWR
+ _02950_ sky130_fd_sc_hd__mux2_1
XFILLER_204_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13662_ deser_B.word_buffer\[98\] deser_B.serial_word\[98\] net123 VGND VGND VPWR
+ VPWR _00499_ sky130_fd_sc_hd__mux2_1
XFILLER_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15401_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[2\] VGND VGND
+ VPWR VPWR _12463_ sky130_fd_sc_hd__and2_1
XFILLER_73_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13593_ deser_B.word_buffer\[29\] deser_B.serial_word\[29\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__mux2_1
XFILLER_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16381_ net67 _03753_ _03755_ systolic_inst.acc_wires\[12\]\[2\] net108 VGND VGND
+ VPWR VPWR _01172_ sky130_fd_sc_hd__a32o_1
X_28367_ clknet_leaf_5_clk _02165_ VGND VGND VPWR VPWR systolic_inst.A_shift\[20\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25579_ systolic_inst.acc_wires\[1\]\[23\] C_out\[55\] net53 VGND VGND VPWR VPWR
+ _02881_ sky130_fd_sc_hd__mux2_1
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18120_ _05307_ _05308_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_26_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27318_ clknet_leaf_289_clk _01116_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_15332_ systolic_inst.acc_wires\[14\]\[26\] systolic_inst.acc_wires\[14\]\[27\] systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12418_ sky130_fd_sc_hd__o21a_1
XFILLER_223_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28298_ clknet_leaf_127_clk _02096_ VGND VGND VPWR VPWR systolic_inst.B_shift\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18051_ _05190_ _05207_ _05205_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__o21a_1
X_15263_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[17\]
+ VGND VGND VPWR VPWR _12360_ sky130_fd_sc_hd__xor2_2
X_27249_ clknet_leaf_275_clk _01047_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_229_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17002_ _04303_ _04304_ _04302_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__a21bo_1
X_14214_ _11402_ _11401_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[5\]
+ net107 VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_158_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15194_ _12292_ _12296_ _12298_ _12299_ VGND VGND VPWR VPWR _12301_ sky130_fd_sc_hd__o211ai_2
XANTENNA_6 systolic_inst.A_outs\[10\]\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14145_ net107 systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[1\] _11335_
+ _11337_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__a22o_1
XFILLER_193_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14076_ deser_B.shift_reg\[110\] deser_B.shift_reg\[111\] deser_B.receiving VGND
+ VGND VPWR VPWR _00902_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18953_ _06050_ _06051_ _06049_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__o21ai_1
XFILLER_193_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17904_ _05086_ _05098_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__xnor2_1
X_18884_ _05992_ _05991_ systolic_inst.acc_wires\[8\]\[12\] net108 VGND VGND VPWR
+ VPWR _01438_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_230_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17835_ _05030_ _05031_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__nand2_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_176_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17766_ _04983_ _04986_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__xor2_1
X_14978_ _12056_ _12058_ _12096_ VGND VGND VPWR VPWR _12099_ sky130_fd_sc_hd__a21o_1
X_19505_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[15\]
+ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__and2_1
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16717_ _04031_ _04037_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__xnor2_1
X_13929_ deser_A.serial_word\[90\] deser_A.shift_reg\[90\] net57 VGND VGND VPWR VPWR
+ _00755_ sky130_fd_sc_hd__mux2_1
X_17697_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[18\]
+ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__or2_1
XFILLER_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19436_ _06486_ _06487_ _06479_ _06483_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__a211o_1
XFILLER_222_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16648_ systolic_inst.A_outs\[11\]\[2\] systolic_inst.B_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\]
+ systolic_inst.A_outs\[11\]\[1\] VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__a22o_1
XFILLER_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_783 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19367_ _06425_ _06426_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__nor2_1
XFILLER_241_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16579_ systolic_inst.A_outs\[11\]\[4\] systolic_inst.A_outs\[10\]\[4\] net118 VGND
+ VGND VPWR VPWR _01206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_214_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18318_ _05481_ _05482_ _05483_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__nand3_1
XFILLER_241_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19298_ _06319_ _06321_ _06358_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__nand3_1
XFILLER_175_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18249_ _05423_ _05424_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21260_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[4\]\[0\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__a22o_1
XFILLER_116_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20211_ systolic_inst.acc_wires\[6\]\[28\] systolic_inst.acc_wires\[6\]\[29\] systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21191_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[12\] _08059_ net117
+ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_239_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20142_ _07111_ _07113_ _07110_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__o21ai_1
XFILLER_131_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_161_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20073_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[6\]\[8\]
+ _07053_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__and3_1
XFILLER_44_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24950_ net111 ser_C.shift_reg\[303\] VGND VGND VPWR VPWR _10945_ sky130_fd_sc_hd__and2_1
XFILLER_170_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23901_ _10483_ systolic_inst.B_shift\[13\]\[2\] net72 VGND VGND VPWR VPWR _01964_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24881_ C_out\[267\] net101 net75 ser_C.shift_reg\[267\] _10910_ VGND VGND VPWR VPWR
+ _02517_ sky130_fd_sc_hd__a221o_1
XFILLER_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26620_ clknet_leaf_22_B_in_serial_clk _00423_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23832_ _11258_ systolic_inst.acc_wires\[0\]\[21\] net64 _10427_ VGND VGND VPWR VPWR
+ _01951_ sky130_fd_sc_hd__a22o_1
XFILLER_214_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23763_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[0\]\[11\]
+ VGND VGND VPWR VPWR _10369_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26551_ clknet_leaf_26_A_in_serial_clk _00354_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20975_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[6\] VGND VGND VPWR
+ VPWR _07849_ sky130_fd_sc_hd__nand2_1
X_25502_ systolic_inst.cycle_cnt\[24\] systolic_inst.cycle_cnt\[23\] _11228_ VGND
+ VGND VPWR VPWR _11231_ sky130_fd_sc_hd__and3_1
XFILLER_214_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22714_ _09386_ _09388_ _09399_ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__and3_1
X_29270_ clknet_leaf_194_clk _03068_ net146 VGND VGND VPWR VPWR C_out\[242\] sky130_fd_sc_hd__dfrtp_1
X_23694_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[0\]\[1\]
+ VGND VGND VPWR VPWR _10310_ sky130_fd_sc_hd__and2_1
X_26482_ clknet_leaf_12_A_in_serial_clk _00285_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28221_ clknet_leaf_99_clk _02019_ VGND VGND VPWR VPWR systolic_inst.B_shift\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25433_ systolic_inst.ce_local _11307_ systolic_inst.cycle_cnt\[0\] VGND VGND VPWR
+ VPWR _02794_ sky130_fd_sc_hd__mux2_1
X_22645_ _09348_ _09352_ _09349_ VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__a21bo_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28152_ clknet_leaf_102_clk _01950_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_118_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25364_ net112 ser_C.shift_reg\[510\] VGND VGND VPWR VPWR _11152_ sky130_fd_sc_hd__and2_1
X_22576_ _09285_ _09291_ _09292_ VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__o21ba_1
XFILLER_139_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27103_ clknet_leaf_10_B_in_serial_clk _00901_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_194_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21527_ _08316_ _08319_ _08337_ VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_114_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24315_ systolic_inst.A_shift\[11\]\[5\] A_in\[45\] net59 VGND VGND VPWR VPWR _10631_
+ sky130_fd_sc_hd__mux2_1
X_28083_ clknet_leaf_115_clk _01881_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25295_ ser_C.parallel_data\[474\] net102 net74 ser_C.shift_reg\[474\] _11117_ VGND
+ VGND VPWR VPWR _02724_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27034_ clknet_leaf_13_B_in_serial_clk _00832_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24246_ _10608_ systolic_inst.A_shift\[18\]\[6\] net70 VGND VGND VPWR VPWR _02184_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21458_ _08288_ _08291_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__or2_1
XFILLER_119_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20409_ _07327_ _07345_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_224_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24177_ systolic_inst.A_shift\[25\]\[0\] net70 net83 systolic_inst.A_shift\[26\]\[0\]
+ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__a22o_1
XFILLER_108_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput10 net10 VGND VGND VPWR VPWR done sky130_fd_sc_hd__buf_1
Xoutput8 net8 VGND VGND VPWR VPWR C_out_serial_clk sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_224_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21389_ _08212_ _08213_ _08218_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__and3_1
XFILLER_162_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23128_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[1\]\[8\]
+ _09788_ VGND VGND VPWR VPWR _09792_ sky130_fd_sc_hd__and3_1
XFILLER_150_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28985_ clknet_leaf_24_clk _02783_ VGND VGND VPWR VPWR systolic_inst.A_shift\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_220_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27936_ clknet_leaf_171_clk _01734_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_23059_ _09731_ _09732_ VGND VGND VPWR VPWR _09734_ sky130_fd_sc_hd__nand2_1
XFILLER_27_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15950_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[30\]
+ VGND VGND VPWR VPWR _12970_ sky130_fd_sc_hd__or2_1
XFILLER_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14901_ _11990_ _12022_ VGND VGND VPWR VPWR _12024_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27867_ clknet_leaf_145_clk _01665_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_15881_ net108 systolic_inst.acc_wires\[13\]\[19\] net67 _12911_ VGND VGND VPWR VPWR
+ _01125_ sky130_fd_sc_hd__a22o_1
XFILLER_40_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29606_ clknet_leaf_23_B_in_serial_clk _03401_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_17620_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[10\]\[7\]
+ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__nand2_1
X_26818_ clknet_leaf_66_clk _00620_ net135 VGND VGND VPWR VPWR B_in\[90\] sky130_fd_sc_hd__dfrtp_1
X_14832_ _11933_ _11955_ VGND VGND VPWR VPWR _11957_ sky130_fd_sc_hd__xnor2_1
X_27798_ clknet_leaf_48_clk _01596_ net137 VGND VGND VPWR VPWR systolic_inst.B_outs\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_64_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29537_ clknet_leaf_256_clk _03335_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[509\]
+ sky130_fd_sc_hd__dfrtp_1
X_17551_ _04776_ _04779_ _04801_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__a21oi_1
X_26749_ clknet_leaf_53_clk _00551_ net143 VGND VGND VPWR VPWR B_in\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14763_ systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[1\] VGND VGND
+ VPWR VPWR _11891_ sky130_fd_sc_hd__nand2_1
XFILLER_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16502_ _03859_ _03858_ systolic_inst.acc_wires\[12\]\[19\] net108 VGND VGND VPWR
+ VPWR _01189_ sky130_fd_sc_hd__a2bb2o_1
X_13714_ B_in\[21\] deser_B.word_buffer\[21\] net86 VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__mux2_1
XFILLER_17_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29468_ clknet_leaf_287_clk _03266_ net136 VGND VGND VPWR VPWR ser_C.parallel_data\[440\]
+ sky130_fd_sc_hd__dfrtp_1
X_17482_ _04701_ _04705_ _04733_ _04735_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__nor4_1
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14694_ _11846_ _11847_ VGND VGND VPWR VPWR _11848_ sky130_fd_sc_hd__or2_1
XFILLER_71_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19221_ _06283_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28419_ clknet_leaf_70_clk _02217_ VGND VGND VPWR VPWR systolic_inst.B_shift\[23\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16433_ _03796_ _03798_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__nand2_1
XFILLER_73_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13645_ deser_B.word_buffer\[81\] deser_B.serial_word\[81\] net123 VGND VGND VPWR
+ VPWR _00482_ sky130_fd_sc_hd__mux2_1
X_29399_ clknet_leaf_239_clk _03197_ net145 VGND VGND VPWR VPWR C_out\[371\] sky130_fd_sc_hd__dfrtp_1
XFILLER_147_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19152_ _06182_ _06217_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16364_ _03741_ _03734_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ net108 VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13576_ deser_B.word_buffer\[12\] deser_B.serial_word\[12\] net124 VGND VGND VPWR
+ VPWR _00413_ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_3__f_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_2_3__leaf_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__inv_2
X_15315_ _12404_ _12403_ systolic_inst.acc_wires\[14\]\[24\] net107 VGND VGND VPWR
+ VPWR _01066_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19083_ systolic_inst.A_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[3\]
+ systolic_inst.B_outs\[7\]\[4\] VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__and4_1
XFILLER_125_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16295_ _03675_ _03674_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__and2b_1
XFILLER_185_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18034_ systolic_inst.A_outs\[9\]\[6\] _05224_ _05223_ VGND VGND VPWR VPWR _05225_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_184_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15246_ _12342_ _12344_ VGND VGND VPWR VPWR _12346_ sky130_fd_sc_hd__or2_1
XFILLER_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15177_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[14\]\[5\]
+ VGND VGND VPWR VPWR _12286_ sky130_fd_sc_hd__and2_1
XFILLER_67_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_947 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14128_ systolic_inst.A_outs\[15\]\[4\] systolic_inst.A_outs\[14\]\[4\] net118 VGND
+ VGND VPWR VPWR _00950_ sky130_fd_sc_hd__mux2_1
X_19985_ _06977_ _06978_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__a21oi_1
XFILLER_193_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_207_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14059_ deser_B.shift_reg\[93\] deser_B.shift_reg\[94\] net126 VGND VGND VPWR VPWR
+ _00885_ sky130_fd_sc_hd__mux2_1
X_18936_ _06035_ _06036_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__and2_1
XFILLER_234_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18867_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[8\]\[11\]
+ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__or2_1
XFILLER_132_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17818_ systolic_inst.A_outs\[9\]\[0\] systolic_inst.A_outs\[9\]\[1\] systolic_inst.B_outs\[9\]\[2\]
+ systolic_inst.B_outs\[9\]\[3\] VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__and4_1
XFILLER_95_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18798_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] _05919_ net117
+ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__mux2_1
XFILLER_94_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17749_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[26\]
+ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__or2_1
XFILLER_70_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20760_ _07667_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__inv_2
XFILLER_90_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19419_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[7\]\[3\]
+ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__and2_1
XFILLER_165_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20691_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[5\]\[11\]
+ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22430_ _09169_ _09168_ VGND VGND VPWR VPWR _09170_ sky130_fd_sc_hd__and2b_1
XFILLER_195_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22361_ _09102_ _09101_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__nand2b_1
XFILLER_163_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24100_ _10559_ systolic_inst.B_shift\[19\]\[5\] net71 VGND VGND VPWR VPWR _02087_
+ sky130_fd_sc_hd__mux2_1
X_21312_ _08166_ _08167_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__or2_1
X_25080_ net112 ser_C.shift_reg\[368\] VGND VGND VPWR VPWR _11010_ sky130_fd_sc_hd__and2_1
X_22292_ _09035_ _09034_ VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__nand2b_1
XFILLER_11_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24031_ systolic_inst.B_shift\[8\]\[3\] B_in\[35\] _00008_ VGND VGND VPWR VPWR _10533_
+ sky130_fd_sc_hd__mux2_1
X_21243_ _08084_ _08107_ _08108_ _08106_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__a31o_1
XFILLER_163_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21174_ _08038_ _08041_ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__or2_1
XFILLER_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20125_ _07100_ _07101_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__nand2_1
XFILLER_131_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_280_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_280_clk
+ sky130_fd_sc_hd__clkbuf_8
X_28770_ clknet_leaf_225_clk _02568_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[318\]
+ sky130_fd_sc_hd__dfrtp_1
X_25982_ systolic_inst.acc_wires\[14\]\[10\] ser_C.parallel_data\[458\] net26 VGND
+ VGND VPWR VPWR _03284_ sky130_fd_sc_hd__mux2_1
XFILLER_217_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27721_ clknet_leaf_189_clk _01519_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20056_ _07042_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__inv_2
XFILLER_58_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24933_ C_out\[293\] net102 net74 ser_C.shift_reg\[293\] _10936_ VGND VGND VPWR VPWR
+ _02543_ sky130_fd_sc_hd__a221o_1
XFILLER_219_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27652_ clknet_leaf_312_clk _01450_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24864_ net110 ser_C.shift_reg\[260\] VGND VGND VPWR VPWR _10902_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26603_ clknet_leaf_16_B_in_serial_clk _00406_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23815_ _10404_ _10406_ _10413_ VGND VGND VPWR VPWR _10414_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27583_ clknet_leaf_219_clk _01381_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_23__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_23__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_24795_ C_out\[224\] net99 net79 ser_C.shift_reg\[224\] _10867_ VGND VGND VPWR VPWR
+ _02474_ sky130_fd_sc_hd__a221o_1
XFILLER_96_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29322_ clknet_leaf_298_clk _03120_ net138 VGND VGND VPWR VPWR C_out\[294\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26534_ clknet_leaf_17_A_in_serial_clk _00337_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_23746_ _10354_ _10353_ systolic_inst.acc_wires\[0\]\[8\] _11258_ VGND VGND VPWR
+ VPWR _01938_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20958_ net108 _07831_ _07832_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__or3b_1
XFILLER_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29253_ clknet_leaf_200_clk _03051_ net147 VGND VGND VPWR VPWR C_out\[225\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26465_ clknet_leaf_1_A_in_serial_clk _00272_ net132 VGND VGND VPWR VPWR deser_A.bit_idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_23677_ _10269_ _10294_ VGND VGND VPWR VPWR _10296_ sky130_fd_sc_hd__or2_1
X_20889_ _07739_ _07745_ _07744_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__a21oi_1
XFILLER_224_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28204_ clknet_leaf_99_clk _02002_ VGND VGND VPWR VPWR systolic_inst.B_shift\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_201_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25416_ _11177_ systolic_inst.A_shift\[1\]\[7\] net71 VGND VGND VPWR VPWR _02785_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ deser_A.bit_idx\[3\] deser_A.bit_idx\[2\] _11309_ deser_A.bit_idx\[4\] VGND
+ VGND VPWR VPWR _11315_ sky130_fd_sc_hd__a31o_1
X_22628_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[24\]
+ VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__and2_1
X_29184_ clknet_leaf_135_clk _02982_ net142 VGND VGND VPWR VPWR C_out\[156\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26396_ clknet_leaf_27_clk _00203_ net137 VGND VGND VPWR VPWR A_in\[64\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28135_ clknet_leaf_127_clk _01933_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13361_ A_in\[70\] deser_A.word_buffer\[70\] net96 VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__mux2_1
X_22559_ net60 _09282_ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__nor2_1
XFILLER_127_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25347_ ser_C.parallel_data\[500\] net98 net78 ser_C.shift_reg\[500\] _11143_ VGND
+ VGND VPWR VPWR _02750_ sky130_fd_sc_hd__a221o_1
XFILLER_220_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15100_ _12146_ _12186_ _12185_ VGND VGND VPWR VPWR _12217_ sky130_fd_sc_hd__a21bo_1
X_28066_ clknet_leaf_120_clk _01864_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_177_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13292_ A_in\[1\] deser_A.word_buffer\[1\] net93 VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__mux2_1
X_16080_ _13044_ _13075_ VGND VGND VPWR VPWR _13076_ sky130_fd_sc_hd__xnor2_1
X_25278_ net111 ser_C.shift_reg\[467\] VGND VGND VPWR VPWR _11109_ sky130_fd_sc_hd__and2_1
XFILLER_177_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27017_ clknet_leaf_22_B_in_serial_clk _00815_ net137 VGND VGND VPWR VPWR deser_B.shift_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_15031_ _12148_ _12149_ VGND VGND VPWR VPWR _12150_ sky130_fd_sc_hd__nor2_1
X_24229_ systolic_inst.A_shift\[20\]\[6\] A_in\[78\] net59 VGND VGND VPWR VPWR _10600_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_271_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_271_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19770_ _06742_ _06771_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__nand2b_1
XFILLER_231_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28968_ clknet_leaf_53_clk _02766_ VGND VGND VPWR VPWR systolic_inst.B_shift\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16982_ _04290_ _04291_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__a21o_1
XFILLER_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18721_ _05813_ _05815_ _05844_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__nand3_1
X_27919_ clknet_leaf_145_clk _01717_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_15933_ net107 systolic_inst.acc_wires\[13\]\[27\] net67 _12955_ VGND VGND VPWR VPWR
+ _01133_ sky130_fd_sc_hd__a22o_1
XFILLER_231_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28899_ clknet_leaf_279_clk _02697_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[447\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_202_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18652_ _05770_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__nand2_1
XFILLER_236_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15864_ net61 _12897_ VGND VGND VPWR VPWR _12898_ sky130_fd_sc_hd__nor2_1
XFILLER_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17603_ _04847_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__inv_2
XFILLER_149_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14815_ _11920_ _11939_ VGND VGND VPWR VPWR _11940_ sky130_fd_sc_hd__nand2_1
XFILLER_236_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18583_ _05709_ _05710_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_194_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[13\]\[7\]
+ VGND VGND VPWR VPWR _12838_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_194_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17534_ _04741_ _04755_ _04753_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__o21a_1
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14746_ systolic_inst.A_outs\[14\]\[6\] systolic_inst.A_outs\[13\]\[6\] net116 VGND
+ VGND VPWR VPWR _01016_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_190_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17465_ _04715_ _04718_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_190_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14677_ _11831_ _11832_ VGND VGND VPWR VPWR _11833_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_211_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19204_ _06266_ _06267_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__xor2_1
XFILLER_242_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16416_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[12\]\[8\]
+ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__xor2_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13628_ deser_B.word_buffer\[64\] deser_B.serial_word\[64\] net123 VGND VGND VPWR
+ VPWR _00465_ sky130_fd_sc_hd__mux2_1
XFILLER_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17396_ _04648_ _04651_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19135_ systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[6\] systolic_inst.A_outs\[7\]\[7\]
+ systolic_inst.B_outs\[7\]\[0\] VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__a22o_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16347_ _03723_ _03724_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__and2b_1
X_13559_ deser_A.shift_reg\[123\] deser_A.shift_reg\[124\] net130 VGND VGND VPWR VPWR
+ _00396_ sky130_fd_sc_hd__mux2_1
XFILLER_185_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19066_ _06133_ _06134_ _06115_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__o21ai_1
XFILLER_118_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16278_ _03516_ _03657_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__nand2_2
XFILLER_145_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18017_ _05169_ _05170_ _05172_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__o21a_1
X_15229_ _12330_ VGND VGND VPWR VPWR _12331_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_209_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_262_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_262_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_87_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19968_ _06962_ _06963_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__nand2b_1
XFILLER_234_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18919_ _06014_ _06017_ _06016_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__o21a_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_143_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19899_ systolic_inst.A_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[5\] systolic_inst.B_outs\[6\]\[6\]
+ systolic_inst.B_outs\[6\]\[7\] VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_143_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1026 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21930_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[3\]\[8\]
+ _08715_ _08714_ VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__a31o_1
XFILLER_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21861_ _08586_ _08648_ _08646_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20812_ _07705_ _07708_ _07707_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__o21a_1
X_23600_ systolic_inst.A_outs\[0\]\[5\] systolic_inst.B_outs\[0\]\[6\] _10193_ _10154_
+ VGND VGND VPWR VPWR _10221_ sky130_fd_sc_hd__a31o_1
X_24580_ net114 ser_C.shift_reg\[118\] VGND VGND VPWR VPWR _10760_ sky130_fd_sc_hd__and2_1
X_21792_ _08563_ _08565_ _08596_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__a21o_1
XFILLER_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20743_ _07644_ _07646_ _07653_ VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__a21oi_1
X_23531_ systolic_inst.B_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[7\]
+ VGND VGND VPWR VPWR _10154_ sky130_fd_sc_hd__and3_2
XFILLER_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23462_ _10077_ _10085_ VGND VGND VPWR VPWR _10087_ sky130_fd_sc_hd__or2_1
X_26250_ clknet_leaf_10_A_in_serial_clk _00058_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_20674_ _07594_ _07593_ systolic_inst.acc_wires\[5\]\[8\] net109 VGND VGND VPWR VPWR
+ _01626_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_177_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22413_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[12\] _09153_ net122
+ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__mux2_1
X_25201_ C_out\[427\] net101 net73 ser_C.shift_reg\[427\] _11070_ VGND VGND VPWR VPWR
+ _02677_ sky130_fd_sc_hd__a221o_1
X_26181_ ser_C.bit_idx\[3\] _11247_ _11249_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__a21oi_1
X_23393_ _09984_ _10018_ VGND VGND VPWR VPWR _10020_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22344_ _09050_ _09051_ _09048_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__a21o_1
X_25132_ net110 ser_C.shift_reg\[394\] VGND VGND VPWR VPWR _11036_ sky130_fd_sc_hd__and2_1
XFILLER_152_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25063_ C_out\[358\] net98 net78 ser_C.shift_reg\[358\] _11001_ VGND VGND VPWR VPWR
+ _02608_ sky130_fd_sc_hd__a221o_1
X_22275_ net122 _09017_ _09018_ _09019_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__a31o_1
XFILLER_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24014_ systolic_inst.B_shift\[7\]\[5\] _11332_ net83 systolic_inst.B_shift\[11\]\[5\]
+ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__a22o_1
XFILLER_219_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21226_ _08089_ _08091_ _08041_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_93_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_253_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_253_clk
+ sky130_fd_sc_hd__clkbuf_8
X_28822_ clknet_leaf_240_clk _02620_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[370\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21157_ _07990_ _07993_ _07996_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20108_ _07085_ _07086_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__and2_1
X_28753_ clknet_leaf_220_clk _02551_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[301\]
+ sky130_fd_sc_hd__dfrtp_1
X_21088_ _07917_ _07958_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__xnor2_1
X_25965_ systolic_inst.acc_wires\[13\]\[25\] ser_C.parallel_data\[441\] net19 VGND
+ VGND VPWR VPWR _03267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27704_ clknet_leaf_191_clk _01502_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20039_ _07021_ _07022_ _07020_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__a21bo_1
XFILLER_4_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24916_ net110 ser_C.shift_reg\[286\] VGND VGND VPWR VPWR _10928_ sky130_fd_sc_hd__and2_1
X_28684_ clknet_leaf_194_clk _02482_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[232\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_115_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25896_ systolic_inst.acc_wires\[11\]\[20\] C_out\[372\] net41 VGND VGND VPWR VPWR
+ _03198_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27635_ clknet_leaf_315_clk _01433_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_215_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24847_ C_out\[250\] net98 net78 ser_C.shift_reg\[250\] _10893_ VGND VGND VPWR VPWR
+ _02500_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_215_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14600_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[15\]\[11\]
+ VGND VGND VPWR VPWR _11767_ sky130_fd_sc_hd__or2_1
XFILLER_160_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15580_ _12611_ _12636_ VGND VGND VPWR VPWR _12637_ sky130_fd_sc_hd__xnor2_1
X_27566_ clknet_leaf_299_clk _01364_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24778_ net113 ser_C.shift_reg\[217\] VGND VGND VPWR VPWR _10859_ sky130_fd_sc_hd__and2_1
XFILLER_233_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29305_ clknet_leaf_325_clk _03103_ net142 VGND VGND VPWR VPWR C_out\[277\] sky130_fd_sc_hd__dfrtp_1
XFILLER_96_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14531_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[15\]\[1\]
+ VGND VGND VPWR VPWR _11708_ sky130_fd_sc_hd__nand2_1
XFILLER_57_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26517_ clknet_leaf_11_A_in_serial_clk _00320_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_23729_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[0\]\[6\]
+ VGND VGND VPWR VPWR _10340_ sky130_fd_sc_hd__nand2_1
XFILLER_18_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27497_ clknet_leaf_226_clk _01295_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29236_ clknet_leaf_182_clk _03034_ net148 VGND VGND VPWR VPWR C_out\[208\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17250_ _04505_ _04508_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26448_ clknet_leaf_347_clk _00255_ net132 VGND VGND VPWR VPWR A_in\[116\] sky130_fd_sc_hd__dfrtp_1
X_14462_ _11641_ _11642_ VGND VGND VPWR VPWR _11644_ sky130_fd_sc_hd__and2_1
XFILLER_105_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16201_ _03582_ _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__nor2_1
X_13413_ A_in\[122\] deser_A.word_buffer\[122\] _00003_ VGND VGND VPWR VPWR _00261_
+ sky130_fd_sc_hd__mux2_1
X_29167_ clknet_leaf_39_clk _02965_ net141 VGND VGND VPWR VPWR C_out\[139\] sky130_fd_sc_hd__dfrtp_1
X_17181_ systolic_inst.A_outs\[10\]\[3\] systolic_inst.A_outs\[9\]\[3\] net120 VGND
+ VGND VPWR VPWR _01269_ sky130_fd_sc_hd__mux2_1
XFILLER_224_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14393_ _11575_ _11576_ VGND VGND VPWR VPWR _11577_ sky130_fd_sc_hd__nand2_1
X_26379_ clknet_leaf_22_clk _00186_ net133 VGND VGND VPWR VPWR A_in\[47\] sky130_fd_sc_hd__dfrtp_1
XFILLER_167_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28118_ clknet_leaf_128_clk _01916_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16132_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[7\]
+ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_42_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13344_ A_in\[53\] deser_A.word_buffer\[53\] net92 VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__mux2_1
X_29098_ clknet_leaf_154_clk _02896_ net150 VGND VGND VPWR VPWR C_out\[70\] sky130_fd_sc_hd__dfrtp_1
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28049_ clknet_leaf_130_clk _01847_ net144 VGND VGND VPWR VPWR systolic_inst.A_outs\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_16063_ _13055_ _13058_ VGND VGND VPWR VPWR _13059_ sky130_fd_sc_hd__xor2_1
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13275_ deser_A.word_buffer\[113\] deser_A.serial_word\[113\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__mux2_1
X_15014_ _12132_ _12133_ VGND VGND VPWR VPWR _12134_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_184_Right_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_244_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_244_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_97_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_204_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19822_ _06783_ _06821_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__nor2_1
XFILLER_116_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_204_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19753_ _06753_ _06754_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__or2_1
X_16965_ _04277_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_200_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15916_ _12936_ _12938_ _12941_ VGND VGND VPWR VPWR _12942_ sky130_fd_sc_hd__a21oi_2
X_18704_ _05792_ _05797_ _05828_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__o21ai_1
X_19684_ _06686_ _06687_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__or2_1
XFILLER_237_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16896_ _04200_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__xnor2_1
XFILLER_225_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18635_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[9\] _05761_
+ _05762_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_192_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[13\]\[13\]
+ _12877_ VGND VGND VPWR VPWR _12883_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18566_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[7\]
+ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__o21ai_2
XFILLER_80_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15778_ _12820_ _12821_ _12822_ VGND VGND VPWR VPWR _12824_ sky130_fd_sc_hd__and3_1
XFILLER_79_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17517_ _04768_ _04769_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14729_ _11866_ _11869_ _11873_ _11876_ VGND VGND VPWR VPWR _11877_ sky130_fd_sc_hd__o31a_1
X_18497_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[5\]
+ systolic_inst.A_outs\[8\]\[6\] VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__and4_1
XFILLER_162_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17448_ _04632_ _04635_ _04666_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__o21ai_1
XFILLER_221_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17379_ _04633_ _04634_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__and2b_1
XFILLER_186_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19118_ _06178_ _06179_ _06183_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__a21o_1
XFILLER_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20390_ _07320_ _07326_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19049_ _06117_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__and2_1
XFILLER_238_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22060_ _08831_ _08832_ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__or2_1
XFILLER_126_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_145_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21011_ systolic_inst.B_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[5\] systolic_inst.A_outs\[4\]\[7\]
+ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_235_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_235_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_173_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25750_ systolic_inst.acc_wires\[7\]\[2\] C_out\[226\] net40 VGND VGND VPWR VPWR
+ _03052_ sky130_fd_sc_hd__mux2_1
XFILLER_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22962_ _09638_ _09639_ VGND VGND VPWR VPWR _09640_ sky130_fd_sc_hd__nand2_1
XFILLER_68_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24701_ C_out\[177\] net100 net80 ser_C.shift_reg\[177\] _10820_ VGND VGND VPWR VPWR
+ _02427_ sky130_fd_sc_hd__a221o_1
XFILLER_215_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21913_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[3\]\[7\]
+ VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__or2_1
X_25681_ systolic_inst.acc_wires\[4\]\[29\] C_out\[157\] net32 VGND VGND VPWR VPWR
+ _02983_ sky130_fd_sc_hd__mux2_1
X_22893_ _09556_ _09572_ VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__or2_1
XFILLER_43_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27420_ clknet_leaf_248_clk _01218_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24632_ net7 ser_C.shift_reg\[144\] VGND VGND VPWR VPWR _10786_ sky130_fd_sc_hd__and2_1
X_21844_ _08620_ _08623_ _08645_ VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__and3_1
XFILLER_97_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27351_ clknet_leaf_233_clk _01149_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_24_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24563_ C_out\[108\] net100 net80 ser_C.shift_reg\[108\] _10751_ VGND VGND VPWR VPWR
+ _02358_ sky130_fd_sc_hd__a221o_1
XFILLER_196_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21775_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[11\] VGND
+ VGND VPWR VPWR _08581_ sky130_fd_sc_hd__and2_1
XFILLER_145_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26302_ clknet_leaf_24_A_in_serial_clk _00110_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_180_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20726_ _07624_ _07630_ _07638_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__a21o_1
XFILLER_168_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23514_ _10094_ _10096_ _10136_ _10137_ VGND VGND VPWR VPWR _10138_ sky130_fd_sc_hd__o211a_1
XFILLER_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27282_ clknet_leaf_323_clk _01080_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_24494_ net113 ser_C.shift_reg\[75\] VGND VGND VPWR VPWR _10717_ sky130_fd_sc_hd__and2_1
XFILLER_180_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29021_ clknet_leaf_93_clk _02819_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_26233_ clknet_leaf_10_A_in_serial_clk _00041_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23445_ _10068_ _10069_ VGND VGND VPWR VPWR _10070_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_134_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20657_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[5\]\[6\]
+ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_134_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23376_ systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[5\]
+ systolic_inst.B_outs\[0\]\[1\] VGND VGND VPWR VPWR _10003_ sky130_fd_sc_hd__a22oi_1
X_26164_ deser_B.serial_word\[119\] deser_B.shift_reg\[119\] net56 VGND VGND VPWR
+ VPWR _03466_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20588_ net120 _07517_ _07519_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_12_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25115_ C_out\[384\] net101 net73 ser_C.shift_reg\[384\] _11027_ VGND VGND VPWR VPWR
+ _02634_ sky130_fd_sc_hd__a221o_1
X_22327_ _09067_ _09068_ VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26095_ deser_B.serial_word\[50\] deser_B.shift_reg\[50\] net55 VGND VGND VPWR VPWR
+ _03397_ sky130_fd_sc_hd__mux2_1
XFILLER_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22258_ _08994_ _09002_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__nand2_1
XFILLER_152_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25046_ net113 ser_C.shift_reg\[351\] VGND VGND VPWR VPWR _10993_ sky130_fd_sc_hd__and2_1
XFILLER_180_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_240_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_240_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21209_ _08075_ _08076_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_226_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_226_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_240_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22189_ _08933_ _08934_ _08922_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__o21bai_1
XFILLER_239_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28805_ clknet_leaf_247_clk _02603_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[353\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26997_ clknet_leaf_18_B_in_serial_clk _00795_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28736_ clknet_leaf_301_clk _02534_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16750_ _04067_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__xnor2_1
X_25948_ systolic_inst.acc_wires\[13\]\[8\] C_out\[424\] net19 VGND VGND VPWR VPWR
+ _03250_ sky130_fd_sc_hd__mux2_1
X_13962_ deser_A.serial_word\[123\] deser_A.shift_reg\[123\] _00002_ VGND VGND VPWR
+ VPWR _00788_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_21_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15701_ _12687_ _12753_ VGND VGND VPWR VPWR _12754_ sky130_fd_sc_hd__nand2_1
X_28667_ clknet_leaf_187_clk _02465_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[215\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16681_ _03997_ _03998_ _04002_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_238_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25879_ systolic_inst.acc_wires\[11\]\[3\] C_out\[355\] net38 VGND VGND VPWR VPWR
+ _03181_ sky130_fd_sc_hd__mux2_1
X_13893_ deser_A.serial_word\[54\] deser_A.shift_reg\[54\] net58 VGND VGND VPWR VPWR
+ _00719_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_238_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18420_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[0\] _05556_
+ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__a21o_1
XFILLER_235_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15632_ _12616_ _12686_ VGND VGND VPWR VPWR _12687_ sky130_fd_sc_hd__xnor2_4
X_27618_ clknet_leaf_318_clk _01416_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_28598_ clknet_leaf_138_clk _02396_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18351_ net66 _05511_ _05512_ systolic_inst.acc_wires\[9\]\[23\] net106 VGND VGND
+ VPWR VPWR _01385_ sky130_fd_sc_hd__a32o_1
XFILLER_15_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15563_ _12616_ _12619_ VGND VGND VPWR VPWR _12620_ sky130_fd_sc_hd__xnor2_1
X_27549_ clknet_leaf_300_clk _01347_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17302_ net118 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[6\] VGND
+ VGND VPWR VPWR _04561_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_44_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _11690_ _11691_ VGND VGND VPWR VPWR _11694_ sky130_fd_sc_hd__and2_1
XFILLER_70_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _05441_ _05444_ _05448_ _05452_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__a211o_1
X_15494_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[7\] VGND VGND
+ VPWR VPWR _12553_ sky130_fd_sc_hd__and2b_1
XFILLER_124_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29219_ clknet_leaf_183_clk _03017_ net146 VGND VGND VPWR VPWR C_out\[191\] sky130_fd_sc_hd__dfrtp_1
X_17233_ _04477_ _04493_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__nor2_1
X_14445_ _11625_ _11626_ VGND VGND VPWR VPWR _11627_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17164_ _04445_ _04447_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14376_ _11447_ _11559_ VGND VGND VPWR VPWR _11560_ sky130_fd_sc_hd__xor2_1
XFILLER_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_185_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16115_ _13072_ _03498_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__xor2_1
XFILLER_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13327_ A_in\[36\] deser_A.word_buffer\[36\] net94 VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__mux2_1
XFILLER_171_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17095_ _04387_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__xor2_1
XFILLER_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16046_ _13034_ _13042_ VGND VGND VPWR VPWR _13043_ sky130_fd_sc_hd__nor2_1
X_13258_ deser_A.word_buffer\[96\] deser_A.serial_word\[96\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__mux2_1
XFILLER_170_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_217_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_217_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_170_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13189_ deser_A.word_buffer\[27\] deser_A.serial_word\[27\] net128 VGND VGND VPWR
+ VPWR _00037_ sky130_fd_sc_hd__mux2_1
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19805_ _06787_ _06804_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__xor2_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17997_ _05150_ _05187_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_140_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19736_ _06710_ _06736_ _06737_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__nor3_1
X_16948_ _04199_ _04262_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__xnor2_1
XFILLER_238_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19667_ _06651_ _06671_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__xnor2_1
X_16879_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[7\] _04167_ _04132_
+ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__a31o_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18618_ _05745_ _05744_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__nand2b_1
X_19598_ _06623_ _06625_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18549_ _05641_ _05677_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_174_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21560_ _08370_ _08369_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__nand2b_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20511_ _07435_ _07443_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_220_Right_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21491_ _08298_ _08305_ VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_170_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23230_ _09858_ _09878_ VGND VGND VPWR VPWR _09879_ sky130_fd_sc_hd__nor2_1
XFILLER_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20442_ _07332_ _07341_ _07340_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__o21ba_1
X_23161_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[1\]\[14\]
+ VGND VGND VPWR VPWR _09820_ sky130_fd_sc_hd__or2_1
XFILLER_140_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20373_ _07307_ _07308_ _07309_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__a21oi_1
Xclkload340 clknet_leaf_0_A_in_serial_clk VGND VGND VPWR VPWR clkload340/Y sky130_fd_sc_hd__clkinv_2
XFILLER_88_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload351 clknet_leaf_26_A_in_serial_clk VGND VGND VPWR VPWR clkload351/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_238_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload362 clknet_leaf_14_A_in_serial_clk VGND VGND VPWR VPWR clkload362/Y sky130_fd_sc_hd__bufinv_16
X_22112_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[2\]
+ systolic_inst.A_outs\[2\]\[3\] VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__nand4_2
Xclkload70 clknet_leaf_347_clk VGND VGND VPWR VPWR clkload70/Y sky130_fd_sc_hd__inv_6
XFILLER_106_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload373 clknet_leaf_27_B_in_serial_clk VGND VGND VPWR VPWR clkload373/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23092_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[1\]\[4\]
+ VGND VGND VPWR VPWR _09761_ sky130_fd_sc_hd__nand2_1
Xclkload384 clknet_leaf_4_B_in_serial_clk VGND VGND VPWR VPWR clkload384/Y sky130_fd_sc_hd__clkinv_4
Xclkload81 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload81/Y sky130_fd_sc_hd__inv_6
Xclkload395 clknet_leaf_17_B_in_serial_clk VGND VGND VPWR VPWR clkload395/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_8_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload92 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload92/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_168_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_208_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_208_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22043_ _08809_ _08811_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__and2_1
XFILLER_47_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26920_ clknet_leaf_4_A_in_serial_clk _00718_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26851_ clknet_leaf_67_clk _00653_ net134 VGND VGND VPWR VPWR B_in\[123\] sky130_fd_sc_hd__dfrtp_1
XFILLER_141_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25802_ systolic_inst.acc_wires\[8\]\[22\] C_out\[278\] net28 VGND VGND VPWR VPWR
+ _03104_ sky130_fd_sc_hd__mux2_1
XFILLER_60_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29570_ clknet_leaf_21_B_in_serial_clk _03365_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26782_ clknet_leaf_56_clk _00584_ net143 VGND VGND VPWR VPWR B_in\[54\] sky130_fd_sc_hd__dfrtp_1
X_23994_ _10522_ systolic_inst.B_shift\[5\]\[0\] _11332_ VGND VGND VPWR VPWR _02018_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28521_ clknet_leaf_154_clk _02319_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25733_ systolic_inst.acc_wires\[6\]\[17\] C_out\[209\] net46 VGND VGND VPWR VPWR
+ _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_112_1355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_867 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22945_ _09515_ _09621_ VGND VGND VPWR VPWR _09623_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28452_ clknet_leaf_131_clk _02250_ net144 VGND VGND VPWR VPWR ser_C.shift_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_112_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25664_ systolic_inst.acc_wires\[4\]\[12\] C_out\[140\] net30 VGND VGND VPWR VPWR
+ _02966_ sky130_fd_sc_hd__mux2_1
XFILLER_44_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22876_ _09554_ _09555_ VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__or2_1
XFILLER_83_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27403_ clknet_leaf_333_clk _01201_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24615_ C_out\[134\] net103 net75 ser_C.shift_reg\[134\] _10777_ VGND VGND VPWR VPWR
+ _02384_ sky130_fd_sc_hd__a221o_1
X_21827_ _08630_ _08629_ VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__and2b_1
XFILLER_169_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28383_ clknet_leaf_31_clk _02181_ VGND VGND VPWR VPWR systolic_inst.A_shift\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_233_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25595_ systolic_inst.acc_wires\[2\]\[7\] C_out\[71\] net34 VGND VGND VPWR VPWR _02897_
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27334_ clknet_leaf_286_clk _01132_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_24546_ net113 ser_C.shift_reg\[101\] VGND VGND VPWR VPWR _10743_ sky130_fd_sc_hd__and2_1
XFILLER_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21758_ _08561_ _08562_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20709_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[5\]\[12\]
+ _07621_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__and3_1
X_27265_ clknet_leaf_282_clk _01063_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_71_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24477_ C_out\[65\] _11302_ net81 ser_C.shift_reg\[65\] _10708_ VGND VGND VPWR VPWR
+ _02315_ sky130_fd_sc_hd__a221o_1
XFILLER_196_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21689_ _08494_ _08495_ VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__xnor2_1
X_29004_ clknet_leaf_104_clk _02802_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14230_ _11415_ _11417_ VGND VGND VPWR VPWR _11418_ sky130_fd_sc_hd__nor2_1
X_26216_ clknet_leaf_12_A_in_serial_clk _00024_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_23428_ _10010_ _10012_ _10052_ _10053_ VGND VGND VPWR VPWR _10054_ sky130_fd_sc_hd__o211a_2
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27196_ clknet_leaf_259_clk _00994_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_153_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_242_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26147_ deser_B.serial_word\[102\] deser_B.shift_reg\[102\] _00001_ VGND VGND VPWR
+ VPWR _03449_ sky130_fd_sc_hd__mux2_1
XFILLER_125_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14161_ _11350_ _11351_ VGND VGND VPWR VPWR _11352_ sky130_fd_sc_hd__or2_1
X_23359_ _09965_ _09985_ VGND VGND VPWR VPWR _09987_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_242_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_242_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13112_ systolic_inst.A_outs\[0\]\[5\] VGND VGND VPWR VPWR _11268_ sky130_fd_sc_hd__inv_2
X_26078_ deser_B.serial_word\[33\] deser_B.shift_reg\[33\] net55 VGND VGND VPWR VPWR
+ _03380_ sky130_fd_sc_hd__mux2_1
X_14092_ deser_B.shift_reg\[126\] deser_B.shift_reg\[127\] net126 VGND VGND VPWR VPWR
+ _00918_ sky130_fd_sc_hd__mux2_1
XFILLER_153_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_180_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xload_slew107 net109 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_16
X_25029_ C_out\[341\] net97 net77 ser_C.shift_reg\[341\] _10984_ VGND VGND VPWR VPWR
+ _02591_ sky130_fd_sc_hd__a221o_1
X_17920_ _11263_ _05113_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17851_ _05027_ _05044_ _05046_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__and3_1
XFILLER_67_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16802_ _04081_ _04083_ _04120_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__and3_1
X_17782_ _04994_ _04998_ _04999_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__a21oi_1
XFILLER_226_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14994_ systolic_inst.A_outs\[14\]\[4\] systolic_inst.B_outs\[14\]\[6\] _11264_ systolic_inst.A_outs\[14\]\[3\]
+ VGND VGND VPWR VPWR _12114_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_66_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19521_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[16\]
+ _06557_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__a21oi_1
X_16733_ systolic_inst.B_outs\[11\]\[7\] _04020_ _04021_ VGND VGND VPWR VPWR _04054_
+ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_178_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13945_ deser_A.serial_word\[106\] deser_A.shift_reg\[106\] net57 VGND VGND VPWR
+ VPWR _00771_ sky130_fd_sc_hd__mux2_1
X_28719_ clknet_leaf_310_clk _02517_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_178_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19452_ _06497_ _06500_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__and2_1
XFILLER_90_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16664_ systolic_inst.A_outs\[11\]\[4\] _03950_ _03968_ _03967_ _03964_ VGND VGND
+ VPWR VPWR _03987_ sky130_fd_sc_hd__a32o_1
XFILLER_234_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13876_ deser_A.serial_word\[37\] deser_A.shift_reg\[37\] net58 VGND VGND VPWR VPWR
+ _00702_ sky130_fd_sc_hd__mux2_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15615_ _12611_ _12636_ _12635_ VGND VGND VPWR VPWR _12671_ sky130_fd_sc_hd__a21boi_1
X_18403_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.A_shift\[16\]\[0\] net121 VGND
+ VGND VPWR VPWR _01394_ sky130_fd_sc_hd__mux2_1
X_19383_ _06441_ _06440_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__and2b_1
XFILLER_37_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16595_ net118 _03922_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__nand2_1
XFILLER_203_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18334_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[21\]
+ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__xnor2_2
XFILLER_43_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15546_ _12565_ _12567_ VGND VGND VPWR VPWR _12604_ sky130_fd_sc_hd__and2_1
XFILLER_15_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18265_ _05438_ _05437_ systolic_inst.acc_wires\[9\]\[11\] net107 VGND VGND VPWR
+ VPWR _01373_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_175_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15477_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[6\] _12536_ net116
+ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__mux2_1
XFILLER_204_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17216_ systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[3\]
+ systolic_inst.B_outs\[10\]\[0\] VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__a22o_1
X_14428_ _11608_ _11609_ VGND VGND VPWR VPWR _11611_ sky130_fd_sc_hd__xnor2_1
X_18196_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[9\]\[1\]
+ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__or2_1
XFILLER_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17147_ _04431_ _04433_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14359_ _11514_ _11543_ VGND VGND VPWR VPWR _11544_ sky130_fd_sc_hd__nand2_1
XFILLER_155_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17078_ _04362_ _04369_ _04370_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__o21ba_1
XFILLER_171_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16029_ _12991_ _13012_ _13014_ VGND VGND VPWR VPWR _13026_ sky130_fd_sc_hd__a21oi_1
XFILLER_100_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19719_ systolic_inst.B_outs\[6\]\[3\] systolic_inst.A_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\]
+ systolic_inst.A_outs\[6\]\[2\] VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__a22oi_1
Xclkbuf_5_4__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_38_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20991_ _07862_ _07863_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22730_ _09393_ _09411_ _09412_ VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__or3_1
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22661_ systolic_inst.acc_wires\[2\]\[28\] systolic_inst.acc_wires\[2\]\[29\] systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__o21ai_1
XFILLER_168_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24400_ net114 ser_C.shift_reg\[28\] VGND VGND VPWR VPWR _10670_ sky130_fd_sc_hd__and2_1
X_21612_ _08418_ _08421_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25380_ _11159_ systolic_inst.B_shift\[14\]\[5\] net70 VGND VGND VPWR VPWR _02767_
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22592_ _09301_ _09303_ _09310_ VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__a21oi_1
XFILLER_200_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24331_ systolic_inst.A_shift\[10\]\[5\] A_in\[37\] net59 VGND VGND VPWR VPWR _10639_
+ sky130_fd_sc_hd__mux2_1
X_21543_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[3\] VGND VGND VPWR
+ VPWR _08355_ sky130_fd_sc_hd__nand2_1
X_27050_ clknet_leaf_24_B_in_serial_clk _00848_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_21474_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.B_shift\[2\]\[2\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__mux2_1
X_24262_ systolic_inst.A_shift\[16\]\[5\] net70 net83 systolic_inst.A_shift\[17\]\[5\]
+ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26001_ systolic_inst.acc_wires\[14\]\[29\] ser_C.parallel_data\[477\] net24 VGND
+ VGND VPWR VPWR _03303_ sky130_fd_sc_hd__mux2_1
X_23213_ _09864_ _09863_ systolic_inst.acc_wires\[1\]\[21\] net109 VGND VGND VPWR
+ VPWR _01895_ sky130_fd_sc_hd__a2bb2o_1
X_20425_ _07322_ _07360_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__nor2_1
XFILLER_140_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1034 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24193_ systolic_inst.B_shift\[22\]\[0\] net72 _11333_ B_in\[112\] VGND VGND VPWR
+ VPWR _02154_ sky130_fd_sc_hd__a22o_1
XFILLER_88_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23144_ net109 systolic_inst.acc_wires\[1\]\[11\] net64 _09805_ VGND VGND VPWR VPWR
+ _01885_ sky130_fd_sc_hd__a22o_1
X_20356_ _07257_ _07292_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__xnor2_1
Xclkload170 clknet_leaf_243_clk VGND VGND VPWR VPWR clkload170/Y sky130_fd_sc_hd__clkinv_2
XFILLER_101_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload181 clknet_leaf_237_clk VGND VGND VPWR VPWR clkload181/Y sky130_fd_sc_hd__bufinv_16
Xclkload192 clknet_leaf_64_clk VGND VGND VPWR VPWR clkload192/Y sky130_fd_sc_hd__inv_6
X_23075_ _09746_ VGND VGND VPWR VPWR _09747_ sky130_fd_sc_hd__inv_2
X_27952_ clknet_leaf_171_clk _01750_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20287_ _07227_ _07226_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[4\]
+ net109 VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_73_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22026_ _08784_ _08791_ _08796_ _08800_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__and4_1
X_26903_ clknet_leaf_16_A_in_serial_clk _00701_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_222_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27883_ clknet_leaf_45_clk _01681_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_49_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26834_ clknet_leaf_89_clk _00636_ net5 VGND VGND VPWR VPWR B_in\[106\] sky130_fd_sc_hd__dfrtp_1
X_29622_ clknet_leaf_8_B_in_serial_clk _03417_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29553_ clknet_leaf_3_B_in_serial_clk _03348_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26765_ clknet_leaf_80_clk _00567_ net153 VGND VGND VPWR VPWR B_in\[37\] sky130_fd_sc_hd__dfrtp_1
XFILLER_151_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_235_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23977_ systolic_inst.B_shift\[12\]\[0\] B_in\[64\] _00008_ VGND VGND VPWR VPWR _10514_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_235_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28504_ clknet_leaf_114_clk _02302_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_13730_ B_in\[37\] deser_B.word_buffer\[37\] net90 VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__mux2_1
X_25716_ systolic_inst.acc_wires\[6\]\[0\] C_out\[192\] net47 VGND VGND VPWR VPWR
+ _03018_ sky130_fd_sc_hd__mux2_1
XFILLER_17_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22928_ _09588_ _09606_ VGND VGND VPWR VPWR _09607_ sky130_fd_sc_hd__xor2_1
X_29484_ clknet_leaf_281_clk _03282_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[456\]
+ sky130_fd_sc_hd__dfrtp_1
X_26696_ clknet_leaf_5_B_in_serial_clk _00499_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_231_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_231_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28435_ clknet_leaf_28_clk _02233_ VGND VGND VPWR VPWR systolic_inst.A_shift\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_231_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25647_ systolic_inst.acc_wires\[3\]\[27\] C_out\[123\] net50 VGND VGND VPWR VPWR
+ _02949_ sky130_fd_sc_hd__mux2_1
X_13661_ deser_B.word_buffer\[97\] deser_B.serial_word\[97\] net123 VGND VGND VPWR
+ VPWR _00498_ sky130_fd_sc_hd__mux2_1
X_22859_ _09464_ _09498_ _09500_ VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15400_ net107 _12460_ _12461_ _12462_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__o31ai_1
XFILLER_25_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16380_ _03754_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__inv_2
X_28366_ clknet_leaf_29_clk _02164_ VGND VGND VPWR VPWR systolic_inst.A_shift\[20\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25578_ systolic_inst.acc_wires\[1\]\[22\] C_out\[54\] net53 VGND VGND VPWR VPWR
+ _02880_ sky130_fd_sc_hd__mux2_1
XFILLER_213_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13592_ deser_B.word_buffer\[28\] deser_B.serial_word\[28\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__mux2_1
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27317_ clknet_leaf_289_clk _01115_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15331_ _12410_ _12414_ VGND VGND VPWR VPWR _12417_ sky130_fd_sc_hd__nor2_1
XFILLER_34_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24529_ C_out\[91\] net100 net82 ser_C.shift_reg\[91\] _10734_ VGND VGND VPWR VPWR
+ _02341_ sky130_fd_sc_hd__a221o_1
XFILLER_185_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28297_ clknet_leaf_123_clk _02095_ VGND VGND VPWR VPWR systolic_inst.B_shift\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18050_ _05222_ _05240_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__xor2_1
X_15262_ net107 systolic_inst.acc_wires\[14\]\[16\] _12357_ _12359_ VGND VGND VPWR
+ VPWR _01058_ sky130_fd_sc_hd__a22o_1
X_27248_ clknet_leaf_271_clk _01046_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_229_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17001_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[11\]\[5\]
+ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_229_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14213_ _11373_ _11375_ _11400_ net107 VGND VGND VPWR VPWR _11402_ sky130_fd_sc_hd__a31o_1
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15193_ _12298_ _12299_ _12292_ _12296_ VGND VGND VPWR VPWR _12300_ sky130_fd_sc_hd__a211o_1
X_27179_ clknet_leaf_248_clk _00977_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_7 systolic_inst.A_outs\[3\]\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14144_ net107 _11336_ VGND VGND VPWR VPWR _11337_ sky130_fd_sc_hd__nor2_1
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14075_ deser_B.shift_reg\[109\] deser_B.shift_reg\[110\] deser_B.receiving VGND
+ VGND VPWR VPWR _00901_ sky130_fd_sc_hd__mux2_1
X_18952_ _06042_ _06043_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__nor2_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17903_ _05065_ _05097_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__xnor2_1
X_18883_ _05984_ _05987_ _05990_ net61 VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__a31o_1
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17834_ systolic_inst.A_outs\[9\]\[1\] systolic_inst.B_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\]
+ systolic_inst.A_outs\[9\]\[0\] VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__a22o_1
XFILLER_79_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14977_ _12097_ VGND VGND VPWR VPWR _12098_ sky130_fd_sc_hd__inv_2
X_17765_ _04984_ _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__nand2_1
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19504_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[15\]
+ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__nor2_1
X_13928_ deser_A.serial_word\[89\] deser_A.shift_reg\[89\] net57 VGND VGND VPWR VPWR
+ _00754_ sky130_fd_sc_hd__mux2_1
X_16716_ _04031_ _04037_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__nor2_1
X_17696_ net106 systolic_inst.acc_wires\[10\]\[17\] net68 _04927_ VGND VGND VPWR VPWR
+ _01315_ sky130_fd_sc_hd__a22o_1
XFILLER_212_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19435_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[7\]\[5\]
+ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__or2_1
X_16647_ systolic_inst.A_outs\[11\]\[2\] systolic_inst.B_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\]
+ systolic_inst.A_outs\[11\]\[1\] VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__a22oi_1
X_13859_ deser_A.serial_word\[20\] deser_A.shift_reg\[20\] net58 VGND VGND VPWR VPWR
+ _00685_ sky130_fd_sc_hd__mux2_1
XFILLER_222_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19366_ _06391_ _06393_ _06424_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__o21a_1
X_16578_ systolic_inst.A_outs\[11\]\[3\] systolic_inst.A_outs\[10\]\[3\] net118 VGND
+ VGND VPWR VPWR _01205_ sky130_fd_sc_hd__mux2_1
XFILLER_222_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18317_ _05482_ _05483_ _05481_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__a21o_1
XFILLER_31_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15529_ systolic_inst.A_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[5\] VGND VGND
+ VPWR VPWR _12587_ sky130_fd_sc_hd__nand2_1
X_19297_ _06319_ _06321_ _06358_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__a21o_1
XFILLER_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18248_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[9\]\[9\]
+ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__nand2_1
XFILLER_124_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18179_ _05317_ _05343_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__and2_1
XFILLER_239_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20210_ net106 systolic_inst.acc_wires\[6\]\[29\] net68 _07173_ VGND VGND VPWR VPWR
+ _01583_ sky130_fd_sc_hd__a22o_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21190_ _08057_ _08058_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__nor2_1
XFILLER_85_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20141_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[19\]
+ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20072_ _07051_ _07053_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__nand2_1
XFILLER_98_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23900_ systolic_inst.B_shift\[17\]\[2\] B_in\[74\] _00008_ VGND VGND VPWR VPWR _10483_
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24880_ net110 ser_C.shift_reg\[268\] VGND VGND VPWR VPWR _10910_ sky130_fd_sc_hd__and2_1
XFILLER_100_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23831_ _10425_ _10426_ VGND VGND VPWR VPWR _10427_ sky130_fd_sc_hd__xor2_1
XFILLER_61_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26550_ clknet_leaf_19_A_in_serial_clk _00353_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_226_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23762_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[0\]\[11\]
+ VGND VGND VPWR VPWR _10368_ sky130_fd_sc_hd__or2_1
XFILLER_214_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20974_ _07844_ _07847_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__xor2_1
XFILLER_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25501_ _11228_ _11230_ systolic_inst.cycle_cnt\[23\] VGND VGND VPWR VPWR _02817_
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22713_ _09392_ _09397_ VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26481_ clknet_leaf_13_A_in_serial_clk _00284_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23693_ net121 _10308_ _10309_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__a21oi_1
XFILLER_213_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28220_ clknet_leaf_99_clk _02018_ VGND VGND VPWR VPWR systolic_inst.B_shift\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25432_ _11185_ systolic_inst.A_shift\[0\]\[7\] net70 VGND VGND VPWR VPWR _02793_
+ sky130_fd_sc_hd__mux2_1
X_22644_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[27\]
+ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__xnor2_1
XFILLER_213_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28151_ clknet_leaf_102_clk _01949_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25363_ ser_C.parallel_data\[508\] net98 net78 ser_C.shift_reg\[508\] _11151_ VGND
+ VGND VPWR VPWR _02758_ sky130_fd_sc_hd__a221o_1
X_22575_ _09281_ _09287_ _09295_ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_118_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27102_ clknet_leaf_9_B_in_serial_clk _00900_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24314_ _10630_ systolic_inst.A_shift\[10\]\[4\] net70 VGND VGND VPWR VPWR _02230_
+ sky130_fd_sc_hd__mux2_1
X_28082_ clknet_leaf_115_clk _01880_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_21526_ _08338_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25294_ net111 ser_C.shift_reg\[475\] VGND VGND VPWR VPWR _11117_ sky130_fd_sc_hd__and2_1
XFILLER_194_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27033_ clknet_leaf_13_B_in_serial_clk _00831_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_182_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24245_ systolic_inst.A_shift\[19\]\[6\] A_in\[70\] net59 VGND VGND VPWR VPWR _10608_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21457_ _08288_ _08291_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20408_ _07342_ _07343_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_224_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21388_ _08231_ _08232_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__and2_1
X_24176_ systolic_inst.A_shift\[26\]\[7\] net70 _10505_ systolic_inst.A_shift\[27\]\[7\]
+ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__a22o_1
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR C_out_serial_data sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_224_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23127_ _09786_ _09788_ VGND VGND VPWR VPWR _09791_ sky130_fd_sc_hd__nand2_1
X_20339_ _07275_ _07276_ _07244_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__a21o_1
XFILLER_150_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28984_ clknet_leaf_58_clk _02782_ VGND VGND VPWR VPWR systolic_inst.A_shift\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27935_ clknet_leaf_180_clk _01733_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_23058_ _09731_ _09732_ VGND VGND VPWR VPWR _09733_ sky130_fd_sc_hd__or2_1
XFILLER_110_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14900_ _11990_ _12022_ VGND VGND VPWR VPWR _12023_ sky130_fd_sc_hd__nand2b_1
X_22009_ net65 _08788_ _08789_ systolic_inst.acc_wires\[3\]\[20\] net106 VGND VGND
+ VPWR VPWR _01766_ sky130_fd_sc_hd__a32o_1
XFILLER_153_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27866_ clknet_leaf_144_clk _01664_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15880_ _12909_ _12910_ VGND VGND VPWR VPWR _12911_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29605_ clknet_leaf_25_B_in_serial_clk _03400_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_14831_ _11933_ _11955_ VGND VGND VPWR VPWR _11956_ sky130_fd_sc_hd__nand2b_1
X_26817_ clknet_leaf_66_clk _00619_ net135 VGND VGND VPWR VPWR B_in\[89\] sky130_fd_sc_hd__dfrtp_1
XFILLER_48_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27797_ clknet_leaf_48_clk _01595_ net137 VGND VGND VPWR VPWR systolic_inst.B_outs\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17550_ _04799_ _04800_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__nand2_1
X_26748_ clknet_leaf_52_clk _00550_ net143 VGND VGND VPWR VPWR B_in\[20\] sky130_fd_sc_hd__dfrtp_1
X_14762_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[1\] _11888_
+ _11890_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__a22o_1
X_29536_ clknet_leaf_257_clk _03334_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[508\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16501_ _03851_ _03855_ _03857_ net61 VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__a31o_1
XFILLER_229_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13713_ B_in\[20\] deser_B.word_buffer\[20\] net86 VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__mux2_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29467_ clknet_leaf_287_clk _03265_ net136 VGND VGND VPWR VPWR C_out\[439\] sky130_fd_sc_hd__dfrtp_1
X_17481_ _04695_ _04697_ _04732_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__a21oi_1
XFILLER_189_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26679_ clknet_leaf_11_B_in_serial_clk _00482_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[81\]
+ sky130_fd_sc_hd__dfrtp_1
X_14693_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[24\]
+ VGND VGND VPWR VPWR _11847_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19220_ systolic_inst.A_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[6\] _11261_ systolic_inst.A_outs\[7\]\[2\]
+ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_28_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16432_ _03796_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__or2_1
XFILLER_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13644_ deser_B.word_buffer\[80\] deser_B.serial_word\[80\] net123 VGND VGND VPWR
+ VPWR _00481_ sky130_fd_sc_hd__mux2_1
X_28418_ clknet_leaf_70_clk _02216_ VGND VGND VPWR VPWR systolic_inst.B_shift\[23\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29398_ clknet_leaf_239_clk _03196_ net145 VGND VGND VPWR VPWR C_out\[370\] sky130_fd_sc_hd__dfrtp_1
XFILLER_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19151_ _06213_ _06216_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16363_ net108 _03730_ _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__or3_1
X_28349_ clknet_leaf_319_clk _02147_ VGND VGND VPWR VPWR systolic_inst.A_shift\[24\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13575_ deser_B.word_buffer\[11\] deser_B.serial_word\[11\] net124 VGND VGND VPWR
+ VPWR _00412_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18102_ _05289_ _05290_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__nand2_1
X_15314_ _12397_ _12399_ _12402_ net61 VGND VGND VPWR VPWR _12404_ sky130_fd_sc_hd__a31o_1
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19082_ _06132_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__xor2_1
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16294_ _03629_ _03645_ _03643_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__o21a_1
XFILLER_160_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18033_ systolic_inst.B_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[7\]
+ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__and3_1
X_15245_ _12342_ _12344_ VGND VGND VPWR VPWR _12345_ sky130_fd_sc_hd__nand2_1
XFILLER_160_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15176_ _11712_ _12283_ _12285_ systolic_inst.acc_wires\[14\]\[4\] net107 VGND VGND
+ VPWR VPWR _01046_ sky130_fd_sc_hd__a32o_1
XFILLER_158_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14127_ systolic_inst.A_outs\[15\]\[3\] systolic_inst.A_outs\[14\]\[3\] net118 VGND
+ VGND VPWR VPWR _00949_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19984_ _11278_ systolic_inst.A_outs\[6\]\[7\] _06928_ _06951_ VGND VGND VPWR VPWR
+ _06979_ sky130_fd_sc_hd__o211a_1
XFILLER_141_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14058_ deser_B.shift_reg\[92\] deser_B.shift_reg\[93\] net126 VGND VGND VPWR VPWR
+ _00884_ sky130_fd_sc_hd__mux2_1
X_18935_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[20\]
+ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_207_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18866_ net63 _05975_ _05976_ systolic_inst.acc_wires\[8\]\[10\] net108 VGND VGND
+ VPWR VPWR _01436_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_199_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17817_ systolic_inst.A_outs\[9\]\[1\] systolic_inst.B_outs\[9\]\[2\] systolic_inst.B_outs\[9\]\[3\]
+ systolic_inst.A_outs\[9\]\[0\] VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__a22oi_1
XFILLER_67_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18797_ _05910_ _05911_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17748_ net69 _04970_ _04971_ systolic_inst.acc_wires\[10\]\[25\] net105 VGND VGND
+ VPWR VPWR _01323_ sky130_fd_sc_hd__a32o_1
XFILLER_223_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17679_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[15\]
+ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__and2_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19418_ net69 _06470_ _06472_ systolic_inst.acc_wires\[7\]\[2\] net105 VGND VGND
+ VPWR VPWR _01492_ sky130_fd_sc_hd__a32o_1
X_20690_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[5\]\[11\]
+ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__or2_1
XFILLER_161_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19349_ _06380_ _06408_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22360_ _09063_ _09065_ _09064_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_14_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_198_Right_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21311_ _08160_ _08163_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__nand2_1
X_22291_ _08995_ _08997_ _08996_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__o21ba_1
XFILLER_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24030_ _10532_ systolic_inst.B_shift\[4\]\[2\] net72 VGND VGND VPWR VPWR _02044_
+ sky130_fd_sc_hd__mux2_1
X_21242_ _08084_ _08106_ _08107_ _08108_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__nand4_1
XFILLER_11_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21173_ _08038_ _08041_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__nand2_1
XFILLER_105_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20124_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[16\]
+ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25981_ systolic_inst.acc_wires\[14\]\[9\] ser_C.parallel_data\[457\] net25 VGND
+ VGND VPWR VPWR _03283_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27720_ clknet_leaf_187_clk _01518_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_209_Left_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20055_ _07038_ _07039_ _07040_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__and3_1
X_24932_ net111 ser_C.shift_reg\[294\] VGND VGND VPWR VPWR _10936_ sky130_fd_sc_hd__and2_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_0_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27651_ clknet_leaf_313_clk _01449_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24863_ C_out\[258\] net101 net73 ser_C.shift_reg\[258\] _10901_ VGND VGND VPWR VPWR
+ _02508_ sky130_fd_sc_hd__a221o_1
XFILLER_6_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26602_ clknet_leaf_18_B_in_serial_clk _00405_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23814_ systolic_inst.acc_wires\[0\]\[16\] systolic_inst.acc_wires\[0\]\[17\] systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _10413_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_68_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27582_ clknet_leaf_219_clk _01380_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24794_ net112 ser_C.shift_reg\[225\] VGND VGND VPWR VPWR _10867_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29321_ clknet_leaf_298_clk _03119_ net138 VGND VGND VPWR VPWR C_out\[293\] sky130_fd_sc_hd__dfrtp_1
XFILLER_199_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26533_ clknet_leaf_17_A_in_serial_clk _00336_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23745_ _10351_ _10352_ net63 VGND VGND VPWR VPWR _10354_ sky130_fd_sc_hd__o21ai_1
XFILLER_96_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20957_ _07796_ _07799_ _07830_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__or3_1
XFILLER_199_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29252_ clknet_leaf_200_clk _03050_ net146 VGND VGND VPWR VPWR C_out\[224\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26464_ clknet_leaf_1_A_in_serial_clk _00271_ net132 VGND VGND VPWR VPWR deser_A.bit_idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_241_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23676_ _10269_ _10294_ VGND VGND VPWR VPWR _10295_ sky130_fd_sc_hd__nand2_1
XFILLER_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20888_ _07756_ _07764_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28203_ clknet_leaf_131_clk _02001_ VGND VGND VPWR VPWR systolic_inst.B_shift\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25415_ systolic_inst.A_shift\[2\]\[7\] A_in\[15\] net59 VGND VGND VPWR VPWR _11177_
+ sky130_fd_sc_hd__mux2_1
X_22627_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[24\]
+ VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_218_Left_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29183_ clknet_leaf_44_clk _02981_ net142 VGND VGND VPWR VPWR C_out\[155\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26395_ clknet_leaf_14_clk _00202_ net133 VGND VGND VPWR VPWR A_in\[63\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28134_ clknet_leaf_128_clk _01932_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25346_ net112 ser_C.shift_reg\[501\] VGND VGND VPWR VPWR _11143_ sky130_fd_sc_hd__and2_1
XFILLER_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13360_ A_in\[69\] deser_A.word_buffer\[69\] net96 VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__mux2_1
XFILLER_224_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22558_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[2\]\[12\]
+ _09278_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__and3_1
XFILLER_195_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28065_ clknet_leaf_120_clk _01863_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_21509_ _08320_ _08321_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13291_ A_in\[0\] deser_A.word_buffer\[0\] net93 VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__mux2_1
X_25277_ ser_C.parallel_data\[465\] net102 net74 ser_C.shift_reg\[465\] _11108_ VGND
+ VGND VPWR VPWR _02715_ sky130_fd_sc_hd__a221o_1
X_22489_ _09219_ _09220_ _09221_ VGND VGND VPWR VPWR _09223_ sky130_fd_sc_hd__and3_1
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27016_ clknet_leaf_22_B_in_serial_clk _00814_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15030_ systolic_inst.A_outs\[14\]\[5\] systolic_inst.B_outs\[14\]\[6\] _11264_ systolic_inst.A_outs\[14\]\[4\]
+ VGND VGND VPWR VPWR _12149_ sky130_fd_sc_hd__o2bb2a_1
X_24228_ _10599_ systolic_inst.A_shift\[19\]\[5\] net70 VGND VGND VPWR VPWR _02175_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24159_ systolic_inst.A_shift\[28\]\[3\] A_in\[99\] net59 VGND VGND VPWR VPWR _10581_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_227_Left_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28967_ clknet_leaf_53_clk _02765_ VGND VGND VPWR VPWR systolic_inst.B_shift\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16981_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[11\]\[0\]
+ _04286_ _04284_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a31o_1
XFILLER_104_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18720_ _05813_ _05815_ _05844_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__a21o_1
X_27918_ clknet_leaf_145_clk _01716_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_15932_ _12953_ _12954_ VGND VGND VPWR VPWR _12955_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_53_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28898_ clknet_leaf_279_clk _02696_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_231_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_202_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ _12894_ _12895_ VGND VGND VPWR VPWR _12897_ sky130_fd_sc_hd__nor2_1
X_18651_ _05775_ _05776_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_202_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27849_ clknet_leaf_179_clk _01647_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14814_ _11934_ _11937_ VGND VGND VPWR VPWR _11939_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17602_ _04844_ _04845_ _04846_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__and3_1
XFILLER_224_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15794_ net67 _12835_ _12837_ systolic_inst.acc_wires\[13\]\[6\] net107 VGND VGND
+ VPWR VPWR _01112_ sky130_fd_sc_hd__a32o_1
X_18582_ _05709_ _05710_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__and2_1
XFILLER_236_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ systolic_inst.A_outs\[14\]\[5\] systolic_inst.A_outs\[13\]\[5\] net116 VGND
+ VGND VPWR VPWR _01015_ sky130_fd_sc_hd__mux2_1
X_29519_ clknet_leaf_247_clk _03317_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[491\]
+ sky130_fd_sc_hd__dfrtp_1
X_17533_ _04742_ _04784_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17464_ _04716_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_190_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14676_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[22\]
+ VGND VGND VPWR VPWR _11832_ sky130_fd_sc_hd__nand2_1
XFILLER_177_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19203_ _06266_ _06267_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__nor2_1
X_16415_ _03780_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__nand2_1
X_13627_ deser_B.word_buffer\[63\] deser_B.serial_word\[63\] net123 VGND VGND VPWR
+ VPWR _00464_ sky130_fd_sc_hd__mux2_1
XFILLER_34_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17395_ _04649_ _04650_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__nor2_1
XFILLER_158_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19134_ _06176_ _06178_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__nand2_1
XFILLER_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16346_ _03724_ _03723_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__and2b_1
XFILLER_203_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13558_ deser_A.shift_reg\[122\] deser_A.shift_reg\[123\] net130 VGND VGND VPWR VPWR
+ _00395_ sky130_fd_sc_hd__mux2_1
XFILLER_242_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19065_ _06130_ _06132_ _06113_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__a21oi_1
XFILLER_195_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16277_ _03516_ _03657_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__or2_1
X_13489_ deser_A.shift_reg\[53\] deser_A.shift_reg\[54\] net130 VGND VGND VPWR VPWR
+ _00326_ sky130_fd_sc_hd__mux2_1
XFILLER_172_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15228_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[14\]\[12\]
+ VGND VGND VPWR VPWR _12330_ sky130_fd_sc_hd__xnor2_1
X_18016_ _05190_ _05207_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__xor2_1
XFILLER_126_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_209_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_209_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15159_ _12269_ _12270_ _12262_ _12265_ VGND VGND VPWR VPWR _12271_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_147_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19967_ _06895_ _06932_ _06931_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_147_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18918_ _06021_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_143_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19898_ systolic_inst.B_outs\[6\]\[5\] systolic_inst.A_outs\[6\]\[6\] VGND VGND VPWR
+ VPWR _06896_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_143_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18849_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[8\]\[8\]
+ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__nand2_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21860_ _08442_ _08582_ _08653_ _08651_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__a31oi_1
XFILLER_55_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20811_ _07710_ VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21791_ _08556_ _08595_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23530_ systolic_inst.B_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[6\] systolic_inst.A_outs\[0\]\[7\]
+ systolic_inst.B_outs\[0\]\[3\] VGND VGND VPWR VPWR _10153_ sky130_fd_sc_hd__a22oi_1
X_20742_ systolic_inst.acc_wires\[5\]\[16\] systolic_inst.acc_wires\[5\]\[17\] systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__o21a_1
XFILLER_24_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23461_ _10077_ _10085_ VGND VGND VPWR VPWR _10086_ sky130_fd_sc_hd__nand2_1
XFILLER_91_1150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20673_ _07591_ _07592_ net64 VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25200_ net110 ser_C.shift_reg\[428\] VGND VGND VPWR VPWR _11070_ sky130_fd_sc_hd__and2_1
X_22412_ _09150_ _09151_ VGND VGND VPWR VPWR _09153_ sky130_fd_sc_hd__xor2_1
XFILLER_108_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26180_ ser_C.bit_idx\[3\] _11303_ _11247_ VGND VGND VPWR VPWR _11249_ sky130_fd_sc_hd__a21oi_1
XFILLER_195_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23392_ _09984_ _10018_ VGND VGND VPWR VPWR _10019_ sky130_fd_sc_hd__nor2_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25131_ C_out\[392\] net101 net73 ser_C.shift_reg\[392\] _11035_ VGND VGND VPWR VPWR
+ _02642_ sky130_fd_sc_hd__a221o_1
X_22343_ _09083_ _09084_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25062_ net112 ser_C.shift_reg\[359\] VGND VGND VPWR VPWR _11001_ sky130_fd_sc_hd__and2_1
X_22274_ net109 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[8\] VGND
+ VGND VPWR VPWR _09019_ sky130_fd_sc_hd__and2_1
XFILLER_178_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24013_ systolic_inst.B_shift\[7\]\[4\] _11332_ net83 systolic_inst.B_shift\[11\]\[4\]
+ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__a22o_1
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21225_ _08041_ _08089_ _08091_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_93_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28821_ clknet_leaf_240_clk _02619_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[369\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_219_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21156_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[11\] _08025_ net117
+ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20107_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[6\]\[14\]
+ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__nand2_1
XFILLER_24_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21087_ _07953_ _07957_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__xnor2_1
X_25964_ systolic_inst.acc_wires\[13\]\[24\] ser_C.parallel_data\[440\] net19 VGND
+ VGND VPWR VPWR _03266_ sky130_fd_sc_hd__mux2_1
X_28752_ clknet_leaf_221_clk _02550_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[300\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27703_ clknet_leaf_192_clk _01501_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_20038_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[6\]\[4\]
+ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24915_ C_out\[284\] net103 net75 ser_C.shift_reg\[284\] _10927_ VGND VGND VPWR VPWR
+ _02534_ sky130_fd_sc_hd__a221o_1
XFILLER_74_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_219_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28683_ clknet_leaf_194_clk _02481_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[231\]
+ sky130_fd_sc_hd__dfrtp_1
X_25895_ systolic_inst.acc_wires\[11\]\[19\] C_out\[371\] net41 VGND VGND VPWR VPWR
+ _03197_ sky130_fd_sc_hd__mux2_1
XFILLER_73_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24846_ net113 ser_C.shift_reg\[251\] VGND VGND VPWR VPWR _10893_ sky130_fd_sc_hd__and2_1
X_27634_ clknet_leaf_324_clk _01432_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_218_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_215_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_215_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_234_Right_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27565_ clknet_leaf_299_clk _01363_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24777_ C_out\[215\] net98 net78 ser_C.shift_reg\[215\] _10858_ VGND VGND VPWR VPWR
+ _02465_ sky130_fd_sc_hd__a221o_1
X_21989_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[18\]
+ VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__or2_1
XFILLER_226_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14530_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[15\]\[1\]
+ VGND VGND VPWR VPWR _11707_ sky130_fd_sc_hd__and2_1
XFILLER_42_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29304_ clknet_leaf_325_clk _03102_ net142 VGND VGND VPWR VPWR C_out\[276\] sky130_fd_sc_hd__dfrtp_1
X_26516_ clknet_leaf_11_A_in_serial_clk _00319_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_230_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23728_ net63 _10337_ _10339_ systolic_inst.acc_wires\[0\]\[5\] _11258_ VGND VGND
+ VPWR VPWR _01935_ sky130_fd_sc_hd__a32o_1
XFILLER_187_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27496_ clknet_leaf_226_clk _01294_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29235_ clknet_leaf_183_clk _03033_ net146 VGND VGND VPWR VPWR C_out\[207\] sky130_fd_sc_hd__dfrtp_1
XFILLER_144_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26447_ clknet_leaf_346_clk _00254_ net132 VGND VGND VPWR VPWR A_in\[115\] sky130_fd_sc_hd__dfrtp_1
X_14461_ _11641_ _11642_ VGND VGND VPWR VPWR _11643_ sky130_fd_sc_hd__nor2_1
XFILLER_109_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23659_ _10244_ _10246_ _10276_ _10277_ VGND VGND VPWR VPWR _10279_ sky130_fd_sc_hd__a211o_1
XFILLER_202_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16200_ _03542_ _03544_ _03581_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__and3_1
XFILLER_35_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13412_ A_in\[121\] deser_A.word_buffer\[121\] _00003_ VGND VGND VPWR VPWR _00260_
+ sky130_fd_sc_hd__mux2_1
XFILLER_230_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29166_ clknet_leaf_39_clk _02964_ net141 VGND VGND VPWR VPWR C_out\[138\] sky130_fd_sc_hd__dfrtp_1
X_17180_ systolic_inst.A_outs\[10\]\[2\] systolic_inst.A_outs\[9\]\[2\] net120 VGND
+ VGND VPWR VPWR _01268_ sky130_fd_sc_hd__mux2_1
XFILLER_224_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14392_ _11573_ _11574_ VGND VGND VPWR VPWR _11576_ sky130_fd_sc_hd__nand2b_1
X_26378_ clknet_leaf_14_clk _00185_ net131 VGND VGND VPWR VPWR A_in\[46\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28117_ clknet_leaf_50_clk _01915_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_161_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16131_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[7\]
+ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__o21a_1
XFILLER_122_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25329_ ser_C.parallel_data\[491\] net97 net77 ser_C.shift_reg\[491\] _11134_ VGND
+ VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a221o_1
X_13343_ A_in\[52\] deser_A.word_buffer\[52\] net92 VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__mux2_1
X_29097_ clknet_leaf_154_clk _02895_ net150 VGND VGND VPWR VPWR C_out\[69\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_94_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28048_ clknet_leaf_131_clk _01846_ net144 VGND VGND VPWR VPWR systolic_inst.A_outs\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_16062_ _13056_ _13057_ VGND VGND VPWR VPWR _13058_ sky130_fd_sc_hd__nor2_1
X_13274_ deser_A.word_buffer\[112\] deser_A.serial_word\[112\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__mux2_1
XFILLER_108_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15013_ _12070_ _12095_ _12094_ VGND VGND VPWR VPWR _12133_ sky130_fd_sc_hd__a21boi_1
XFILLER_237_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19821_ _06789_ _06791_ _06788_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__o21ba_1
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_204_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19752_ systolic_inst.A_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[4\]
+ systolic_inst.B_outs\[6\]\[3\] VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__a22oi_1
XFILLER_42_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16964_ _04197_ _04257_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18703_ _05792_ _05797_ _05828_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_196_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15915_ _12939_ _12940_ VGND VGND VPWR VPWR _12941_ sky130_fd_sc_hd__or2_1
XFILLER_231_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19683_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[4\]
+ systolic_inst.A_outs\[6\]\[5\] VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__and4_1
XFILLER_77_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16895_ _04210_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__nand2_1
XFILLER_209_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18634_ _05724_ _05727_ _05760_ net108 VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__a31oi_1
XFILLER_237_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_192_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _12879_ _12880_ VGND VGND VPWR VPWR _12882_ sky130_fd_sc_hd__nand2_1
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_201_Right_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18565_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[7\]
+ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__o21a_1
XFILLER_18_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15777_ _12820_ _12821_ _12822_ VGND VGND VPWR VPWR _12823_ sky130_fd_sc_hd__a21o_1
XFILLER_221_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17516_ _04766_ _04767_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14728_ systolic_inst.acc_wires\[15\]\[28\] systolic_inst.acc_wires\[15\]\[29\] systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _11876_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18496_ systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[5\] systolic_inst.A_outs\[8\]\[6\]
+ systolic_inst.B_outs\[8\]\[0\] VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__a22oi_1
XFILLER_220_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14659_ _11816_ _11817_ VGND VGND VPWR VPWR _11818_ sky130_fd_sc_hd__xnor2_1
X_17447_ _04699_ _04700_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_180_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_180_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17378_ _04634_ _04633_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__and2b_1
XFILLER_14_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19117_ _06178_ _06179_ _06183_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__nand3_2
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16329_ _03676_ _03678_ _03708_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__o21a_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19048_ _06115_ _06116_ _06106_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__a21o_1
XFILLER_106_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21010_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[6\] VGND VGND VPWR
+ VPWR _07883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22961_ _09599_ _09601_ _09637_ VGND VGND VPWR VPWR _09639_ sky130_fd_sc_hd__nand3_1
XFILLER_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24700_ net113 ser_C.shift_reg\[178\] VGND VGND VPWR VPWR _10820_ sky130_fd_sc_hd__and2_1
XFILLER_210_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21912_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[3\]\[7\]
+ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__nand2_1
X_25680_ systolic_inst.acc_wires\[4\]\[28\] C_out\[156\] net32 VGND VGND VPWR VPWR
+ _02982_ sky130_fd_sc_hd__mux2_1
X_22892_ _09570_ _09571_ VGND VGND VPWR VPWR _09572_ sky130_fd_sc_hd__xnor2_1
X_24631_ C_out\[142\] net104 _10643_ ser_C.shift_reg\[142\] _10785_ VGND VGND VPWR
+ VPWR _02392_ sky130_fd_sc_hd__a221o_1
XFILLER_55_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21843_ _08620_ _08623_ _08645_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27350_ clknet_leaf_234_clk _01148_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_24562_ net113 ser_C.shift_reg\[109\] VGND VGND VPWR VPWR _10751_ sky130_fd_sc_hd__and2_1
XFILLER_208_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21774_ _08544_ _08548_ _08578_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__o21ai_1
XFILLER_184_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26301_ clknet_leaf_23_A_in_serial_clk _00109_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23513_ _10134_ _10135_ _10068_ _10071_ VGND VGND VPWR VPWR _10137_ sky130_fd_sc_hd__a211o_1
X_20725_ _07634_ _07635_ _07629_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__or3b_1
XFILLER_145_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27281_ clknet_leaf_321_clk _01079_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_93_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24493_ C_out\[73\] _11302_ net81 ser_C.shift_reg\[73\] _10716_ VGND VGND VPWR VPWR
+ _02323_ sky130_fd_sc_hd__a221o_1
XFILLER_211_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_171_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_171_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29020_ clknet_leaf_93_clk _02818_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_221_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26232_ clknet_leaf_6_A_in_serial_clk _00040_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_225_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23444_ _10066_ _10067_ _10065_ VGND VGND VPWR VPWR _10069_ sky130_fd_sc_hd__o21a_1
XFILLER_196_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20656_ net64 _07577_ _07579_ systolic_inst.acc_wires\[5\]\[5\] net109 VGND VGND
+ VPWR VPWR _01623_ sky130_fd_sc_hd__a32o_1
XFILLER_149_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26163_ deser_B.serial_word\[118\] deser_B.shift_reg\[118\] net56 VGND VGND VPWR
+ VPWR _03465_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23375_ _09998_ _10001_ VGND VGND VPWR VPWR _10002_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_59_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20587_ _07487_ _07516_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_95_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25114_ net110 ser_C.shift_reg\[385\] VGND VGND VPWR VPWR _11027_ sky130_fd_sc_hd__and2_1
X_22326_ _09068_ _09067_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__nand2b_1
XFILLER_125_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26094_ deser_B.serial_word\[49\] deser_B.shift_reg\[49\] net55 VGND VGND VPWR VPWR
+ _03396_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25045_ C_out\[349\] net98 net78 ser_C.shift_reg\[349\] _10992_ VGND VGND VPWR VPWR
+ _02599_ sky130_fd_sc_hd__a221o_1
X_22257_ _08999_ _09000_ VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_240_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_240_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21208_ _08071_ _08074_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_240_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22188_ _08933_ _08934_ _08922_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__or3b_1
XFILLER_160_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28804_ clknet_leaf_247_clk _02602_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[352\]
+ sky130_fd_sc_hd__dfrtp_1
X_21139_ _08006_ _08007_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_50_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26996_ clknet_leaf_18_B_in_serial_clk _00794_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13961_ deser_A.serial_word\[122\] deser_A.shift_reg\[122\] _00002_ VGND VGND VPWR
+ VPWR _00787_ sky130_fd_sc_hd__mux2_1
X_28735_ clknet_leaf_302_clk _02533_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[283\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25947_ systolic_inst.acc_wires\[13\]\[7\] C_out\[423\] net19 VGND VGND VPWR VPWR
+ _03249_ sky130_fd_sc_hd__mux2_1
XFILLER_8_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15700_ _12751_ _12752_ VGND VGND VPWR VPWR _12753_ sky130_fd_sc_hd__and2_1
XFILLER_234_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16680_ _03997_ _03998_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__nand3_2
XFILLER_235_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28666_ clknet_leaf_176_clk _02464_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[214\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25878_ systolic_inst.acc_wires\[11\]\[2\] C_out\[354\] net38 VGND VGND VPWR VPWR
+ _03180_ sky130_fd_sc_hd__mux2_1
X_13892_ deser_A.serial_word\[53\] deser_A.shift_reg\[53\] _00002_ VGND VGND VPWR
+ VPWR _00718_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_238_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_238_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24829_ C_out\[241\] net98 net78 ser_C.shift_reg\[241\] _10884_ VGND VGND VPWR VPWR
+ _02491_ sky130_fd_sc_hd__a221o_1
X_15631_ _12648_ _12685_ systolic_inst.A_outs\[13\]\[7\] VGND VGND VPWR VPWR _12686_
+ sky130_fd_sc_hd__and3b_1
X_27617_ clknet_leaf_321_clk _01415_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_28597_ clknet_leaf_41_clk _02395_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[145\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18350_ _05503_ _05507_ _05510_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__a21o_1
X_15562_ _12617_ _12618_ VGND VGND VPWR VPWR _12619_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_48_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27548_ clknet_leaf_299_clk _01346_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14513_ _11690_ _11691_ VGND VGND VPWR VPWR _11693_ sky130_fd_sc_hd__or2_1
X_17301_ _04558_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27479_ clknet_leaf_307_clk _01277_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15493_ systolic_inst.A_outs\[13\]\[2\] systolic_inst.B_outs\[13\]\[5\] VGND VGND
+ VPWR VPWR _12552_ sky130_fd_sc_hd__nand2_1
X_18281_ _05445_ _05448_ _05452_ _05447_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_162_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_162_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29218_ clknet_leaf_181_clk _03016_ net148 VGND VGND VPWR VPWR C_out\[190\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14444_ systolic_inst.B_outs\[15\]\[5\] systolic_inst.A_outs\[15\]\[7\] VGND VGND
+ VPWR VPWR _11626_ sky130_fd_sc_hd__nand2_1
X_17232_ _04475_ _04492_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17163_ _04440_ _04443_ _04442_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__o21a_1
X_29149_ clknet_leaf_174_clk _02947_ net150 VGND VGND VPWR VPWR C_out\[121\] sky130_fd_sc_hd__dfrtp_1
XFILLER_156_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14375_ systolic_inst.A_outs\[15\]\[6\] _11558_ _11557_ VGND VGND VPWR VPWR _11559_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_196_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16114_ _13072_ _03498_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_185_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13326_ A_in\[35\] deser_A.word_buffer\[35\] net94 VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__mux2_1
XFILLER_171_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17094_ _04379_ _04381_ _04388_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16045_ _13035_ _13040_ VGND VGND VPWR VPWR _13042_ sky130_fd_sc_hd__xor2_1
X_13257_ deser_A.word_buffer\[95\] deser_A.serial_word\[95\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__mux2_1
XFILLER_170_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13188_ deser_A.word_buffer\[26\] deser_A.serial_word\[26\] net128 VGND VGND VPWR
+ VPWR _00036_ sky130_fd_sc_hd__mux2_1
XFILLER_69_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19804_ _06787_ _06804_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__or2_1
XFILLER_97_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17996_ _05150_ _05187_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_140_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19735_ _06736_ _06737_ _06710_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16947_ _04260_ _04261_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__nor2_1
XFILLER_77_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19666_ _06653_ _06669_ _06670_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16878_ net119 _04193_ _04194_ _04195_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__a31o_1
XFILLER_53_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18617_ systolic_inst.A_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[5\] _05707_ _05706_
+ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__a31oi_1
X_15829_ _12843_ _12866_ _12856_ _12865_ VGND VGND VPWR VPWR _12867_ sky130_fd_sc_hd__o2bb2a_1
X_19597_ _06618_ _06621_ _06620_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__o21a_1
XFILLER_53_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18548_ _05641_ _05677_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__or2_1
XFILLER_80_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_153_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_153_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18479_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[3\] _05607_ _05608_
+ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_99_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20510_ _07435_ _07443_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_170_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21490_ _08302_ _08303_ _08304_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__a21o_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20441_ _07368_ _07376_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload330 clknet_leaf_174_clk VGND VGND VPWR VPWR clkload330/Y sky130_fd_sc_hd__clkinv_4
X_23160_ _09815_ _09817_ _09819_ systolic_inst.acc_wires\[1\]\[13\] net109 VGND VGND
+ VPWR VPWR _01887_ sky130_fd_sc_hd__a32o_1
X_20372_ _07307_ _07308_ _07309_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__and3_1
XFILLER_49_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload341 clknet_leaf_1_A_in_serial_clk VGND VGND VPWR VPWR clkload341/Y sky130_fd_sc_hd__bufinv_16
XFILLER_118_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload352 clknet_leaf_3_A_in_serial_clk VGND VGND VPWR VPWR clkload352/Y sky130_fd_sc_hd__clkinv_8
X_22111_ _08859_ _08860_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__nor2_1
XFILLER_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload60 clknet_leaf_1_clk VGND VGND VPWR VPWR clkload60/Y sky130_fd_sc_hd__clkinv_8
Xclkload363 clknet_leaf_16_A_in_serial_clk VGND VGND VPWR VPWR clkload363/X sky130_fd_sc_hd__clkbuf_4
XFILLER_238_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload374 clknet_leaf_28_B_in_serial_clk VGND VGND VPWR VPWR clkload374/Y sky130_fd_sc_hd__bufinv_16
Xclkload71 clknet_leaf_348_clk VGND VGND VPWR VPWR clkload71/Y sky130_fd_sc_hd__inv_8
X_23091_ net64 _09758_ _09760_ systolic_inst.acc_wires\[1\]\[3\] _11258_ VGND VGND
+ VPWR VPWR _01877_ sky130_fd_sc_hd__a32o_1
Xclkload385 clknet_leaf_5_B_in_serial_clk VGND VGND VPWR VPWR clkload385/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload82 clknet_leaf_28_clk VGND VGND VPWR VPWR clkload82/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload93 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload93/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22042_ systolic_inst.acc_wires\[3\]\[24\] systolic_inst.acc_wires\[3\]\[25\] systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__o21a_1
XFILLER_173_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26850_ clknet_leaf_66_clk _00652_ net134 VGND VGND VPWR VPWR B_in\[122\] sky130_fd_sc_hd__dfrtp_1
XFILLER_87_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25801_ systolic_inst.acc_wires\[8\]\[21\] C_out\[277\] net28 VGND VGND VPWR VPWR
+ _03103_ sky130_fd_sc_hd__mux2_1
XFILLER_87_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26781_ clknet_leaf_54_clk _00583_ net137 VGND VGND VPWR VPWR B_in\[53\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23993_ systolic_inst.B_shift\[9\]\[0\] B_in\[8\] _00008_ VGND VGND VPWR VPWR _10522_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28520_ clknet_leaf_155_clk _02318_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[68\]
+ sky130_fd_sc_hd__dfrtp_1
X_25732_ systolic_inst.acc_wires\[6\]\[16\] C_out\[208\] net46 VGND VGND VPWR VPWR
+ _03034_ sky130_fd_sc_hd__mux2_1
X_22944_ _09515_ _09621_ VGND VGND VPWR VPWR _09622_ sky130_fd_sc_hd__or2_1
XFILLER_25_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25663_ systolic_inst.acc_wires\[4\]\[11\] C_out\[139\] net30 VGND VGND VPWR VPWR
+ _02965_ sky130_fd_sc_hd__mux2_1
XFILLER_44_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28451_ clknet_leaf_35_clk _02249_ VGND VGND VPWR VPWR systolic_inst.A_shift\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_22875_ _09515_ _09553_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__and2_1
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27402_ clknet_leaf_333_clk _01200_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_24614_ net110 ser_C.shift_reg\[135\] VGND VGND VPWR VPWR _10777_ sky130_fd_sc_hd__and2_1
XFILLER_188_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21826_ _08585_ _08599_ _08597_ VGND VGND VPWR VPWR _08630_ sky130_fd_sc_hd__o21a_1
X_28382_ clknet_leaf_33_clk _02180_ VGND VGND VPWR VPWR systolic_inst.A_shift\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_233_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25594_ systolic_inst.acc_wires\[2\]\[6\] C_out\[70\] net34 VGND VGND VPWR VPWR _02896_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_159_Left_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_233_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27333_ clknet_leaf_286_clk _01131_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24545_ C_out\[99\] net99 net79 ser_C.shift_reg\[99\] _10742_ VGND VGND VPWR VPWR
+ _02349_ sky130_fd_sc_hd__a221o_1
XFILLER_145_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21757_ _08562_ _08561_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_144_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20708_ _07615_ _07616_ _07623_ VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__a21o_1
XFILLER_129_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27264_ clknet_leaf_269_clk _01062_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24476_ net112 ser_C.shift_reg\[66\] VGND VGND VPWR VPWR _10708_ sky130_fd_sc_hd__and2_1
X_21688_ _08495_ _08494_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__nand2b_1
XFILLER_145_1198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29003_ clknet_leaf_104_clk _02801_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_26215_ clknet_leaf_12_A_in_serial_clk _00023_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23427_ _10033_ _10051_ VGND VGND VPWR VPWR _10053_ sky130_fd_sc_hd__nand2_1
X_20639_ _07562_ _07563_ _07564_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__and3_1
X_27195_ clknet_leaf_254_clk _00993_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26146_ deser_B.serial_word\[101\] deser_B.shift_reg\[101\] _00001_ VGND VGND VPWR
+ VPWR _03448_ sky130_fd_sc_hd__mux2_1
X_14160_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[0\] systolic_inst.B_outs\[15\]\[3\]
+ systolic_inst.A_outs\[15\]\[3\] VGND VGND VPWR VPWR _11351_ sky130_fd_sc_hd__and4_1
X_23358_ _09965_ _09985_ VGND VGND VPWR VPWR _09986_ sky130_fd_sc_hd__nand2b_1
XFILLER_50_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_242_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13111_ systolic_inst.A_outs\[0\]\[4\] VGND VGND VPWR VPWR _11267_ sky130_fd_sc_hd__inv_2
XFILLER_125_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_242_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22309_ _09047_ _09050_ _09051_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__and3_1
X_26077_ deser_B.serial_word\[32\] deser_B.shift_reg\[32\] net55 VGND VGND VPWR VPWR
+ _03379_ sky130_fd_sc_hd__mux2_1
X_14091_ deser_B.shift_reg\[125\] deser_B.shift_reg\[126\] net126 VGND VGND VPWR VPWR
+ _00917_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_168_Left_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23289_ net121 _09920_ VGND VGND VPWR VPWR _09921_ sky130_fd_sc_hd__nand2_1
XFILLER_152_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25028_ net112 ser_C.shift_reg\[342\] VGND VGND VPWR VPWR _10984_ sky130_fd_sc_hd__and2_1
XFILLER_156_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xload_slew108 _11258_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_16
XFILLER_65_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17850_ _05044_ _05046_ _05027_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16801_ _04081_ _04083_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__a21o_1
XFILLER_117_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17781_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[31\]
+ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__xnor2_1
X_26979_ clknet_leaf_28_A_in_serial_clk _00777_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_14993_ systolic_inst.A_outs\[14\]\[3\] systolic_inst.A_outs\[14\]\[4\] systolic_inst.B_outs\[14\]\[6\]
+ systolic_inst.B_outs\[14\]\[7\] VGND VGND VPWR VPWR _12113_ sky130_fd_sc_hd__and4b_1
XFILLER_208_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19520_ _06559_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__inv_2
XFILLER_8_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28718_ clknet_leaf_314_clk _02516_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[266\]
+ sky130_fd_sc_hd__dfrtp_1
X_16732_ _03990_ _04025_ _04024_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a21bo_1
XFILLER_219_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13944_ deser_A.serial_word\[105\] deser_A.shift_reg\[105\] net57 VGND VGND VPWR
+ VPWR _00770_ sky130_fd_sc_hd__mux2_1
X_29698_ clknet_5_21__leaf_clk VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_178_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19451_ net62 _06499_ _06500_ systolic_inst.acc_wires\[7\]\[7\] net105 VGND VGND
+ VPWR VPWR _01497_ sky130_fd_sc_hd__a32o_1
X_28649_ clknet_leaf_202_clk _02447_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[197\]
+ sky130_fd_sc_hd__dfrtp_1
X_16663_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[5\] _03985_
+ _03986_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__a22o_1
X_13875_ deser_A.serial_word\[36\] deser_A.shift_reg\[36\] net58 VGND VGND VPWR VPWR
+ _00701_ sky130_fd_sc_hd__mux2_1
XFILLER_235_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_177_Left_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18402_ _05555_ _05554_ systolic_inst.acc_wires\[9\]\[31\] net105 VGND VGND VPWR
+ VPWR _01393_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15614_ _12613_ _12668_ VGND VGND VPWR VPWR _12670_ sky130_fd_sc_hd__xnor2_1
X_19382_ _06375_ _06418_ _06417_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__o21a_1
X_16594_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[1\]
+ systolic_inst.B_outs\[11\]\[0\] VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__a22o_1
X_18333_ net64 _05496_ _05497_ systolic_inst.acc_wires\[9\]\[20\] net106 VGND VGND
+ VPWR VPWR _01382_ sky130_fd_sc_hd__a32o_1
XFILLER_203_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15545_ _12573_ _12602_ VGND VGND VPWR VPWR _12603_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_135_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_37_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15476_ _12504_ _12535_ VGND VGND VPWR VPWR _12536_ sky130_fd_sc_hd__xnor2_1
X_18264_ _05430_ _05432_ _05436_ _11713_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__a31o_1
XFILLER_204_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14427_ _11609_ _11608_ VGND VGND VPWR VPWR _11610_ sky130_fd_sc_hd__and2b_1
X_17215_ _04465_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__or2_1
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18195_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[9\]\[1\]
+ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__nand2_1
XFILLER_200_1115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17146_ _04424_ _04426_ _04432_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__a21o_1
X_14358_ _11541_ _11542_ VGND VGND VPWR VPWR _11543_ sky130_fd_sc_hd__and2_1
XFILLER_239_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13309_ A_in\[18\] deser_A.word_buffer\[18\] net91 VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__mux2_1
XFILLER_170_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17077_ _04358_ _04365_ _04371_ _04364_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__a211o_1
XFILLER_239_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14289_ _11439_ _11441_ VGND VGND VPWR VPWR _11475_ sky130_fd_sc_hd__or2_1
XFILLER_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16028_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[5\] VGND
+ VGND VPWR VPWR _13025_ sky130_fd_sc_hd__and2_1
XFILLER_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17979_ _05154_ _05171_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__or2_1
XFILLER_84_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19718_ systolic_inst.A_outs\[6\]\[2\] systolic_inst.B_outs\[6\]\[3\] systolic_inst.A_outs\[6\]\[3\]
+ systolic_inst.B_outs\[6\]\[4\] VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__and4_1
X_20990_ _07863_ _07862_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__nand2b_1
XFILLER_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19649_ systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[3\]
+ systolic_inst.B_outs\[6\]\[0\] VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__a22o_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22660_ net109 systolic_inst.acc_wires\[2\]\[29\] net65 _09367_ VGND VGND VPWR VPWR
+ _01839_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_172_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21611_ _08387_ _08419_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22591_ systolic_inst.acc_wires\[2\]\[16\] systolic_inst.acc_wires\[2\]\[17\] systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__o21a_1
XFILLER_179_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_126_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_61_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24330_ _10638_ systolic_inst.A_shift\[9\]\[4\] net70 VGND VGND VPWR VPWR _02238_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21542_ systolic_inst.A_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[5\] VGND VGND VPWR
+ VPWR _08354_ sky130_fd_sc_hd__nand2_1
XFILLER_166_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24261_ systolic_inst.A_shift\[16\]\[4\] net70 net83 systolic_inst.A_shift\[17\]\[4\]
+ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__a22o_1
X_21473_ systolic_inst.B_outs\[2\]\[1\] systolic_inst.B_shift\[2\]\[1\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__mux2_1
XFILLER_222_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26000_ systolic_inst.acc_wires\[14\]\[28\] ser_C.parallel_data\[476\] net24 VGND
+ VGND VPWR VPWR _03302_ sky130_fd_sc_hd__mux2_1
XFILLER_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23212_ _09854_ _09860_ _09861_ _11713_ VGND VGND VPWR VPWR _09864_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_116_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20424_ _07287_ _07329_ _07328_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__o21ba_1
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24192_ systolic_inst.A_shift\[24\]\[7\] net70 _10505_ systolic_inst.A_shift\[25\]\[7\]
+ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__a22o_1
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23143_ _09803_ _09804_ VGND VGND VPWR VPWR _09805_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20355_ _07257_ _07292_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__and2_1
XFILLER_135_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload160 clknet_leaf_219_clk VGND VGND VPWR VPWR clkload160/Y sky130_fd_sc_hd__clkinv_8
XFILLER_135_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload171 clknet_leaf_244_clk VGND VGND VPWR VPWR clkload171/Y sky130_fd_sc_hd__bufinv_16
XFILLER_88_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload182 clknet_leaf_238_clk VGND VGND VPWR VPWR clkload182/Y sky130_fd_sc_hd__bufinv_16
Xclkload193 clknet_leaf_65_clk VGND VGND VPWR VPWR clkload193/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_162_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23074_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[1\]\[0\]
+ _09744_ _09745_ VGND VGND VPWR VPWR _09746_ sky130_fd_sc_hd__and4_1
X_27951_ clknet_leaf_171_clk _01749_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_129_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20286_ _07207_ _07224_ _07225_ net109 VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_73_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22025_ net106 systolic_inst.acc_wires\[3\]\[23\] net65 _08802_ VGND VGND VPWR VPWR
+ _01769_ sky130_fd_sc_hd__a22o_1
X_26902_ clknet_leaf_16_A_in_serial_clk _00700_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_222_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27882_ clknet_leaf_45_clk _01680_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29621_ clknet_leaf_6_B_in_serial_clk _03416_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26833_ clknet_leaf_89_clk _00635_ net5 VGND VGND VPWR VPWR B_in\[105\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29552_ clknet_leaf_3_B_in_serial_clk _03347_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_217_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26764_ clknet_leaf_80_clk _00566_ net144 VGND VGND VPWR VPWR B_in\[36\] sky130_fd_sc_hd__dfrtp_1
X_23976_ _10513_ systolic_inst.B_shift\[9\]\[7\] _11332_ VGND VGND VPWR VPWR _02009_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_235_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_235_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28503_ clknet_leaf_113_clk _02301_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22927_ _09603_ _09604_ VGND VGND VPWR VPWR _09606_ sky130_fd_sc_hd__xor2_1
X_25715_ systolic_inst.acc_wires\[5\]\[31\] C_out\[191\] net43 VGND VGND VPWR VPWR
+ _03017_ sky130_fd_sc_hd__mux2_1
XFILLER_57_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26695_ clknet_leaf_5_B_in_serial_clk _00498_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_29483_ clknet_leaf_271_clk _03281_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_231_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13660_ deser_B.word_buffer\[96\] deser_B.serial_word\[96\] net123 VGND VGND VPWR
+ VPWR _00497_ sky130_fd_sc_hd__mux2_1
XFILLER_72_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28434_ clknet_leaf_28_clk _02232_ VGND VGND VPWR VPWR systolic_inst.A_shift\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_231_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25646_ systolic_inst.acc_wires\[3\]\[26\] C_out\[122\] net50 VGND VGND VPWR VPWR
+ _02948_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22858_ _09520_ _09538_ VGND VGND VPWR VPWR _09539_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21809_ _08612_ _08613_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__nor2_1
XFILLER_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25577_ systolic_inst.acc_wires\[1\]\[21\] C_out\[53\] net53 VGND VGND VPWR VPWR
+ _02879_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_117_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13591_ deser_B.word_buffer\[27\] deser_B.serial_word\[27\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__mux2_1
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28365_ clknet_leaf_29_clk _02163_ VGND VGND VPWR VPWR systolic_inst.A_shift\[20\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_22789_ _09448_ _09470_ _09471_ VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__nand3_1
XFILLER_25_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15330_ net107 systolic_inst.acc_wires\[14\]\[27\] _11712_ _12416_ VGND VGND VPWR
+ VPWR _01069_ sky130_fd_sc_hd__a22o_1
X_24528_ net114 ser_C.shift_reg\[92\] VGND VGND VPWR VPWR _10734_ sky130_fd_sc_hd__and2_1
XFILLER_200_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27316_ clknet_leaf_290_clk _01114_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_169_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28296_ clknet_leaf_121_clk _02094_ VGND VGND VPWR VPWR systolic_inst.B_shift\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15261_ net61 _12358_ VGND VGND VPWR VPWR _12359_ sky130_fd_sc_hd__nor2_1
X_24459_ C_out\[56\] net100 net82 ser_C.shift_reg\[56\] _10699_ VGND VGND VPWR VPWR
+ _02306_ sky130_fd_sc_hd__a221o_1
XFILLER_201_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27247_ clknet_leaf_274_clk _01045_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_229_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14212_ _11373_ _11375_ _11400_ VGND VGND VPWR VPWR _11401_ sky130_fd_sc_hd__a21oi_1
X_17000_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[11\]\[5\]
+ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__nand2_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15192_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[14\]\[7\]
+ VGND VGND VPWR VPWR _12299_ sky130_fd_sc_hd__or2_1
X_27178_ clknet_leaf_247_clk _00976_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_165_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_8 systolic_inst.A_outs\[5\]\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26129_ deser_B.serial_word\[84\] deser_B.shift_reg\[84\] net56 VGND VGND VPWR VPWR
+ _03431_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14143_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[1\]
+ systolic_inst.B_outs\[15\]\[1\] VGND VGND VPWR VPWR _11336_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_39_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14074_ deser_B.shift_reg\[108\] deser_B.shift_reg\[109\] deser_B.receiving VGND
+ VGND VPWR VPWR _00900_ sky130_fd_sc_hd__mux2_1
X_18951_ systolic_inst.acc_wires\[8\]\[20\] systolic_inst.acc_wires\[8\]\[21\] systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__o21a_1
XFILLER_98_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17902_ _05091_ _05095_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__xor2_1
X_18882_ _05984_ _05987_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__a21oi_1
XFILLER_239_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17833_ systolic_inst.A_outs\[9\]\[0\] systolic_inst.A_outs\[9\]\[1\] systolic_inst.B_outs\[9\]\[3\]
+ systolic_inst.B_outs\[9\]\[4\] VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__nand4_1
XFILLER_0_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17764_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[28\]
+ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__nand2_1
X_14976_ _12056_ _12058_ _12096_ VGND VGND VPWR VPWR _12097_ sky130_fd_sc_hd__and3_1
XFILLER_212_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19503_ net62 _06544_ _06545_ systolic_inst.acc_wires\[7\]\[14\] net105 VGND VGND
+ VPWR VPWR _01504_ sky130_fd_sc_hd__a32o_1
XFILLER_35_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16715_ _04001_ _04036_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__xnor2_1
X_13927_ deser_A.serial_word\[88\] deser_A.shift_reg\[88\] net57 VGND VGND VPWR VPWR
+ _00753_ sky130_fd_sc_hd__mux2_1
X_17695_ _04924_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19434_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[7\]\[5\]
+ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__nand2_1
XFILLER_39_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_179_Right_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16646_ systolic_inst.A_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[2\] systolic_inst.B_outs\[11\]\[3\]
+ systolic_inst.B_outs\[11\]\[4\] VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__and4_1
XFILLER_165_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13858_ deser_A.serial_word\[19\] deser_A.shift_reg\[19\] net58 VGND VGND VPWR VPWR
+ _00684_ sky130_fd_sc_hd__mux2_1
XFILLER_62_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19365_ _06391_ _06393_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_108_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16577_ systolic_inst.A_outs\[11\]\[2\] systolic_inst.A_outs\[10\]\[2\] net118 VGND
+ VGND VPWR VPWR _01204_ sky130_fd_sc_hd__mux2_1
XFILLER_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13789_ B_in\[96\] deser_B.word_buffer\[96\] net89 VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__mux2_1
XFILLER_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18316_ _05474_ _05476_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__nand2_1
X_15528_ _12584_ _12585_ VGND VGND VPWR VPWR _12586_ sky130_fd_sc_hd__xnor2_1
X_19296_ _06348_ _06356_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18247_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[9\]\[9\]
+ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__nor2_1
XFILLER_30_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15459_ systolic_inst.A_outs\[13\]\[1\] systolic_inst.B_outs\[13\]\[5\] systolic_inst.B_outs\[13\]\[6\]
+ systolic_inst.A_outs\[13\]\[0\] VGND VGND VPWR VPWR _12519_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_152_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18178_ _05362_ _05363_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17129_ _04374_ _04375_ _04397_ _04417_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__a211o_1
XFILLER_143_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20140_ net106 systolic_inst.acc_wires\[6\]\[18\] net62 _07114_ VGND VGND VPWR VPWR
+ _01572_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_165_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20071_ _07050_ _07053_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__nand2_1
XFILLER_44_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23830_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[20\]
+ _10424_ VGND VGND VPWR VPWR _10426_ sky130_fd_sc_hd__a21bo_1
XFILLER_57_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23761_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[0\]\[11\]
+ VGND VGND VPWR VPWR _10367_ sky130_fd_sc_hd__nor2_1
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_347_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_347_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20973_ systolic_inst.B_outs\[4\]\[5\] _07845_ _07846_ VGND VGND VPWR VPWR _07847_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_38_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25500_ _00008_ _11228_ VGND VGND VPWR VPWR _11230_ sky130_fd_sc_hd__nor2_1
XFILLER_214_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22712_ _09392_ _09397_ VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__nand2_1
XFILLER_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26480_ clknet_leaf_13_A_in_serial_clk _00283_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_23692_ net121 systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[0\]\[0\]
+ VGND VGND VPWR VPWR _10309_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25431_ systolic_inst.A_shift\[1\]\[7\] A_in\[7\] net59 VGND VGND VPWR VPWR _11185_
+ sky130_fd_sc_hd__mux2_1
X_22643_ net109 systolic_inst.acc_wires\[2\]\[26\] net65 _09353_ VGND VGND VPWR VPWR
+ _01836_ sky130_fd_sc_hd__a22o_1
XFILLER_213_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28150_ clknet_leaf_108_clk _01948_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25362_ net112 ser_C.shift_reg\[509\] VGND VGND VPWR VPWR _11151_ sky130_fd_sc_hd__and2_1
XFILLER_90_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22574_ _09291_ _09292_ _09286_ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_118_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27101_ clknet_leaf_8_B_in_serial_clk _00899_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_178_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24313_ systolic_inst.A_shift\[11\]\[4\] A_in\[44\] net59 VGND VGND VPWR VPWR _10630_
+ sky130_fd_sc_hd__mux2_1
X_28081_ clknet_leaf_115_clk _01879_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_194_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21525_ _08316_ _08319_ _08337_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__a21o_1
XFILLER_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25293_ ser_C.parallel_data\[473\] net102 net74 ser_C.shift_reg\[473\] _11116_ VGND
+ VGND VPWR VPWR _02723_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27032_ clknet_leaf_12_B_in_serial_clk _00830_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_193_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24244_ _10607_ systolic_inst.A_shift\[18\]\[5\] net70 VGND VGND VPWR VPWR _02183_
+ sky130_fd_sc_hd__mux2_1
X_21456_ _08289_ _08290_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20407_ _07342_ _07343_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__or2_1
X_24175_ systolic_inst.A_shift\[26\]\[6\] net70 _10505_ systolic_inst.A_shift\[27\]\[6\]
+ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__a22o_1
XFILLER_108_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_224_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21387_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[20\]
+ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_224_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23126_ _09785_ _09788_ VGND VGND VPWR VPWR _09790_ sky130_fd_sc_hd__nand2_1
XFILLER_190_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20338_ _07244_ _07275_ _07276_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__nand3_1
X_28983_ clknet_leaf_57_clk _02781_ VGND VGND VPWR VPWR systolic_inst.A_shift\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27934_ clknet_leaf_180_clk _01732_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_23057_ _09679_ _09684_ _09706_ _09708_ VGND VGND VPWR VPWR _09732_ sky130_fd_sc_hd__o31a_1
XFILLER_163_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20269_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.A_outs\[5\]\[1\] systolic_inst.B_outs\[5\]\[3\]
+ systolic_inst.B_outs\[5\]\[4\] VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__nand4_1
XFILLER_62_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22008_ _08786_ _08787_ _08784_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__o21ai_2
XFILLER_131_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27865_ clknet_leaf_143_clk _01663_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29604_ clknet_leaf_25_B_in_serial_clk _03399_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_26816_ clknet_leaf_63_clk _00618_ net135 VGND VGND VPWR VPWR B_in\[88\] sky130_fd_sc_hd__dfrtp_1
X_14830_ _11953_ _11954_ VGND VGND VPWR VPWR _11955_ sky130_fd_sc_hd__and2_1
XFILLER_76_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27796_ clknet_leaf_45_clk _01594_ net137 VGND VGND VPWR VPWR systolic_inst.B_outs\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29535_ clknet_leaf_258_clk _03333_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[507\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26747_ clknet_leaf_52_clk _00549_ net143 VGND VGND VPWR VPWR B_in\[19\] sky130_fd_sc_hd__dfrtp_1
X_14761_ net118 _11889_ VGND VGND VPWR VPWR _11890_ sky130_fd_sc_hd__and2_1
XFILLER_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23959_ systolic_inst.B_shift\[11\]\[6\] _11332_ net83 systolic_inst.B_shift\[15\]\[6\]
+ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_338_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_338_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_45_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16500_ _03851_ _03855_ _03857_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__a21oi_1
X_13712_ B_in\[19\] deser_B.word_buffer\[19\] net86 VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__mux2_1
XFILLER_17_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29466_ clknet_leaf_287_clk _03264_ net136 VGND VGND VPWR VPWR C_out\[438\] sky130_fd_sc_hd__dfrtp_1
X_14692_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[24\]
+ VGND VGND VPWR VPWR _11846_ sky130_fd_sc_hd__nor2_1
X_17480_ _04733_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__inv_2
XFILLER_232_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26678_ clknet_leaf_11_B_in_serial_clk _00481_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28417_ clknet_leaf_70_clk _02215_ VGND VGND VPWR VPWR systolic_inst.B_shift\[23\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16431_ _03784_ _03785_ _03790_ _03797_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__a31o_1
X_25629_ systolic_inst.acc_wires\[3\]\[9\] C_out\[105\] net48 VGND VGND VPWR VPWR
+ _02931_ sky130_fd_sc_hd__mux2_1
X_13643_ deser_B.word_buffer\[79\] deser_B.serial_word\[79\] net123 VGND VGND VPWR
+ VPWR _00480_ sky130_fd_sc_hd__mux2_1
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29397_ clknet_leaf_241_clk _03195_ net145 VGND VGND VPWR VPWR C_out\[369\] sky130_fd_sc_hd__dfrtp_1
XFILLER_147_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19150_ _06181_ _06214_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13574_ deser_B.word_buffer\[10\] deser_B.serial_word\[10\] net124 VGND VGND VPWR
+ VPWR _00411_ sky130_fd_sc_hd__mux2_1
X_16362_ _03736_ _03739_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28348_ clknet_leaf_319_clk _02146_ VGND VGND VPWR VPWR systolic_inst.A_shift\[24\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18101_ _05149_ _05288_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__nand2_1
X_15313_ _12397_ _12399_ _12402_ VGND VGND VPWR VPWR _12403_ sky130_fd_sc_hd__a21oi_2
XFILLER_34_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19081_ _06145_ _06148_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__xor2_1
XFILLER_125_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16293_ _03660_ _03673_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__xor2_1
XFILLER_201_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28279_ clknet_leaf_130_clk _02077_ VGND VGND VPWR VPWR systolic_inst.B_shift\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18032_ systolic_inst.B_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[6\] systolic_inst.A_outs\[9\]\[7\]
+ systolic_inst.B_outs\[9\]\[3\] VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__a22o_1
XFILLER_173_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15244_ _12329_ _12337_ _12343_ VGND VGND VPWR VPWR _12344_ sky130_fd_sc_hd__o21ai_1
XFILLER_173_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15175_ _12284_ VGND VGND VPWR VPWR _12285_ sky130_fd_sc_hd__inv_2
XFILLER_201_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14126_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.A_outs\[14\]\[2\] net118 VGND
+ VGND VPWR VPWR _00948_ sky130_fd_sc_hd__mux2_1
X_19983_ systolic_inst.B_outs\[6\]\[5\] systolic_inst.B_outs\[6\]\[6\] systolic_inst.A_outs\[6\]\[7\]
+ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__nand3_1
XFILLER_158_1175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1006 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14057_ deser_B.shift_reg\[91\] deser_B.shift_reg\[92\] net126 VGND VGND VPWR VPWR
+ _00883_ sky130_fd_sc_hd__mux2_1
X_18934_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[20\]
+ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__or2_1
XFILLER_45_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_207_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18865_ _05967_ _05971_ _05974_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_105_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17816_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[2\] _05013_
+ _05014_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__a22o_1
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18796_ _05909_ _05917_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__nand2_1
XFILLER_227_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17747_ _04965_ _04967_ _04969_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_329_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_329_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_47_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14959_ systolic_inst.A_outs\[14\]\[4\] systolic_inst.B_outs\[14\]\[5\] VGND VGND
+ VPWR VPWR _12080_ sky130_fd_sc_hd__nand2_1
XFILLER_130_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17678_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[15\]
+ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_158_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19417_ _06471_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__inv_2
XFILLER_35_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16629_ _03952_ _03953_ _03935_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19348_ _06406_ _06407_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__nor2_1
XFILLER_17_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_114_Left_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19279_ net119 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[11\] VGND
+ VGND VPWR VPWR _06341_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_14_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21310_ _08164_ _08165_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__and2b_1
XFILLER_191_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22290_ _09030_ _09033_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21241_ _08052_ _08053_ _08083_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__or3_1
XFILLER_144_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21172_ _07923_ _08040_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_70_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20123_ _07098_ _07099_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__and2_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Left_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25980_ systolic_inst.acc_wires\[14\]\[8\] ser_C.parallel_data\[456\] net25 VGND
+ VGND VPWR VPWR _03282_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_215_Right_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_A_in_serial_clk clknet_2_1__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_19_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20054_ _07038_ _07039_ _07040_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__a21o_1
XFILLER_113_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24931_ C_out\[292\] net102 net74 ser_C.shift_reg\[292\] _10935_ VGND VGND VPWR VPWR
+ _02542_ sky130_fd_sc_hd__a221o_1
XFILLER_58_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27650_ clknet_leaf_326_clk _01448_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_24862_ net110 ser_C.shift_reg\[259\] VGND VGND VPWR VPWR _10901_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_107_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26601_ clknet_leaf_18_B_in_serial_clk _00404_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23813_ _10410_ _10411_ VGND VGND VPWR VPWR _10412_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24793_ C_out\[223\] net99 net79 ser_C.shift_reg\[223\] _10866_ VGND VGND VPWR VPWR
+ _02473_ sky130_fd_sc_hd__a221o_1
X_27581_ clknet_leaf_220_clk _01379_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_68_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29320_ clknet_leaf_298_clk _03118_ net138 VGND VGND VPWR VPWR C_out\[292\] sky130_fd_sc_hd__dfrtp_1
X_23744_ _10351_ _10352_ VGND VGND VPWR VPWR _10353_ sky130_fd_sc_hd__and2_1
X_26532_ clknet_leaf_5_A_in_serial_clk _00335_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_217_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20956_ _07796_ _07799_ _07830_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__o21a_1
XFILLER_214_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29251_ clknet_leaf_184_clk _03049_ net146 VGND VGND VPWR VPWR C_out\[223\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23675_ _10292_ _10293_ VGND VGND VPWR VPWR _10294_ sky130_fd_sc_hd__and2_1
X_26463_ clknet_leaf_1_A_in_serial_clk _00270_ net132 VGND VGND VPWR VPWR deser_A.bit_idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_132_Left_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20887_ _07762_ _07763_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__nand2_1
XFILLER_242_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28202_ clknet_leaf_129_clk _02000_ VGND VGND VPWR VPWR systolic_inst.B_shift\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_22626_ _09319_ _09338_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__nor2_1
XFILLER_198_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25414_ _11176_ systolic_inst.A_shift\[1\]\[6\] net70 VGND VGND VPWR VPWR _02784_
+ sky130_fd_sc_hd__mux2_1
X_29182_ clknet_leaf_44_clk _02980_ net142 VGND VGND VPWR VPWR C_out\[154\] sky130_fd_sc_hd__dfrtp_1
XFILLER_139_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26394_ clknet_leaf_12_clk _00201_ net134 VGND VGND VPWR VPWR A_in\[62\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28133_ clknet_leaf_128_clk _01931_ net144 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_25345_ ser_C.parallel_data\[499\] net102 net77 ser_C.shift_reg\[499\] _11142_ VGND
+ VGND VPWR VPWR _02749_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_12_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22557_ _09272_ _09273_ _09280_ VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__a21o_1
XFILLER_107_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21508_ _08320_ _08321_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__and2b_1
X_28064_ clknet_leaf_120_clk _01862_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25276_ net111 ser_C.shift_reg\[466\] VGND VGND VPWR VPWR _11108_ sky130_fd_sc_hd__and2_1
X_13290_ deser_A.serial_toggle deser_A.serial_word_ready VGND VGND VPWR VPWR _00138_
+ sky130_fd_sc_hd__xor2_1
X_22488_ _09219_ _09220_ _09221_ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__a21o_1
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27015_ clknet_leaf_22_B_in_serial_clk _00813_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_24227_ systolic_inst.A_shift\[20\]\[5\] A_in\[77\] net59 VGND VGND VPWR VPWR _10599_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21439_ _08269_ _08273_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__nor2_1
XFILLER_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24158_ _10580_ systolic_inst.A_shift\[27\]\[2\] net70 VGND VGND VPWR VPWR _02124_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_141_Left_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23109_ _09773_ _09774_ _09775_ VGND VGND VPWR VPWR _09776_ sky130_fd_sc_hd__a21o_1
XFILLER_194_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28966_ clknet_leaf_52_clk _02764_ VGND VGND VPWR VPWR systolic_inst.B_shift\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24089_ systolic_inst.B_shift\[23\]\[0\] B_in\[56\] net59 VGND VGND VPWR VPWR _10554_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16980_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[11\]\[2\]
+ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__or2_1
XFILLER_150_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27917_ clknet_leaf_145_clk _01715_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_15931_ _12947_ _12951_ _12948_ VGND VGND VPWR VPWR _12954_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_53_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28897_ clknet_leaf_284_clk _02695_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[445\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _05776_ _05775_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__nand2b_1
XFILLER_231_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27848_ clknet_leaf_179_clk _01646_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15862_ _12894_ _12895_ VGND VGND VPWR VPWR _12896_ sky130_fd_sc_hd__nand2_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17601_ _04839_ _04840_ _04838_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__a21bo_1
XFILLER_190_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14813_ _11937_ _11934_ VGND VGND VPWR VPWR _11938_ sky130_fd_sc_hd__nand2b_1
XFILLER_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18581_ systolic_inst.A_outs\[8\]\[2\] systolic_inst.B_outs\[8\]\[5\] _05673_ _05672_
+ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__a31o_1
X_27779_ clknet_leaf_186_clk _01577_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_15793_ _12836_ VGND VGND VPWR VPWR _12837_ sky130_fd_sc_hd__inv_2
XFILLER_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29518_ clknet_leaf_247_clk _03316_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[490\]
+ sky130_fd_sc_hd__dfrtp_1
X_17532_ _04781_ _04782_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__xor2_1
X_14744_ systolic_inst.A_outs\[14\]\[4\] systolic_inst.A_outs\[13\]\[4\] net116 VGND
+ VGND VPWR VPWR _01014_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_150_Left_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_190_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29449_ clknet_leaf_293_clk _03247_ net139 VGND VGND VPWR VPWR C_out\[421\] sky130_fd_sc_hd__dfrtp_1
X_17463_ systolic_inst.A_outs\[10\]\[5\] systolic_inst.B_outs\[10\]\[6\] _11275_ systolic_inst.A_outs\[10\]\[4\]
+ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__o2bb2a_1
X_14675_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[22\]
+ VGND VGND VPWR VPWR _11831_ sky130_fd_sc_hd__or2_1
X_19202_ _06226_ _06228_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__nor2_1
X_16414_ net67 _03782_ _03783_ systolic_inst.acc_wires\[12\]\[7\] net108 VGND VGND
+ VPWR VPWR _01177_ sky130_fd_sc_hd__a32o_1
XFILLER_60_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13626_ deser_B.word_buffer\[62\] deser_B.serial_word\[62\] net123 VGND VGND VPWR
+ VPWR _00463_ sky130_fd_sc_hd__mux2_1
X_17394_ systolic_inst.A_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[6\] _11275_ systolic_inst.A_outs\[10\]\[2\]
+ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_34_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19133_ _06147_ _06174_ _06173_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16345_ _03660_ _03702_ _03701_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__o21a_1
XFILLER_125_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13557_ deser_A.shift_reg\[121\] deser_A.shift_reg\[122\] net130 VGND VGND VPWR VPWR
+ _00394_ sky130_fd_sc_hd__mux2_1
XFILLER_157_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19064_ _06113_ _06130_ _06132_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__and3_1
X_16276_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[7\] _03630_ _03594_
+ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__a31o_1
X_13488_ deser_A.shift_reg\[52\] deser_A.shift_reg\[53\] net130 VGND VGND VPWR VPWR
+ _00325_ sky130_fd_sc_hd__mux2_1
XFILLER_185_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18015_ _05205_ _05206_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__nand2_1
X_15227_ _12317_ _12326_ _12327_ _12328_ VGND VGND VPWR VPWR _12329_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_209_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15158_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[14\]\[2\]
+ VGND VGND VPWR VPWR _12270_ sky130_fd_sc_hd__or2_1
XFILLER_236_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14109_ systolic_inst.B_shift\[12\]\[1\] net72 _11333_ B_in\[97\] VGND VGND VPWR
+ VPWR _00931_ sky130_fd_sc_hd__a22o_1
X_19966_ _06960_ _06961_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15089_ systolic_inst.A_outs\[14\]\[6\] _11264_ VGND VGND VPWR VPWR _12206_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_147_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18917_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[17\]
+ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__xor2_2
XFILLER_80_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19897_ _06825_ _06894_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_143_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18848_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[8\]\[8\]
+ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__or2_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18779_ _05835_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20810_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[29\]
+ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__xor2_1
XFILLER_36_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21790_ _08592_ _08593_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20741_ _07650_ _07651_ VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__nand2_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23460_ _10082_ _10083_ VGND VGND VPWR VPWR _10085_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20672_ _07591_ _07592_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__and2_1
XFILLER_52_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22411_ _09085_ _09088_ _09118_ _09150_ _09116_ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__o311a_1
XFILLER_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23391_ _09968_ _10016_ VGND VGND VPWR VPWR _10018_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_108_1394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25130_ net110 ser_C.shift_reg\[393\] VGND VGND VPWR VPWR _11035_ sky130_fd_sc_hd__and2_1
X_22342_ _09083_ _09084_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__nor2_1
XFILLER_163_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25061_ C_out\[357\] net98 net78 ser_C.shift_reg\[357\] _11000_ VGND VGND VPWR VPWR
+ _02607_ sky130_fd_sc_hd__a221o_1
X_22273_ _09015_ _09016_ VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__nand2b_1
XFILLER_219_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24012_ systolic_inst.B_shift\[7\]\[3\] _11332_ net83 systolic_inst.B_shift\[11\]\[3\]
+ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21224_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.B_outs\[4\]\[6\] systolic_inst.A_outs\[4\]\[7\]
+ _08090_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__a31oi_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28820_ clknet_leaf_239_clk _02618_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[368\]
+ sky130_fd_sc_hd__dfrtp_1
X_21155_ _08023_ _08024_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_109_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20106_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[6\]\[14\]
+ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__or2_1
XFILLER_28_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28751_ clknet_leaf_221_clk _02549_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21086_ _07954_ _07956_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__nand2_1
XFILLER_28_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25963_ systolic_inst.acc_wires\[13\]\[23\] C_out\[439\] net19 VGND VGND VPWR VPWR
+ _03265_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_97_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27702_ clknet_leaf_198_clk _01500_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20037_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[6\]\[4\]
+ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__nand2_1
XFILLER_4_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24914_ net110 ser_C.shift_reg\[285\] VGND VGND VPWR VPWR _10927_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_219_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28682_ clknet_leaf_196_clk _02480_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_115_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25894_ systolic_inst.acc_wires\[11\]\[18\] C_out\[370\] net41 VGND VGND VPWR VPWR
+ _03196_ sky130_fd_sc_hd__mux2_1
XFILLER_160_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27633_ clknet_leaf_324_clk _01431_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24845_ C_out\[249\] net98 net78 ser_C.shift_reg\[249\] _10892_ VGND VGND VPWR VPWR
+ _02499_ sky130_fd_sc_hd__a221o_1
XFILLER_234_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_215_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27564_ clknet_leaf_299_clk _01362_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_21988_ net106 systolic_inst.acc_wires\[3\]\[17\] net65 _08771_ VGND VGND VPWR VPWR
+ _01763_ sky130_fd_sc_hd__a22o_1
X_24776_ net113 ser_C.shift_reg\[216\] VGND VGND VPWR VPWR _10858_ sky130_fd_sc_hd__and2_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29303_ clknet_leaf_325_clk _03101_ net142 VGND VGND VPWR VPWR C_out\[275\] sky130_fd_sc_hd__dfrtp_1
XFILLER_215_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26515_ clknet_leaf_11_A_in_serial_clk _00318_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_23727_ _10338_ VGND VGND VPWR VPWR _10339_ sky130_fd_sc_hd__inv_2
X_20939_ _07810_ _07813_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__xor2_1
X_27495_ clknet_leaf_227_clk _01293_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_215_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29234_ clknet_leaf_205_clk _03032_ net146 VGND VGND VPWR VPWR C_out\[206\] sky130_fd_sc_hd__dfrtp_1
XFILLER_42_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26446_ clknet_leaf_346_clk _00253_ net132 VGND VGND VPWR VPWR A_in\[114\] sky130_fd_sc_hd__dfrtp_1
X_14460_ _11554_ _11611_ _11610_ VGND VGND VPWR VPWR _11642_ sky130_fd_sc_hd__a21oi_1
XFILLER_241_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23658_ _10276_ _10277_ _10244_ _10246_ VGND VGND VPWR VPWR _10278_ sky130_fd_sc_hd__o211ai_1
XFILLER_144_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ A_in\[120\] deser_A.word_buffer\[120\] _00003_ VGND VGND VPWR VPWR _00259_
+ sky130_fd_sc_hd__mux2_1
X_22609_ net109 systolic_inst.acc_wires\[2\]\[21\] net65 _09324_ VGND VGND VPWR VPWR
+ _01831_ sky130_fd_sc_hd__a22o_1
XFILLER_167_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29165_ clknet_leaf_39_clk _02963_ net141 VGND VGND VPWR VPWR C_out\[137\] sky130_fd_sc_hd__dfrtp_1
X_14391_ _11574_ _11573_ VGND VGND VPWR VPWR _11575_ sky130_fd_sc_hd__nand2b_1
XFILLER_168_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23589_ _10167_ _10170_ _10210_ VGND VGND VPWR VPWR _10211_ sky130_fd_sc_hd__o21a_1
X_26377_ clknet_leaf_29_clk _00184_ net133 VGND VGND VPWR VPWR A_in\[45\] sky130_fd_sc_hd__dfrtp_1
XFILLER_128_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_195_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28116_ clknet_leaf_128_clk _01914_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_16130_ _13095_ _13097_ _13096_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__o21bai_1
X_13342_ A_in\[51\] deser_A.word_buffer\[51\] net95 VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25328_ net112 ser_C.shift_reg\[492\] VGND VGND VPWR VPWR _11134_ sky130_fd_sc_hd__and2_1
X_29096_ clknet_leaf_155_clk _02894_ net150 VGND VGND VPWR VPWR C_out\[68\] sky130_fd_sc_hd__dfrtp_1
XFILLER_182_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28047_ clknet_leaf_130_clk _01845_ net144 VGND VGND VPWR VPWR systolic_inst.A_outs\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_16061_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[5\]
+ systolic_inst.A_outs\[12\]\[6\] VGND VGND VPWR VPWR _13057_ sky130_fd_sc_hd__and4_1
X_13273_ deser_A.word_buffer\[111\] deser_A.serial_word\[111\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__mux2_1
X_25259_ ser_C.parallel_data\[456\] net102 net74 ser_C.shift_reg\[456\] _11099_ VGND
+ VGND VPWR VPWR _02706_ sky130_fd_sc_hd__a221o_1
XFILLER_237_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15012_ _12130_ _12131_ VGND VGND VPWR VPWR _12132_ sky130_fd_sc_hd__nand2_1
XFILLER_170_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19820_ _06780_ _06786_ _06785_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_183_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_204_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19751_ systolic_inst.B_outs\[6\]\[3\] systolic_inst.A_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\]
+ systolic_inst.A_outs\[6\]\[4\] VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__and4_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28949_ clknet_leaf_261_clk _02747_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[497\]
+ sky130_fd_sc_hd__dfrtp_1
X_16963_ _04200_ _04262_ _04260_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_88_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
X_18702_ _05826_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_196_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15914_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[24\]
+ VGND VGND VPWR VPWR _12940_ sky130_fd_sc_hd__and2_1
XFILLER_42_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_196_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19682_ systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[5\]
+ systolic_inst.B_outs\[6\]\[0\] VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__a22oi_1
XFILLER_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16894_ _04176_ _04178_ _04209_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__nand3_1
XFILLER_231_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18633_ _05724_ _05727_ _05760_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__a21o_1
XFILLER_225_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15845_ _12879_ _12880_ VGND VGND VPWR VPWR _12881_ sky130_fd_sc_hd__and2_1
XFILLER_237_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18564_ _05665_ _05667_ _05666_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__o21bai_1
X_15776_ _12815_ _12816_ _12814_ VGND VGND VPWR VPWR _12822_ sky130_fd_sc_hd__a21bo_1
XFILLER_220_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17515_ _04701_ _04705_ _04735_ _04766_ _04734_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_16_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ net105 systolic_inst.acc_wires\[15\]\[29\] net69 _11875_ VGND VGND VPWR VPWR
+ _01007_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18495_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[3\] _05609_ _05607_
+ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__a31o_1
XFILLER_221_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17446_ _04699_ _04700_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__nor2_1
X_14658_ _11812_ _11814_ _11811_ VGND VGND VPWR VPWR _11817_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13609_ deser_B.word_buffer\[45\] deser_B.serial_word\[45\] net124 VGND VGND VPWR
+ VPWR _00446_ sky130_fd_sc_hd__mux2_1
X_17377_ _04595_ _04596_ _04594_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__a21oi_1
XFILLER_242_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14589_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[15\]\[8\]
+ _11754_ VGND VGND VPWR VPWR _11758_ sky130_fd_sc_hd__and3_1
XFILLER_158_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
X_19116_ _06180_ _06182_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__nor2_1
XFILLER_119_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16328_ _03659_ _03707_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__xnor2_1
XFILLER_229_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19047_ _06106_ _06115_ _06116_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__nand3_1
XFILLER_174_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16259_ _03632_ _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_149_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19949_ _06944_ _06945_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__and2_1
XFILLER_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_79_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_214_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22960_ _09599_ _09601_ _09637_ VGND VGND VPWR VPWR _09638_ sky130_fd_sc_hd__a21o_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21911_ net68 _08703_ _08705_ systolic_inst.acc_wires\[3\]\[6\] net106 VGND VGND
+ VPWR VPWR _01752_ sky130_fd_sc_hd__a32o_1
XFILLER_56_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22891_ _09525_ _09534_ _09533_ VGND VGND VPWR VPWR _09571_ sky130_fd_sc_hd__o21ba_1
XFILLER_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21842_ _08643_ _08644_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__or2_1
X_24630_ net7 ser_C.shift_reg\[143\] VGND VGND VPWR VPWR _10785_ sky130_fd_sc_hd__and2_1
XFILLER_167_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24561_ C_out\[107\] net100 net80 ser_C.shift_reg\[107\] _10750_ VGND VGND VPWR VPWR
+ _02357_ sky130_fd_sc_hd__a221o_1
XFILLER_93_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21773_ _08544_ _08548_ _08578_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_121_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26300_ clknet_leaf_23_A_in_serial_clk _00108_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_184_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20724_ net64 _07636_ _07637_ systolic_inst.acc_wires\[5\]\[15\] net109 VGND VGND
+ VPWR VPWR _01633_ sky130_fd_sc_hd__a32o_1
X_23512_ _10068_ _10071_ _10134_ _10135_ VGND VGND VPWR VPWR _10136_ sky130_fd_sc_hd__o211ai_4
XFILLER_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24492_ net112 ser_C.shift_reg\[74\] VGND VGND VPWR VPWR _10716_ sky130_fd_sc_hd__and2_1
X_27280_ clknet_leaf_323_clk _01078_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_223_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23443_ _10065_ _10066_ _10067_ VGND VGND VPWR VPWR _10068_ sky130_fd_sc_hd__nor3_2
X_26231_ clknet_leaf_6_A_in_serial_clk _00039_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20655_ _07578_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__inv_2
XFILLER_177_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23374_ _09999_ _10000_ VGND VGND VPWR VPWR _10001_ sky130_fd_sc_hd__or2_1
X_26162_ deser_B.serial_word\[117\] deser_B.shift_reg\[117\] net56 VGND VGND VPWR
+ VPWR _03464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20586_ _07491_ _07516_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22325_ _09030_ _09032_ _09031_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__o21ba_1
X_25113_ C_out\[383\] net97 net77 ser_C.shift_reg\[383\] _11026_ VGND VGND VPWR VPWR
+ _02633_ sky130_fd_sc_hd__a221o_1
XFILLER_30_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26093_ deser_B.serial_word\[48\] deser_B.shift_reg\[48\] net55 VGND VGND VPWR VPWR
+ _03395_ sky130_fd_sc_hd__mux2_1
XFILLER_178_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25044_ net113 ser_C.shift_reg\[350\] VGND VGND VPWR VPWR _10992_ sky130_fd_sc_hd__and2_1
X_22256_ _09000_ _08999_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__nand2b_1
XFILLER_191_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_240_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21207_ _08071_ _08074_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__and2_1
XFILLER_219_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_240_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22187_ _08931_ _08932_ _08903_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28803_ clknet_leaf_244_clk _02601_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_152_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21138_ _08006_ _08007_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__and2_1
XFILLER_78_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26995_ clknet_leaf_18_B_in_serial_clk _00793_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28734_ clknet_leaf_302_clk _02532_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[282\]
+ sky130_fd_sc_hd__dfrtp_1
X_21069_ _07939_ _07940_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__nor2_1
X_25946_ systolic_inst.acc_wires\[13\]\[6\] C_out\[422\] net26 VGND VGND VPWR VPWR
+ _03248_ sky130_fd_sc_hd__mux2_1
X_13960_ deser_A.serial_word\[121\] deser_A.shift_reg\[121\] _00002_ VGND VGND VPWR
+ VPWR _00786_ sky130_fd_sc_hd__mux2_1
XFILLER_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28665_ clknet_leaf_176_clk _02463_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[213\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_150_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25877_ systolic_inst.acc_wires\[11\]\[1\] C_out\[353\] net39 VGND VGND VPWR VPWR
+ _03179_ sky130_fd_sc_hd__mux2_1
X_13891_ deser_A.serial_word\[52\] deser_A.shift_reg\[52\] net58 VGND VGND VPWR VPWR
+ _00717_ sky130_fd_sc_hd__mux2_1
XFILLER_235_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_238_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_238_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ systolic_inst.B_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\] VGND VGND
+ VPWR VPWR _12685_ sky130_fd_sc_hd__or2_1
X_27616_ clknet_leaf_321_clk _01414_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24828_ net113 ser_C.shift_reg\[242\] VGND VGND VPWR VPWR _10884_ sky130_fd_sc_hd__and2_1
X_28596_ clknet_leaf_41_clk _02394_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[144\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_222_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ systolic_inst.B_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[5\]
+ systolic_inst.A_outs\[13\]\[6\] VGND VGND VPWR VPWR _12618_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_48_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27547_ clknet_leaf_35_clk _01345_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_203_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24759_ C_out\[206\] net99 net79 ser_C.shift_reg\[206\] _10849_ VGND VGND VPWR VPWR
+ _02456_ sky130_fd_sc_hd__a221o_1
XFILLER_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17300_ _04502_ _04528_ _04527_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14512_ _11690_ _11691_ VGND VGND VPWR VPWR _11692_ sky130_fd_sc_hd__nor2_1
X_18280_ _05450_ _05451_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__nand2_1
X_27478_ clknet_leaf_306_clk _01276_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15492_ _12547_ _12550_ VGND VGND VPWR VPWR _12551_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29217_ clknet_leaf_179_clk _03015_ net148 VGND VGND VPWR VPWR C_out\[189\] sky130_fd_sc_hd__dfrtp_1
X_17231_ _04476_ _04490_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__a21oi_1
X_26429_ clknet_leaf_3_clk _00236_ net131 VGND VGND VPWR VPWR A_in\[97\] sky130_fd_sc_hd__dfrtp_1
X_14443_ _11623_ _11624_ VGND VGND VPWR VPWR _11625_ sky130_fd_sc_hd__nor2_1
XFILLER_230_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29148_ clknet_leaf_175_clk _02946_ net150 VGND VGND VPWR VPWR C_out\[120\] sky130_fd_sc_hd__dfrtp_1
XFILLER_156_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17162_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__inv_2
XFILLER_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14374_ systolic_inst.B_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[7\]
+ VGND VGND VPWR VPWR _11558_ sky130_fd_sc_hd__and3_1
XFILLER_156_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16113_ _13072_ _03498_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_185_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13325_ A_in\[34\] deser_A.word_buffer\[34\] net94 VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__mux2_1
X_29079_ clknet_leaf_114_clk _02877_ net150 VGND VGND VPWR VPWR C_out\[51\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_185_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17093_ systolic_inst.acc_wires\[11\]\[16\] systolic_inst.acc_wires\[11\]\[17\] systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__o21a_1
XFILLER_122_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16044_ _13035_ _13040_ VGND VGND VPWR VPWR _13041_ sky130_fd_sc_hd__nand2b_1
XFILLER_143_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13256_ deser_A.word_buffer\[94\] deser_A.serial_word\[94\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13187_ deser_A.word_buffer\[25\] deser_A.serial_word\[25\] net128 VGND VGND VPWR
+ VPWR _00035_ sky130_fd_sc_hd__mux2_1
XFILLER_124_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19803_ _06802_ _06803_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17995_ _05156_ _05158_ _05155_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__o21ba_1
XFILLER_97_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19734_ _06734_ _06735_ _06704_ _06707_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__o211a_1
X_16946_ _04234_ _04236_ _04259_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__and3_1
XFILLER_133_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_38_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19665_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[3\]
+ systolic_inst.A_outs\[6\]\[4\] VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__and4_1
XFILLER_42_1178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16877_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[11\] VGND
+ VGND VPWR VPWR _04195_ sky130_fd_sc_hd__and2_1
XFILLER_20_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18616_ _05740_ _05743_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__xnor2_1
X_15828_ _12849_ _12865_ VGND VGND VPWR VPWR _12866_ sky130_fd_sc_hd__nor2_1
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19596_ _06623_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__inv_2
XFILLER_231_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18547_ _05669_ _05675_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_138_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15759_ net66 _12806_ _12807_ systolic_inst.acc_wires\[13\]\[1\] net107 VGND VGND
+ VPWR VPWR _01107_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_138_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18478_ _05607_ _05609_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[3\]
+ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_99_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17429_ _04648_ _04650_ _04649_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__o21ba_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20440_ _07373_ _07374_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload320 clknet_leaf_155_clk VGND VGND VPWR VPWR clkload320/Y sky130_fd_sc_hd__clkinv_2
X_20371_ _07273_ _07275_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__nand2_1
XFILLER_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload331 clknet_leaf_159_clk VGND VGND VPWR VPWR clkload331/Y sky130_fd_sc_hd__clkinv_4
XFILLER_174_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload342 clknet_leaf_2_A_in_serial_clk VGND VGND VPWR VPWR clkload342/Y sky130_fd_sc_hd__clkinv_4
X_22110_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.A_outs\[2\]\[1\] systolic_inst.B_outs\[2\]\[2\]
+ systolic_inst.B_outs\[2\]\[3\] VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__and4_1
XFILLER_162_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload50 clknet_leaf_291_clk VGND VGND VPWR VPWR clkload50/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload353 clknet_leaf_4_A_in_serial_clk VGND VGND VPWR VPWR clkload353/Y sky130_fd_sc_hd__bufinv_16
XFILLER_106_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23090_ _09759_ VGND VGND VPWR VPWR _09760_ sky130_fd_sc_hd__inv_2
Xclkload61 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload61/Y sky130_fd_sc_hd__clkinv_4
Xclkload364 clknet_leaf_17_A_in_serial_clk VGND VGND VPWR VPWR clkload364/Y sky130_fd_sc_hd__clkinv_2
Xclkload375 clknet_leaf_29_B_in_serial_clk VGND VGND VPWR VPWR clkload375/Y sky130_fd_sc_hd__bufinv_16
Xclkload72 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload72/Y sky130_fd_sc_hd__clkinv_2
Xclkload386 clknet_leaf_6_B_in_serial_clk VGND VGND VPWR VPWR clkload386/Y sky130_fd_sc_hd__bufinv_16
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload83 clknet_leaf_29_clk VGND VGND VPWR VPWR clkload83/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload94 clknet_leaf_35_clk VGND VGND VPWR VPWR clkload94/X sky130_fd_sc_hd__clkbuf_4
X_22041_ _08814_ _08815_ VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_168_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25800_ systolic_inst.acc_wires\[8\]\[20\] C_out\[276\] net22 VGND VGND VPWR VPWR
+ _03102_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26780_ clknet_leaf_54_clk _00582_ net143 VGND VGND VPWR VPWR B_in\[52\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23992_ _10521_ systolic_inst.B_shift\[8\]\[7\] net72 VGND VGND VPWR VPWR _02017_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25731_ systolic_inst.acc_wires\[6\]\[15\] C_out\[207\] net43 VGND VGND VPWR VPWR
+ _03033_ sky130_fd_sc_hd__mux2_1
X_22943_ systolic_inst.A_outs\[1\]\[6\] _09590_ _09591_ _09557_ VGND VGND VPWR VPWR
+ _09621_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_123_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28450_ clknet_leaf_35_clk _02248_ VGND VGND VPWR VPWR systolic_inst.A_shift\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25662_ systolic_inst.acc_wires\[4\]\[10\] C_out\[138\] net29 VGND VGND VPWR VPWR
+ _02964_ sky130_fd_sc_hd__mux2_1
XFILLER_216_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22874_ _09515_ _09553_ VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__nor2_1
XFILLER_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27401_ clknet_leaf_332_clk _01199_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24613_ C_out\[133\] net103 net75 ser_C.shift_reg\[133\] _10776_ VGND VGND VPWR VPWR
+ _02383_ sky130_fd_sc_hd__a221o_1
XFILLER_110_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21825_ _08586_ _08628_ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__xnor2_1
X_28381_ clknet_leaf_34_clk _02179_ VGND VGND VPWR VPWR systolic_inst.A_shift\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25593_ systolic_inst.acc_wires\[2\]\[5\] C_out\[69\] net34 VGND VGND VPWR VPWR _02895_
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_233_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_233_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27332_ clknet_leaf_287_clk _01130_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_24544_ net113 ser_C.shift_reg\[100\] VGND VGND VPWR VPWR _10742_ sky130_fd_sc_hd__and2_1
X_21756_ _08522_ _08524_ _08523_ VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__o21ba_1
XFILLER_197_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_894 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20707_ _07617_ _07621_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__nand2b_1
XFILLER_106_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27263_ clknet_leaf_269_clk _01061_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_24475_ C_out\[64\] _11302_ net81 ser_C.shift_reg\[64\] _10707_ VGND VGND VPWR VPWR
+ _02314_ sky130_fd_sc_hd__a221o_1
X_21687_ _08453_ _08455_ _08454_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__o21ba_1
XFILLER_106_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29002_ clknet_leaf_103_clk _02800_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26214_ clknet_leaf_12_A_in_serial_clk _00022_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload0 clknet_5_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_8
X_23426_ _10033_ _10051_ VGND VGND VPWR VPWR _10052_ sky130_fd_sc_hd__or2_2
X_20638_ _07557_ _07558_ _07556_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__a21bo_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27194_ clknet_leaf_256_clk _00992_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_165_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26145_ deser_B.serial_word\[100\] deser_B.shift_reg\[100\] _00001_ VGND VGND VPWR
+ VPWR _03447_ sky130_fd_sc_hd__mux2_1
X_23357_ _09982_ _09983_ VGND VGND VPWR VPWR _09985_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20569_ _07499_ _07500_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__and2_1
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_242_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_242_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22308_ _09048_ _09049_ VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__nor2_1
X_13110_ systolic_inst.A_outs\[0\]\[2\] VGND VGND VPWR VPWR _11266_ sky130_fd_sc_hd__inv_2
X_14090_ deser_B.shift_reg\[124\] deser_B.shift_reg\[125\] net126 VGND VGND VPWR VPWR
+ _00916_ sky130_fd_sc_hd__mux2_1
X_26076_ deser_B.serial_word\[31\] deser_B.shift_reg\[31\] net55 VGND VGND VPWR VPWR
+ _03378_ sky130_fd_sc_hd__mux2_1
X_23288_ systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[1\] systolic_inst.A_outs\[0\]\[1\]
+ systolic_inst.B_outs\[0\]\[0\] VGND VGND VPWR VPWR _09920_ sky130_fd_sc_hd__a22o_1
XFILLER_124_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22239_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[7\]
+ VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_180_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25027_ C_out\[340\] net97 net77 ser_C.shift_reg\[340\] _10983_ VGND VGND VPWR VPWR
+ _02590_ sky130_fd_sc_hd__a221o_1
XFILLER_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_29__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_29__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_121_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xload_slew109 _11258_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_37_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16800_ _04092_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17780_ net62 _04997_ _04998_ systolic_inst.acc_wires\[10\]\[30\] net105 VGND VGND
+ VPWR VPWR _01328_ sky130_fd_sc_hd__a32o_1
XFILLER_232_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26978_ clknet_leaf_28_A_in_serial_clk _00776_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_14992_ systolic_inst.B_outs\[14\]\[5\] systolic_inst.A_outs\[14\]\[5\] VGND VGND
+ VPWR VPWR _12112_ sky130_fd_sc_hd__nand2_1
X_28717_ clknet_leaf_314_clk _02515_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[265\]
+ sky130_fd_sc_hd__dfrtp_1
X_16731_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[7\] _04052_ net119
+ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__mux2_1
X_25929_ systolic_inst.acc_wires\[12\]\[21\] C_out\[405\] net17 VGND VGND VPWR VPWR
+ _03231_ sky130_fd_sc_hd__mux2_1
X_13943_ deser_A.serial_word\[104\] deser_A.shift_reg\[104\] net57 VGND VGND VPWR
+ VPWR _00769_ sky130_fd_sc_hd__mux2_1
X_29697_ clknet_leaf_106_clk _00007_ net151 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_178_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_178_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19450_ _06491_ _06495_ _06497_ _06498_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__o211ai_2
X_28648_ clknet_leaf_202_clk _02446_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[196\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16662_ _03983_ _03984_ net119 VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__o21a_1
XFILLER_234_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13874_ deser_A.serial_word\[35\] deser_A.shift_reg\[35\] net58 VGND VGND VPWR VPWR
+ _00700_ sky130_fd_sc_hd__mux2_1
XFILLER_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18401_ _05548_ _05552_ _05553_ net60 VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__a31o_1
XFILLER_90_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15613_ _12613_ _12668_ VGND VGND VPWR VPWR _12669_ sky130_fd_sc_hd__nand2_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19381_ _06375_ _06439_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__xnor2_1
X_28579_ clknet_leaf_168_clk _02377_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_16593_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.A_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\]
+ systolic_inst.A_outs\[11\]\[1\] VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__and4_1
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18332_ _05494_ _05495_ _05491_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__o21ai_2
X_15544_ _12599_ _12600_ VGND VGND VPWR VPWR _12602_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18263_ _05430_ _05432_ _05436_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__a21oi_1
XFILLER_230_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15475_ _12533_ _12534_ VGND VGND VPWR VPWR _12535_ sky130_fd_sc_hd__nor2_1
XFILLER_188_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17214_ systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[3\] VGND VGND
+ VPWR VPWR _04476_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14426_ _11556_ _11572_ _11571_ VGND VGND VPWR VPWR _11609_ sky130_fd_sc_hd__o21ba_1
XFILLER_198_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18194_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[9\]\[1\]
+ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__and2_1
XFILLER_204_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17145_ systolic_inst.acc_wires\[11\]\[24\] systolic_inst.acc_wires\[11\]\[25\] systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__o21a_1
X_14357_ _11498_ _11500_ _11540_ VGND VGND VPWR VPWR _11542_ sky130_fd_sc_hd__or3_1
XFILLER_200_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13308_ A_in\[17\] deser_A.word_buffer\[17\] net91 VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__mux2_1
XFILLER_171_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17076_ _04373_ _04372_ systolic_inst.acc_wires\[11\]\[15\] net105 VGND VGND VPWR
+ VPWR _01249_ sky130_fd_sc_hd__a2bb2o_1
X_14288_ _11406_ _11445_ _11444_ VGND VGND VPWR VPWR _11474_ sky130_fd_sc_hd__a21o_1
XFILLER_100_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16027_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[4\] _13024_
+ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__a21bo_1
XFILLER_100_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13239_ deser_A.word_buffer\[77\] deser_A.serial_word\[77\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__mux2_1
XFILLER_174_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17978_ _05169_ _05170_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__xnor2_1
XFILLER_215_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19717_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[4\] VGND VGND VPWR
+ VPWR _06720_ sky130_fd_sc_hd__nand2_1
X_16929_ _04242_ _04243_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__and2b_1
XFILLER_211_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19648_ _06642_ _06653_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__or2_1
XFILLER_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19579_ systolic_inst.acc_wires\[7\]\[24\] systolic_inst.acc_wires\[7\]\[25\] systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__o21a_1
XFILLER_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21610_ systolic_inst.A_outs\[3\]\[1\] systolic_inst.B_outs\[3\]\[6\] _08419_ VGND
+ VGND VPWR VPWR _08420_ sky130_fd_sc_hd__and3_1
XFILLER_90_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22590_ _09307_ _09308_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__nand2_1
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21541_ _08331_ _08351_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24260_ systolic_inst.A_shift\[16\]\[3\] net70 net83 systolic_inst.A_shift\[17\]\[3\]
+ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__a22o_1
X_21472_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_shift\[2\]\[0\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__mux2_1
XFILLER_53_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23211_ _09854_ _09860_ _09861_ VGND VGND VPWR VPWR _09863_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20423_ _07320_ _07326_ _07325_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_116_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24191_ systolic_inst.A_shift\[24\]\[6\] net70 _10505_ systolic_inst.A_shift\[25\]\[6\]
+ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23142_ _09796_ _09798_ _09794_ VGND VGND VPWR VPWR _09804_ sky130_fd_sc_hd__a21bo_1
XFILLER_119_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20354_ _07285_ _07291_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__xor2_1
XFILLER_31_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload150 clknet_leaf_298_clk VGND VGND VPWR VPWR clkload150/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload161 clknet_leaf_220_clk VGND VGND VPWR VPWR clkload161/Y sky130_fd_sc_hd__inv_8
XFILLER_49_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload172 clknet_leaf_245_clk VGND VGND VPWR VPWR clkload172/Y sky130_fd_sc_hd__bufinv_16
XFILLER_162_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload183 clknet_leaf_239_clk VGND VGND VPWR VPWR clkload183/X sky130_fd_sc_hd__clkbuf_8
X_23073_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[1\]\[1\]
+ VGND VGND VPWR VPWR _09745_ sky130_fd_sc_hd__or2_1
X_27950_ clknet_leaf_180_clk _01748_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload194 clknet_leaf_66_clk VGND VGND VPWR VPWR clkload194/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_129_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20285_ _07224_ _07225_ _07207_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_129_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22024_ _08800_ _08801_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__xor2_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26901_ clknet_leaf_16_A_in_serial_clk _00699_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_161_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27881_ clknet_leaf_46_clk _01679_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_222_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29620_ clknet_leaf_6_B_in_serial_clk _03415_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26832_ clknet_leaf_87_clk _00634_ net144 VGND VGND VPWR VPWR B_in\[104\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29551_ clknet_leaf_110_clk _03346_ net151 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26763_ clknet_leaf_80_clk _00565_ net144 VGND VGND VPWR VPWR B_in\[35\] sky130_fd_sc_hd__dfrtp_1
XFILLER_151_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23975_ systolic_inst.B_shift\[13\]\[7\] B_in\[47\] _00008_ VGND VGND VPWR VPWR _10513_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_235_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28502_ clknet_leaf_113_clk _02300_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_235_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25714_ systolic_inst.acc_wires\[5\]\[30\] C_out\[190\] net46 VGND VGND VPWR VPWR
+ _03016_ sky130_fd_sc_hd__mux2_1
XFILLER_5_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22926_ _09603_ _09604_ VGND VGND VPWR VPWR _09605_ sky130_fd_sc_hd__nand2b_1
X_29482_ clknet_leaf_271_clk _03280_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[454\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26694_ clknet_leaf_1_B_in_serial_clk _00497_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28433_ clknet_leaf_28_clk _02231_ VGND VGND VPWR VPWR systolic_inst.A_shift\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_231_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25645_ systolic_inst.acc_wires\[3\]\[25\] C_out\[121\] net50 VGND VGND VPWR VPWR
+ _02947_ sky130_fd_sc_hd__mux2_1
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22857_ _09535_ _09536_ VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21808_ _08610_ _08611_ VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__nor2_1
X_28364_ clknet_leaf_29_clk _02162_ VGND VGND VPWR VPWR systolic_inst.A_shift\[20\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25576_ systolic_inst.acc_wires\[1\]\[20\] C_out\[52\] net53 VGND VGND VPWR VPWR
+ _02878_ sky130_fd_sc_hd__mux2_1
X_13590_ deser_B.word_buffer\[26\] deser_B.serial_word\[26\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__mux2_1
X_22788_ _09468_ _09469_ _09438_ VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__a21o_1
XFILLER_40_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27315_ clknet_leaf_290_clk _01113_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24527_ C_out\[90\] net100 net82 ser_C.shift_reg\[90\] _10733_ VGND VGND VPWR VPWR
+ _02340_ sky130_fd_sc_hd__a221o_1
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28295_ clknet_leaf_121_clk _02093_ VGND VGND VPWR VPWR systolic_inst.B_shift\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_21739_ _08473_ _08477_ _08507_ _08509_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__o31a_1
XFILLER_157_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15260_ _12355_ _12356_ VGND VGND VPWR VPWR _12358_ sky130_fd_sc_hd__nor2_1
X_27246_ clknet_leaf_274_clk _01044_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24458_ net114 ser_C.shift_reg\[57\] VGND VGND VPWR VPWR _10699_ sky130_fd_sc_hd__and2_1
XFILLER_36_1291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14211_ _11378_ _11398_ VGND VGND VPWR VPWR _11400_ sky130_fd_sc_hd__xnor2_1
X_23409_ systolic_inst.B_outs\[0\]\[3\] systolic_inst.A_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[4\]
+ systolic_inst.A_outs\[0\]\[4\] VGND VGND VPWR VPWR _10035_ sky130_fd_sc_hd__and4_1
XFILLER_138_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15191_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[14\]\[7\]
+ VGND VGND VPWR VPWR _12298_ sky130_fd_sc_hd__nand2_1
X_27177_ clknet_leaf_248_clk _00975_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_229_Right_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24389_ C_out\[21\] net104 _10643_ ser_C.shift_reg\[21\] _10664_ VGND VGND VPWR VPWR
+ _02271_ sky130_fd_sc_hd__a221o_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_9 systolic_inst.A_outs\[6\]\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26128_ deser_B.serial_word\[83\] deser_B.shift_reg\[83\] net56 VGND VGND VPWR VPWR
+ _03430_ sky130_fd_sc_hd__mux2_1
X_14142_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[1\]
+ systolic_inst.A_outs\[15\]\[0\] VGND VGND VPWR VPWR _11335_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14073_ deser_B.shift_reg\[107\] deser_B.shift_reg\[108\] net126 VGND VGND VPWR VPWR
+ _00899_ sky130_fd_sc_hd__mux2_1
X_26059_ deser_B.serial_word\[14\] deser_B.shift_reg\[14\] net55 VGND VGND VPWR VPWR
+ _03361_ sky130_fd_sc_hd__mux2_1
X_18950_ _06047_ _06048_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__and2_1
XFILLER_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_18_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17901_ _05091_ _05092_ _05094_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__or3_1
X_18881_ _05988_ _05989_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__nand2_1
XFILLER_117_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17832_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[2\] VGND VGND VPWR
+ VPWR _05029_ sky130_fd_sc_hd__and2_1
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17763_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[28\]
+ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__or2_1
X_14975_ _12070_ _12095_ VGND VGND VPWR VPWR _12096_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19502_ _06541_ _06543_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__or2_1
XFILLER_75_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16714_ _04032_ _04035_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__xnor2_1
X_13926_ deser_A.serial_word\[87\] deser_A.shift_reg\[87\] net57 VGND VGND VPWR VPWR
+ _00752_ sky130_fd_sc_hd__mux2_1
X_17694_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[16\]
+ _04922_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19433_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[7\]\[5\]
+ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__and2_1
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16645_ _03951_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__xor2_1
XFILLER_223_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13857_ deser_A.serial_word\[18\] deser_A.shift_reg\[18\] net58 VGND VGND VPWR VPWR
+ _00683_ sky130_fd_sc_hd__mux2_1
XFILLER_63_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19364_ _06374_ _06423_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16576_ systolic_inst.A_outs\[11\]\[1\] systolic_inst.A_outs\[10\]\[1\] net118 VGND
+ VGND VPWR VPWR _01203_ sky130_fd_sc_hd__mux2_1
X_13788_ B_in\[95\] deser_B.word_buffer\[95\] net89 VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__mux2_1
X_18315_ systolic_inst.acc_wires\[9\]\[16\] systolic_inst.acc_wires\[9\]\[17\] systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__o21ai_1
XFILLER_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15527_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[6\] VGND VGND
+ VPWR VPWR _12585_ sky130_fd_sc_hd__nand2_1
X_19295_ _06348_ _06356_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__nand2_1
XFILLER_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18246_ net66 _05421_ _05422_ systolic_inst.acc_wires\[9\]\[8\] net107 VGND VGND
+ VPWR VPWR _01370_ sky130_fd_sc_hd__a32o_1
XFILLER_31_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15458_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[4\] _12515_ _12516_
+ VGND VGND VPWR VPWR _12518_ sky130_fd_sc_hd__a22o_1
XFILLER_176_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14409_ _11558_ _11591_ systolic_inst.A_outs\[15\]\[7\] VGND VGND VPWR VPWR _11592_
+ sky130_fd_sc_hd__and3b_1
XFILLER_117_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18177_ _05363_ _05362_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__nand2b_1
XFILLER_239_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15389_ _12450_ _12451_ VGND VGND VPWR VPWR _12452_ sky130_fd_sc_hd__nor2_1
XFILLER_50_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_27_A_in_serial_clk clknet_2_0__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_27_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_17128_ _04396_ _04403_ _04408_ _04413_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__nand4_1
XFILLER_237_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_292_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_292_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17059_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[11\]\[12\]
+ _04355_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_111_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20070_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[6\]\[8\]
+ _07051_ _07053_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__a211o_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_12__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_12__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_174_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23760_ _11258_ systolic_inst.acc_wires\[0\]\[10\] net63 _10366_ VGND VGND VPWR VPWR
+ _01940_ sky130_fd_sc_hd__a22o_1
XFILLER_122_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20972_ systolic_inst.A_outs\[4\]\[2\] systolic_inst.B_outs\[4\]\[5\] systolic_inst.A_outs\[4\]\[6\]
+ systolic_inst.B_outs\[4\]\[1\] VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__a22o_1
XFILLER_122_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22711_ _09395_ _09396_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__and2_1
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23691_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[0\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _10308_ sky130_fd_sc_hd__a21o_1
XFILLER_26_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25430_ _11184_ systolic_inst.A_shift\[0\]\[6\] net70 VGND VGND VPWR VPWR _02792_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22642_ _09350_ _09352_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1002 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22573_ net65 _09293_ _09294_ systolic_inst.acc_wires\[2\]\[15\] net109 VGND VGND
+ VPWR VPWR _01825_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_118_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25361_ ser_C.parallel_data\[507\] net98 net78 ser_C.shift_reg\[507\] _11150_ VGND
+ VGND VPWR VPWR _02757_ sky130_fd_sc_hd__a221o_1
XFILLER_222_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27100_ clknet_leaf_7_B_in_serial_clk _00898_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_196_Left_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24312_ _10629_ systolic_inst.A_shift\[10\]\[3\] net70 VGND VGND VPWR VPWR _02229_
+ sky130_fd_sc_hd__mux2_1
X_28080_ clknet_leaf_114_clk _01878_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_21524_ _08329_ _08335_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25292_ net111 ser_C.shift_reg\[474\] VGND VGND VPWR VPWR _11116_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27031_ clknet_leaf_12_B_in_serial_clk _00829_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_194_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21455_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[30\]
+ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__or2_1
X_24243_ systolic_inst.A_shift\[19\]\[5\] A_in\[69\] net59 VGND VGND VPWR VPWR _10607_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20406_ systolic_inst.B_outs\[5\]\[7\] _07235_ _07267_ _07304_ VGND VGND VPWR VPWR
+ _07343_ sky130_fd_sc_hd__o31a_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24174_ systolic_inst.A_shift\[26\]\[5\] net70 _10505_ systolic_inst.A_shift\[27\]\[5\]
+ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__a22o_1
XFILLER_135_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21386_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[20\]
+ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_224_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_224_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23125_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[1\]\[8\]
+ _09786_ _09788_ VGND VGND VPWR VPWR _09789_ sky130_fd_sc_hd__a211o_1
X_20337_ _07273_ _07274_ _07262_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__a21o_1
X_28982_ clknet_leaf_60_clk _02780_ VGND VGND VPWR VPWR systolic_inst.A_shift\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23056_ _09728_ _09729_ VGND VGND VPWR VPWR _09731_ sky130_fd_sc_hd__xnor2_1
X_27933_ clknet_leaf_180_clk _01731_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_20268_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[2\] VGND VGND VPWR
+ VPWR _07209_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_34_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22007_ _08784_ _08786_ _08787_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__or3_1
XFILLER_114_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27864_ clknet_leaf_147_clk _01662_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_118_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20199_ systolic_inst.acc_wires\[6\]\[26\] systolic_inst.acc_wires\[6\]\[27\] systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__o21a_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29603_ clknet_leaf_20_B_in_serial_clk _03398_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_26815_ clknet_leaf_62_clk _00617_ net135 VGND VGND VPWR VPWR B_in\[87\] sky130_fd_sc_hd__dfrtp_1
X_27795_ clknet_leaf_45_clk _01593_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_29_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29534_ clknet_leaf_258_clk _03332_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[506\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26746_ clknet_leaf_51_clk _00548_ net143 VGND VGND VPWR VPWR B_in\[18\] sky130_fd_sc_hd__dfrtp_1
X_14760_ systolic_inst.A_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[1\]
+ systolic_inst.B_outs\[14\]\[0\] VGND VGND VPWR VPWR _11889_ sky130_fd_sc_hd__a22o_1
X_23958_ systolic_inst.B_shift\[11\]\[5\] _11332_ net83 systolic_inst.B_shift\[15\]\[5\]
+ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__a22o_1
XFILLER_57_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13711_ B_in\[18\] deser_B.word_buffer\[18\] net86 VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__mux2_1
X_22909_ _09586_ _09587_ VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__or2_1
X_29465_ clknet_leaf_287_clk _03263_ net136 VGND VGND VPWR VPWR C_out\[437\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26677_ clknet_leaf_11_B_in_serial_clk _00480_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_14691_ _11824_ _11844_ VGND VGND VPWR VPWR _11845_ sky130_fd_sc_hd__nor2_1
X_23889_ _10472_ _10475_ VGND VGND VPWR VPWR _10476_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28416_ clknet_leaf_69_clk _02214_ VGND VGND VPWR VPWR systolic_inst.B_shift\[23\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16430_ _03789_ _03792_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__or2_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13642_ deser_B.word_buffer\[78\] deser_B.serial_word\[78\] net123 VGND VGND VPWR
+ VPWR _00479_ sky130_fd_sc_hd__mux2_1
X_25628_ systolic_inst.acc_wires\[3\]\[8\] C_out\[104\] net48 VGND VGND VPWR VPWR
+ _02930_ sky130_fd_sc_hd__mux2_1
XFILLER_189_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29396_ clknet_leaf_237_clk _03194_ net145 VGND VGND VPWR VPWR C_out\[368\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16361_ _03737_ _03738_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__xnor2_1
X_28347_ clknet_leaf_342_clk _02145_ VGND VGND VPWR VPWR systolic_inst.A_shift\[25\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25559_ systolic_inst.acc_wires\[1\]\[3\] C_out\[35\] net36 VGND VGND VPWR VPWR _02861_
+ sky130_fd_sc_hd__mux2_1
X_13573_ deser_B.word_buffer\[9\] deser_B.serial_word\[9\] net124 VGND VGND VPWR VPWR
+ _00410_ sky130_fd_sc_hd__mux2_1
XFILLER_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18100_ _05149_ _05288_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_213_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15312_ _12400_ _12401_ VGND VGND VPWR VPWR _12402_ sky130_fd_sc_hd__or2_1
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19080_ _06146_ _06147_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__nor2_1
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28278_ clknet_leaf_130_clk _02076_ VGND VGND VPWR VPWR systolic_inst.B_shift\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16292_ _03671_ _03672_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__nand2_1
XFILLER_157_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18031_ _05220_ _05221_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__or2_1
XFILLER_184_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15243_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[14\]\[13\]
+ _12338_ VGND VGND VPWR VPWR _12343_ sky130_fd_sc_hd__a21oi_1
X_27229_ clknet_leaf_252_clk _01027_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_201_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15174_ _12274_ _12278_ _12281_ _12282_ VGND VGND VPWR VPWR _12284_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_274_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_274_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14125_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.A_outs\[14\]\[1\] net118 VGND
+ VGND VPWR VPWR _00947_ sky130_fd_sc_hd__mux2_1
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19982_ systolic_inst.B_outs\[6\]\[5\] systolic_inst.A_outs\[6\]\[7\] _06955_ _06954_
+ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__a31o_1
XFILLER_207_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14056_ deser_B.shift_reg\[90\] deser_B.shift_reg\[91\] deser_B.receiving VGND VGND
+ VPWR VPWR _00882_ sky130_fd_sc_hd__mux2_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18933_ _06034_ _06033_ systolic_inst.acc_wires\[8\]\[19\] net108 VGND VGND VPWR
+ VPWR _01445_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18864_ _05967_ _05971_ _05974_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__nand3_1
XFILLER_223_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17815_ _05011_ _05012_ net116 VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_199_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18795_ _05913_ _05916_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_199_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17746_ _04965_ _04967_ _04969_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__or3_1
X_14958_ _12075_ _12078_ VGND VGND VPWR VPWR _12079_ sky130_fd_sc_hd__xnor2_1
XFILLER_242_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13909_ deser_A.serial_word\[70\] deser_A.shift_reg\[70\] net57 VGND VGND VPWR VPWR
+ _00735_ sky130_fd_sc_hd__mux2_1
XFILLER_78_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17677_ _11712_ _04910_ _04911_ systolic_inst.acc_wires\[10\]\[14\] net105 VGND VGND
+ VPWR VPWR _01312_ sky130_fd_sc_hd__a32o_1
X_14889_ _12005_ _12011_ VGND VGND VPWR VPWR _12012_ sky130_fd_sc_hd__nor2_1
XFILLER_208_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19416_ _06461_ _06464_ _06468_ _06469_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__o211a_1
XFILLER_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16628_ _03949_ _03951_ _03933_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19347_ _06404_ _06405_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_154_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16559_ _03907_ _03906_ systolic_inst.acc_wires\[12\]\[28\] net108 VGND VGND VPWR
+ VPWR _01198_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19278_ _06340_ _06338_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[10\]
+ net105 VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_14_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18229_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[9\]\[6\]
+ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__and2_1
XFILLER_164_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21240_ _08057_ _08085_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__nand2_1
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_265_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_265_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21171_ _07884_ _08039_ systolic_inst.A_outs\[4\]\[7\] VGND VGND VPWR VPWR _08040_
+ sky130_fd_sc_hd__and3b_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20122_ _07086_ _07093_ _07094_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__o21ba_1
XFILLER_137_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20053_ _07033_ _07034_ _07032_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__a21bo_1
X_24930_ net111 ser_C.shift_reg\[293\] VGND VGND VPWR VPWR _10935_ sky130_fd_sc_hd__and2_1
XFILLER_219_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24861_ C_out\[257\] net101 net73 ser_C.shift_reg\[257\] _10900_ VGND VGND VPWR VPWR
+ _02507_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26600_ clknet_leaf_18_B_in_serial_clk _00403_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23812_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[18\]
+ VGND VGND VPWR VPWR _10411_ sky130_fd_sc_hd__nand2_1
XFILLER_6_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27580_ clknet_leaf_220_clk _01378_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24792_ net112 ser_C.shift_reg\[224\] VGND VGND VPWR VPWR _10866_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26531_ clknet_leaf_5_A_in_serial_clk _00334_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_217_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23743_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[0\]\[8\]
+ VGND VGND VPWR VPWR _10352_ sky130_fd_sc_hd__xor2_1
XFILLER_226_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20955_ _07828_ _07829_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__nor2_1
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29250_ clknet_leaf_184_clk _03048_ net146 VGND VGND VPWR VPWR C_out\[222\] sky130_fd_sc_hd__dfrtp_1
XFILLER_242_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26462_ clknet_leaf_1_A_in_serial_clk _00269_ net132 VGND VGND VPWR VPWR deser_A.bit_idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23674_ _10266_ _10272_ _10291_ VGND VGND VPWR VPWR _10293_ sky130_fd_sc_hd__or3_1
X_20886_ _07760_ _07761_ _07742_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28201_ clknet_leaf_128_clk _01999_ VGND VGND VPWR VPWR systolic_inst.B_shift\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_25413_ systolic_inst.A_shift\[2\]\[6\] A_in\[14\] net59 VGND VGND VPWR VPWR _11176_
+ sky130_fd_sc_hd__mux2_1
X_22625_ systolic_inst.acc_wires\[2\]\[20\] systolic_inst.acc_wires\[2\]\[21\] systolic_inst.acc_wires\[2\]\[22\]
+ systolic_inst.acc_wires\[2\]\[23\] systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__o41a_1
X_29181_ clknet_leaf_44_clk _02979_ net142 VGND VGND VPWR VPWR C_out\[153\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26393_ clknet_leaf_16_clk _00200_ net132 VGND VGND VPWR VPWR A_in\[61\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28132_ clknet_leaf_128_clk _01930_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25344_ net112 ser_C.shift_reg\[500\] VGND VGND VPWR VPWR _11142_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22556_ _09274_ _09278_ VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__nand2b_1
XFILLER_22_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28063_ clknet_leaf_121_clk _01861_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21507_ _08299_ _08305_ _08308_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25275_ ser_C.parallel_data\[464\] net102 net74 ser_C.shift_reg\[464\] _11107_ VGND
+ VGND VPWR VPWR _02714_ sky130_fd_sc_hd__a221o_1
X_22487_ _09214_ _09215_ _09213_ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__a21bo_1
XFILLER_181_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27014_ clknet_leaf_21_B_in_serial_clk _00812_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24226_ _10598_ systolic_inst.A_shift\[19\]\[4\] net70 VGND VGND VPWR VPWR _02174_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21438_ _11258_ systolic_inst.acc_wires\[4\]\[27\] net63 _08275_ VGND VGND VPWR VPWR
+ _01709_ sky130_fd_sc_hd__a22o_1
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_256_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_256_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21369_ _11258_ systolic_inst.acc_wires\[4\]\[16\] _08215_ _08217_ VGND VGND VPWR
+ VPWR _01698_ sky130_fd_sc_hd__a22o_1
X_24157_ systolic_inst.A_shift\[28\]\[2\] A_in\[98\] net59 VGND VGND VPWR VPWR _10580_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23108_ _09768_ _09769_ _09767_ VGND VGND VPWR VPWR _09775_ sky130_fd_sc_hd__a21bo_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28965_ clknet_leaf_78_clk _02763_ VGND VGND VPWR VPWR systolic_inst.B_shift\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_24088_ systolic_inst.B_shift\[2\]\[7\] net70 net83 systolic_inst.B_shift\[6\]\[7\]
+ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__a22o_1
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15930_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[27\]
+ VGND VGND VPWR VPWR _12953_ sky130_fd_sc_hd__xnor2_1
X_27916_ clknet_leaf_145_clk _01714_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_23039_ _11277_ systolic_inst.A_outs\[1\]\[7\] _09660_ _09686_ VGND VGND VPWR VPWR
+ _09714_ sky130_fd_sc_hd__o211ai_1
XFILLER_114_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28896_ clknet_leaf_284_clk _02694_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[444\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27847_ clknet_leaf_180_clk _01645_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_15861_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[16\]
+ VGND VGND VPWR VPWR _12895_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_202_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_202_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[10\]\[4\]
+ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__or2_1
X_14812_ _11935_ _11936_ VGND VGND VPWR VPWR _11937_ sky130_fd_sc_hd__or2_1
XFILLER_92_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18580_ _05705_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27778_ clknet_leaf_176_clk _01576_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_15792_ _12832_ _12833_ _12834_ VGND VGND VPWR VPWR _12836_ sky130_fd_sc_hd__and3_1
XFILLER_224_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17531_ _04781_ _04782_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_194_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26729_ clknet_leaf_73_clk _00531_ net144 VGND VGND VPWR VPWR B_in\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14743_ systolic_inst.A_outs\[14\]\[3\] systolic_inst.A_outs\[13\]\[3\] net116 VGND
+ VGND VPWR VPWR _01013_ sky130_fd_sc_hd__mux2_1
X_29517_ clknet_leaf_255_clk _03315_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[489\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29448_ clknet_leaf_293_clk _03246_ net139 VGND VGND VPWR VPWR C_out\[420\] sky130_fd_sc_hd__dfrtp_1
X_17462_ systolic_inst.A_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[5\] systolic_inst.B_outs\[10\]\[6\]
+ systolic_inst.B_outs\[10\]\[7\] VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__and4b_1
XFILLER_229_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14674_ _11830_ _11829_ systolic_inst.acc_wires\[15\]\[21\] net107 VGND VGND VPWR
+ VPWR _00999_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19201_ _06234_ _06264_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__xor2_1
X_16413_ _03775_ _03778_ _03780_ _03781_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__o211ai_2
X_13625_ deser_B.word_buffer\[61\] deser_B.serial_word\[61\] net123 VGND VGND VPWR
+ VPWR _00462_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29379_ clknet_leaf_244_clk _03177_ net145 VGND VGND VPWR VPWR C_out\[351\] sky130_fd_sc_hd__dfrtp_1
X_17393_ systolic_inst.A_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[6\]
+ systolic_inst.B_outs\[10\]\[7\] VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__and4b_1
XFILLER_60_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19132_ _06168_ _06191_ _06190_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__a21boi_1
XFILLER_9_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16344_ _03660_ _03722_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13556_ deser_A.shift_reg\[120\] deser_A.shift_reg\[121\] net130 VGND VGND VPWR VPWR
+ _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_80_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19063_ systolic_inst.A_outs\[7\]\[4\] _06131_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__nand2_1
XFILLER_186_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16275_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[11\] _03656_ net115
+ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__mux2_1
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13487_ deser_A.shift_reg\[51\] deser_A.shift_reg\[52\] net130 VGND VGND VPWR VPWR
+ _00324_ sky130_fd_sc_hd__mux2_1
XFILLER_218_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18014_ _05166_ _05168_ _05204_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__nand3_1
XFILLER_199_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15226_ _12314_ _12320_ _12322_ VGND VGND VPWR VPWR _12328_ sky130_fd_sc_hd__o21a_1
XFILLER_173_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_247_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_247_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_172_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15157_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[14\]\[2\]
+ VGND VGND VPWR VPWR _12269_ sky130_fd_sc_hd__nand2_1
X_14108_ systolic_inst.B_shift\[12\]\[0\] net72 _11333_ B_in\[96\] VGND VGND VPWR
+ VPWR _00930_ sky130_fd_sc_hd__a22o_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19965_ _06895_ _06959_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_147_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15088_ systolic_inst.B_outs\[14\]\[6\] systolic_inst.A_outs\[14\]\[7\] VGND VGND
+ VPWR VPWR _12205_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14039_ deser_B.shift_reg\[73\] deser_B.shift_reg\[74\] deser_B.receiving VGND VGND
+ VPWR VPWR _00865_ sky130_fd_sc_hd__mux2_1
X_18916_ net63 _06018_ _06020_ systolic_inst.acc_wires\[8\]\[16\] net108 VGND VGND
+ VPWR VPWR _01442_ sky130_fd_sc_hd__a32o_1
X_19896_ _06858_ _06893_ systolic_inst.A_outs\[6\]\[7\] VGND VGND VPWR VPWR _06894_
+ sky130_fd_sc_hd__and3b_1
X_18847_ net63 _05959_ _05960_ systolic_inst.acc_wires\[8\]\[7\] net108 VGND VGND
+ VPWR VPWR _01433_ sky130_fd_sc_hd__a32o_1
XFILLER_95_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18778_ _05899_ _05900_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__nor2_1
XFILLER_227_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17729_ _11712_ _04954_ _04955_ systolic_inst.acc_wires\[10\]\[22\] net105 VGND VGND
+ VPWR VPWR _01320_ sky130_fd_sc_hd__a32o_1
XFILLER_63_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20740_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[18\]
+ VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20671_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[5\]\[8\]
+ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__xor2_1
XFILLER_177_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22410_ _09085_ _09088_ _09118_ _09116_ VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__o31a_1
XFILLER_91_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23390_ _09968_ _10016_ VGND VGND VPWR VPWR _10017_ sky130_fd_sc_hd__or2_1
XFILLER_91_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22341_ _09020_ _09045_ _09044_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__a21boi_1
XFILLER_137_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22272_ _09016_ _09015_ VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__nand2b_1
X_25060_ net112 ser_C.shift_reg\[358\] VGND VGND VPWR VPWR _11000_ sky130_fd_sc_hd__and2_1
XFILLER_178_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24011_ systolic_inst.B_shift\[7\]\[2\] net70 net83 systolic_inst.B_shift\[11\]\[2\]
+ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21223_ systolic_inst.A_outs\[4\]\[6\] _07852_ _08060_ _08062_ VGND VGND VPWR VPWR
+ _08090_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_238_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_238_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21154_ _07982_ _07986_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__nor2_1
XFILLER_132_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20105_ _07080_ _07082_ _07084_ systolic_inst.acc_wires\[6\]\[13\] net106 VGND VGND
+ VPWR VPWR _01567_ sky130_fd_sc_hd__a32o_1
X_28750_ clknet_leaf_222_clk _02548_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[298\]
+ sky130_fd_sc_hd__dfrtp_1
X_21085_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\] systolic_inst.A_outs\[4\]\[6\]
+ systolic_inst.A_outs\[4\]\[7\] VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__nand4_1
X_25962_ systolic_inst.acc_wires\[13\]\[22\] C_out\[438\] net19 VGND VGND VPWR VPWR
+ _03264_ sky130_fd_sc_hd__mux2_1
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27701_ clknet_leaf_198_clk _01499_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20036_ net68 _07023_ _07025_ systolic_inst.acc_wires\[6\]\[3\] net106 VGND VGND
+ VPWR VPWR _01557_ sky130_fd_sc_hd__a32o_1
X_24913_ C_out\[283\] net103 net75 ser_C.shift_reg\[283\] _10926_ VGND VGND VPWR VPWR
+ _02533_ sky130_fd_sc_hd__a221o_1
XFILLER_219_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28681_ clknet_leaf_195_clk _02479_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[229\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25893_ systolic_inst.acc_wires\[11\]\[17\] C_out\[369\] net39 VGND VGND VPWR VPWR
+ _03195_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_219_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_29_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_115_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27632_ clknet_leaf_324_clk _01430_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24844_ net113 ser_C.shift_reg\[250\] VGND VGND VPWR VPWR _10892_ sky130_fd_sc_hd__and2_1
XFILLER_46_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_215_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27563_ clknet_leaf_218_clk _01361_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_73_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24775_ C_out\[214\] net98 net78 ser_C.shift_reg\[214\] _10857_ VGND VGND VPWR VPWR
+ _02464_ sky130_fd_sc_hd__a221o_1
X_21987_ _08768_ _08770_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__xnor2_1
X_29302_ clknet_leaf_325_clk _03100_ net142 VGND VGND VPWR VPWR C_out\[274\] sky130_fd_sc_hd__dfrtp_1
XFILLER_148_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26514_ clknet_leaf_11_A_in_serial_clk _00317_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_23726_ _10334_ _10335_ _10336_ VGND VGND VPWR VPWR _10338_ sky130_fd_sc_hd__and3_1
XFILLER_226_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27494_ clknet_leaf_227_clk _01292_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_20938_ _07811_ _07812_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__nand2_1
XFILLER_242_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29233_ clknet_leaf_204_clk _03031_ net147 VGND VGND VPWR VPWR C_out\[205\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26445_ clknet_leaf_348_clk _00252_ net132 VGND VGND VPWR VPWR A_in\[113\] sky130_fd_sc_hd__dfrtp_1
X_23657_ _10274_ _10275_ _10224_ _10227_ VGND VGND VPWR VPWR _10277_ sky130_fd_sc_hd__o211a_1
XFILLER_35_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20869_ _07739_ _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__xnor2_1
XFILLER_224_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13410_ A_in\[119\] deser_A.word_buffer\[119\] net92 VGND VGND VPWR VPWR _00258_
+ sky130_fd_sc_hd__mux2_1
X_22608_ _09322_ _09323_ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__xor2_1
XFILLER_169_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29164_ clknet_leaf_39_clk _02962_ net142 VGND VGND VPWR VPWR C_out\[136\] sky130_fd_sc_hd__dfrtp_1
XFILLER_179_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14390_ _11521_ _11522_ _11539_ _11538_ _11537_ VGND VGND VPWR VPWR _11574_ sky130_fd_sc_hd__o32a_1
X_26376_ clknet_leaf_28_clk _00183_ net133 VGND VGND VPWR VPWR A_in\[44\] sky130_fd_sc_hd__dfrtp_1
XFILLER_195_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23588_ _10208_ _10209_ VGND VGND VPWR VPWR _10210_ sky130_fd_sc_hd__nor2_1
XFILLER_10_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28115_ clknet_leaf_47_clk _01913_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_128_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25327_ ser_C.parallel_data\[490\] net97 net77 ser_C.shift_reg\[490\] _11133_ VGND
+ VGND VPWR VPWR _02740_ sky130_fd_sc_hd__a221o_1
XFILLER_70_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13341_ A_in\[50\] deser_A.word_buffer\[50\] net92 VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__mux2_1
X_29095_ clknet_leaf_155_clk _02893_ net150 VGND VGND VPWR VPWR C_out\[67\] sky130_fd_sc_hd__dfrtp_1
X_22539_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[2\]\[11\]
+ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__or2_1
XFILLER_183_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28046_ clknet_leaf_127_clk _01844_ net144 VGND VGND VPWR VPWR systolic_inst.A_outs\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_16060_ systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[5\] systolic_inst.A_outs\[12\]\[6\]
+ systolic_inst.B_outs\[12\]\[0\] VGND VGND VPWR VPWR _13056_ sky130_fd_sc_hd__a22oi_1
XFILLER_143_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25258_ net111 ser_C.shift_reg\[457\] VGND VGND VPWR VPWR _11099_ sky130_fd_sc_hd__and2_1
X_13272_ deser_A.word_buffer\[110\] deser_A.serial_word\[110\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__mux2_1
XFILLER_108_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15011_ _12072_ _12129_ VGND VGND VPWR VPWR _12131_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_229_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_229_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_237_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24209_ systolic_inst.A_shift\[21\]\[4\] A_in\[84\] net59 VGND VGND VPWR VPWR _10590_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25189_ C_out\[421\] net102 net74 ser_C.shift_reg\[421\] _11064_ VGND VGND VPWR VPWR
+ _02671_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_204_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_204_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19750_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[5\] VGND VGND VPWR
+ VPWR _06752_ sky130_fd_sc_hd__nand2_1
XFILLER_68_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28948_ clknet_leaf_260_clk _02746_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[496\]
+ sky130_fd_sc_hd__dfrtp_1
X_16962_ _04056_ _04196_ _04267_ _04265_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__a31o_1
XFILLER_111_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18701_ _05787_ _05789_ _05824_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__a21oi_1
X_15913_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[24\]
+ VGND VGND VPWR VPWR _12939_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_196_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19681_ _06663_ _06665_ _06664_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__a21bo_1
XFILLER_49_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16893_ _04176_ _04178_ _04209_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__a21o_1
XFILLER_103_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_196_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28879_ clknet_leaf_289_clk _02677_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[427\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_1349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15844_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[13\]\[14\]
+ VGND VGND VPWR VPWR _12880_ sky130_fd_sc_hd__nand2_1
XFILLER_65_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18632_ _05757_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__nand2_1
XFILLER_225_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15775_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[13\]\[4\]
+ VGND VGND VPWR VPWR _12821_ sky130_fd_sc_hd__or2_1
X_18563_ systolic_inst.B_outs\[8\]\[7\] _05658_ _05659_ VGND VGND VPWR VPWR _05692_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_224_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14726_ _11872_ _11874_ VGND VGND VPWR VPWR _11875_ sky130_fd_sc_hd__xnor2_1
X_17514_ _04701_ _04705_ _04735_ _04734_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__o31a_1
X_18494_ systolic_inst.A_outs\[8\]\[4\] _05587_ _05605_ _05604_ _05601_ VGND VGND
+ VPWR VPWR _05625_ sky130_fd_sc_hd__a32o_1
XFILLER_91_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17445_ _04638_ _04663_ _04662_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__a21boi_1
X_14657_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[19\]
+ VGND VGND VPWR VPWR _11816_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13608_ deser_B.word_buffer\[44\] deser_B.serial_word\[44\] net124 VGND VGND VPWR
+ VPWR _00445_ sky130_fd_sc_hd__mux2_1
XFILLER_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17376_ _04630_ _04631_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__xor2_1
X_14588_ _11752_ _11754_ VGND VGND VPWR VPWR _11757_ sky130_fd_sc_hd__nand2_1
XFILLER_220_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19115_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.A_outs\[7\]\[1\] systolic_inst.B_outs\[7\]\[5\]
+ systolic_inst.B_outs\[7\]\[6\] VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__and4_1
XFILLER_14_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16327_ _03705_ _03706_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__nor2_1
XFILLER_158_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13539_ deser_A.shift_reg\[103\] deser_A.shift_reg\[104\] net129 VGND VGND VPWR VPWR
+ _00376_ sky130_fd_sc_hd__mux2_1
XFILLER_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19046_ systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[3\]
+ systolic_inst.B_outs\[7\]\[0\] VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__a22o_1
XFILLER_12_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16258_ _03637_ _03638_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_149_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15209_ _12309_ _12311_ _12313_ systolic_inst.acc_wires\[14\]\[9\] net107 VGND VGND
+ VPWR VPWR _01051_ sky130_fd_sc_hd__a32o_1
XFILLER_133_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16189_ _03564_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19948_ _06942_ _06943_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19879_ _06875_ _06876_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21910_ _08704_ VGND VGND VPWR VPWR _08705_ sky130_fd_sc_hd__inv_2
XFILLER_110_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22890_ _09561_ _09569_ VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21841_ _08556_ _08642_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__and2_1
XFILLER_93_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24560_ net113 ser_C.shift_reg\[108\] VGND VGND VPWR VPWR _10750_ sky130_fd_sc_hd__and2_1
XFILLER_130_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21772_ _08575_ _08577_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__nor2_1
XFILLER_230_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23511_ _10132_ _10133_ _10089_ _10092_ VGND VGND VPWR VPWR _10135_ sky130_fd_sc_hd__o211ai_2
X_20723_ _07634_ _07635_ _07628_ _07632_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__o211ai_1
X_24491_ C_out\[72\] _11302_ net81 ser_C.shift_reg\[72\] _10715_ VGND VGND VPWR VPWR
+ _02322_ sky130_fd_sc_hd__a221o_1
XFILLER_184_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26230_ clknet_leaf_7_A_in_serial_clk _00038_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23442_ systolic_inst.A_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[5\] _10025_ VGND
+ VGND VPWR VPWR _10067_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20654_ _07574_ _07575_ _07576_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__and3_1
XFILLER_17_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26161_ deser_B.serial_word\[116\] deser_B.shift_reg\[116\] net56 VGND VGND VPWR
+ VPWR _03463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20585_ _07487_ _07491_ _07516_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__or3_1
X_23373_ systolic_inst.B_outs\[0\]\[3\] systolic_inst.A_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[4\]
+ systolic_inst.A_outs\[0\]\[2\] VGND VGND VPWR VPWR _10000_ sky130_fd_sc_hd__a22oi_1
XFILLER_149_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25112_ net110 ser_C.shift_reg\[384\] VGND VGND VPWR VPWR _11026_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_95_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22324_ _09063_ _09066_ VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26092_ deser_B.serial_word\[47\] deser_B.shift_reg\[47\] net55 VGND VGND VPWR VPWR
+ _03394_ sky130_fd_sc_hd__mux2_1
XFILLER_165_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25043_ C_out\[348\] net98 net78 ser_C.shift_reg\[348\] _10991_ VGND VGND VPWR VPWR
+ _02598_ sky130_fd_sc_hd__a221o_1
X_22255_ systolic_inst.A_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[5\] _08963_ _08962_
+ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__a31oi_2
XFILLER_219_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21206_ _07991_ _08072_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_240_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22186_ _08903_ _08931_ _08932_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__and3_1
XFILLER_132_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_240_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28802_ clknet_leaf_244_clk _02600_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[350\]
+ sky130_fd_sc_hd__dfrtp_1
X_21137_ systolic_inst.A_outs\[4\]\[4\] systolic_inst.B_outs\[4\]\[6\] _07964_ _07965_
+ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__a31o_1
XFILLER_238_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26994_ clknet_leaf_1_A_in_serial_clk _00792_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_132_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21068_ _07922_ _07938_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__and2_1
X_25945_ systolic_inst.acc_wires\[13\]\[5\] C_out\[421\] net26 VGND VGND VPWR VPWR
+ _03247_ sky130_fd_sc_hd__mux2_1
X_28733_ clknet_leaf_302_clk _02531_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20019_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[6\]\[0\]
+ _07009_ _07010_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__and4_1
XFILLER_115_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28664_ clknet_leaf_176_clk _02462_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[212\]
+ sky130_fd_sc_hd__dfrtp_1
X_25876_ systolic_inst.acc_wires\[11\]\[0\] C_out\[352\] net39 VGND VGND VPWR VPWR
+ _03178_ sky130_fd_sc_hd__mux2_1
X_13890_ deser_A.serial_word\[51\] deser_A.shift_reg\[51\] net58 VGND VGND VPWR VPWR
+ _00716_ sky130_fd_sc_hd__mux2_1
XFILLER_235_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_238_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24827_ C_out\[240\] net99 net79 ser_C.shift_reg\[240\] _10883_ VGND VGND VPWR VPWR
+ _02490_ sky130_fd_sc_hd__a221o_1
X_27615_ clknet_leaf_324_clk _01413_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_238_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28595_ clknet_leaf_43_clk _02393_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[143\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15560_ systolic_inst.B_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[5\] systolic_inst.A_outs\[13\]\[6\]
+ systolic_inst.B_outs\[13\]\[3\] VGND VGND VPWR VPWR _12617_ sky130_fd_sc_hd__a22oi_1
X_27546_ clknet_leaf_34_clk _01344_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_199_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24758_ net113 ser_C.shift_reg\[207\] VGND VGND VPWR VPWR _10849_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14511_ _11620_ _11669_ _11667_ VGND VGND VPWR VPWR _11691_ sky130_fd_sc_hd__a21oi_1
X_23709_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[0\]\[3\]
+ VGND VGND VPWR VPWR _10323_ sky130_fd_sc_hd__or2_1
XFILLER_226_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27477_ clknet_leaf_307_clk _01275_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_15491_ _12548_ _12549_ VGND VGND VPWR VPWR _12550_ sky130_fd_sc_hd__or2_1
X_24689_ C_out\[171\] net104 net76 ser_C.shift_reg\[171\] _10814_ VGND VGND VPWR VPWR
+ _02421_ sky130_fd_sc_hd__a221o_1
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17230_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[3\]
+ systolic_inst.A_outs\[10\]\[4\] VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__and4_1
X_29216_ clknet_leaf_179_clk _03014_ net148 VGND VGND VPWR VPWR C_out\[188\] sky130_fd_sc_hd__dfrtp_1
X_26428_ clknet_leaf_3_clk _00235_ net131 VGND VGND VPWR VPWR A_in\[96\] sky130_fd_sc_hd__dfrtp_1
X_14442_ systolic_inst.A_outs\[15\]\[5\] systolic_inst.B_outs\[15\]\[6\] systolic_inst.A_outs\[15\]\[6\]
+ systolic_inst.B_outs\[15\]\[7\] VGND VGND VPWR VPWR _11624_ sky130_fd_sc_hd__and4b_1
XFILLER_187_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_189_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29147_ clknet_leaf_175_clk _02945_ net150 VGND VGND VPWR VPWR C_out\[119\] sky130_fd_sc_hd__dfrtp_1
XFILLER_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17161_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[29\]
+ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_189_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26359_ clknet_leaf_66_clk _00166_ net134 VGND VGND VPWR VPWR A_in\[27\] sky130_fd_sc_hd__dfrtp_1
X_14373_ systolic_inst.B_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[6\] systolic_inst.A_outs\[15\]\[7\]
+ systolic_inst.B_outs\[15\]\[3\] VGND VGND VPWR VPWR _11557_ sky130_fd_sc_hd__a22o_1
XFILLER_183_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16112_ _13099_ _03496_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__xnor2_1
X_13324_ A_in\[33\] deser_A.word_buffer\[33\] net94 VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__mux2_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29078_ clknet_leaf_113_clk _02876_ net150 VGND VGND VPWR VPWR C_out\[50\] sky130_fd_sc_hd__dfrtp_1
XFILLER_196_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17092_ _04385_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__nand2_1
XFILLER_155_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28029_ clknet_leaf_161_clk _01827_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_202_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16043_ _13036_ _13039_ VGND VGND VPWR VPWR _13040_ sky130_fd_sc_hd__xnor2_1
X_13255_ deser_A.word_buffer\[93\] deser_A.serial_word\[93\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13186_ deser_A.word_buffer\[24\] deser_A.serial_word\[24\] net128 VGND VGND VPWR
+ VPWR _00034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19802_ _06727_ _06761_ _06763_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17994_ _05147_ _05153_ _05152_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__a21o_1
XFILLER_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19733_ _06704_ _06707_ _06734_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__a211oi_2
XFILLER_133_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16945_ _04234_ _04236_ _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__a21oi_1
X_19664_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.A_outs\[6\]\[4\] VGND VGND VPWR
+ VPWR _06669_ sky130_fd_sc_hd__nand2_1
X_16876_ _04155_ _04161_ _04192_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__o21ai_1
XFILLER_231_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18615_ _05741_ _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__nor2_1
XFILLER_168_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15827_ _12855_ _12860_ _12861_ VGND VGND VPWR VPWR _12865_ sky130_fd_sc_hd__nand3_1
XFILLER_25_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19595_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[29\]
+ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__xor2_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15758_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[13\]\[0\]
+ _12803_ _12804_ VGND VGND VPWR VPWR _12807_ sky130_fd_sc_hd__a22o_1
X_18546_ _05669_ _05675_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__nor2_1
XFILLER_33_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14709_ net105 systolic_inst.acc_wires\[15\]\[26\] net69 _11860_ VGND VGND VPWR VPWR
+ _01004_ sky130_fd_sc_hd__a22o_1
XFILLER_127_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15689_ _12741_ _12742_ VGND VGND VPWR VPWR _12743_ sky130_fd_sc_hd__nand2_1
X_18477_ systolic_inst.A_outs\[8\]\[2\] systolic_inst.B_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\]
+ systolic_inst.A_outs\[8\]\[1\] VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17428_ _04679_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17359_ _04612_ _04615_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload310 clknet_leaf_120_clk VGND VGND VPWR VPWR clkload310/Y sky130_fd_sc_hd__inv_6
XFILLER_179_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20370_ _07294_ _07306_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__nand2_1
Xclkload321 clknet_leaf_156_clk VGND VGND VPWR VPWR clkload321/Y sky130_fd_sc_hd__inv_8
XFILLER_88_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload332 clknet_leaf_160_clk VGND VGND VPWR VPWR clkload332/Y sky130_fd_sc_hd__inv_6
XFILLER_88_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload40 clknet_leaf_339_clk VGND VGND VPWR VPWR clkload40/Y sky130_fd_sc_hd__bufinv_16
Xclkload343 clknet_leaf_27_A_in_serial_clk VGND VGND VPWR VPWR clkload343/X sky130_fd_sc_hd__clkbuf_8
XFILLER_238_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19029_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.A_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\]
+ systolic_inst.A_outs\[7\]\[1\] VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__and4_1
Xclkload51 clknet_leaf_301_clk VGND VGND VPWR VPWR clkload51/Y sky130_fd_sc_hd__inv_8
Xclkload354 clknet_leaf_5_A_in_serial_clk VGND VGND VPWR VPWR clkload354/Y sky130_fd_sc_hd__clkinv_2
Xclkload62 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload62/Y sky130_fd_sc_hd__inv_6
Xclkload365 clknet_leaf_18_A_in_serial_clk VGND VGND VPWR VPWR clkload365/Y sky130_fd_sc_hd__inv_8
Xclkload376 clknet_leaf_30_B_in_serial_clk VGND VGND VPWR VPWR clkload376/Y sky130_fd_sc_hd__inv_6
Xclkload73 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload73/Y sky130_fd_sc_hd__inv_6
X_22040_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[26\]
+ VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__nand2_1
Xclkload387 clknet_leaf_7_B_in_serial_clk VGND VGND VPWR VPWR clkload387/Y sky130_fd_sc_hd__bufinv_16
Xclkload84 clknet_leaf_30_clk VGND VGND VPWR VPWR clkload84/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_90_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload95 clknet_leaf_139_clk VGND VGND VPWR VPWR clkload95/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_8_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1087 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23991_ systolic_inst.B_shift\[12\]\[7\] B_in\[71\] _00008_ VGND VGND VPWR VPWR _10521_
+ sky130_fd_sc_hd__mux2_1
XFILLER_130_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25730_ systolic_inst.acc_wires\[6\]\[14\] C_out\[206\] net45 VGND VGND VPWR VPWR
+ _03032_ sky130_fd_sc_hd__mux2_1
X_22942_ _09620_ _09618_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[10\]
+ net109 VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_151_1374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25661_ systolic_inst.acc_wires\[4\]\[9\] C_out\[137\] net29 VGND VGND VPWR VPWR
+ _02963_ sky130_fd_sc_hd__mux2_1
X_22873_ _09480_ _09522_ _09521_ VGND VGND VPWR VPWR _09553_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_30_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27400_ clknet_leaf_334_clk _01198_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24612_ net110 ser_C.shift_reg\[134\] VGND VGND VPWR VPWR _10776_ sky130_fd_sc_hd__and2_1
XFILLER_231_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21824_ _08625_ _08626_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__xor2_1
XFILLER_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28380_ clknet_leaf_31_clk _02178_ VGND VGND VPWR VPWR systolic_inst.A_shift\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25592_ systolic_inst.acc_wires\[2\]\[4\] C_out\[68\] net34 VGND VGND VPWR VPWR _02894_
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_233_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27331_ clknet_leaf_288_clk _01129_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_233_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24543_ C_out\[98\] net99 net79 ser_C.shift_reg\[98\] _10741_ VGND VGND VPWR VPWR
+ _02348_ sky130_fd_sc_hd__a221o_1
XFILLER_180_1003 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21755_ _08557_ _08560_ VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__xnor2_1
X_20706_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[5\]\[12\]
+ _07619_ _07621_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__a211o_1
X_27262_ clknet_leaf_270_clk _01060_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_24474_ net112 ser_C.shift_reg\[65\] VGND VGND VPWR VPWR _10707_ sky130_fd_sc_hd__and2_1
XFILLER_157_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21686_ _08490_ _08493_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29001_ clknet_leaf_93_clk _02799_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_200_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26213_ clknet_leaf_13_A_in_serial_clk _00021_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23425_ _10048_ _10049_ VGND VGND VPWR VPWR _10051_ sky130_fd_sc_hd__xor2_1
Xclkload1 clknet_5_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_12
XFILLER_149_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20637_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[5\]\[3\]
+ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__or2_1
X_27193_ clknet_leaf_254_clk _00991_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26144_ deser_B.serial_word\[99\] deser_B.shift_reg\[99\] _00001_ VGND VGND VPWR
+ VPWR _03446_ sky130_fd_sc_hd__mux2_1
XFILLER_165_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23356_ _09982_ _09983_ VGND VGND VPWR VPWR _09984_ sky130_fd_sc_hd__nand2b_1
XFILLER_166_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20568_ _07467_ _07470_ _07498_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__or3_1
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_242_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22307_ _09013_ _09014_ _09017_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__o21a_1
XFILLER_153_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26075_ deser_B.serial_word\[30\] deser_B.shift_reg\[30\] net55 VGND VGND VPWR VPWR
+ _03377_ sky130_fd_sc_hd__mux2_1
X_23287_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[1\]
+ systolic_inst.A_outs\[0\]\[1\] VGND VGND VPWR VPWR _09919_ sky130_fd_sc_hd__and4_1
X_20499_ systolic_inst.B_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\] VGND VGND VPWR
+ VPWR _07433_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_180_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25026_ net112 ser_C.shift_reg\[341\] VGND VGND VPWR VPWR _10983_ sky130_fd_sc_hd__and2_1
XFILLER_69_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22238_ _08955_ _08957_ _08956_ VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_180_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22169_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[3\] _08900_ _08898_
+ VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_37_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14991_ _12075_ _12110_ VGND VGND VPWR VPWR _12111_ sky130_fd_sc_hd__xor2_1
X_26977_ clknet_leaf_28_A_in_serial_clk _00775_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13942_ deser_A.serial_word\[103\] deser_A.shift_reg\[103\] net57 VGND VGND VPWR
+ VPWR _00768_ sky130_fd_sc_hd__mux2_1
X_28716_ clknet_leaf_314_clk _02514_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[264\]
+ sky130_fd_sc_hd__dfrtp_1
X_16730_ _04050_ _04051_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__xor2_1
X_25928_ systolic_inst.acc_wires\[12\]\[20\] C_out\[404\] net17 VGND VGND VPWR VPWR
+ _03230_ sky130_fd_sc_hd__mux2_1
X_29696_ clknet_leaf_11_clk _03491_ VGND VGND VPWR VPWR systolic_inst.A_shift\[30\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16661_ _03983_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__nand2_1
X_28647_ clknet_leaf_202_clk _02445_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[195\]
+ sky130_fd_sc_hd__dfrtp_1
X_25859_ systolic_inst.acc_wires\[10\]\[15\] C_out\[335\] net12 VGND VGND VPWR VPWR
+ _03161_ sky130_fd_sc_hd__mux2_1
XFILLER_35_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13873_ deser_A.serial_word\[34\] deser_A.shift_reg\[34\] net58 VGND VGND VPWR VPWR
+ _00699_ sky130_fd_sc_hd__mux2_1
XFILLER_234_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18400_ _05548_ _05552_ _05553_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__a21oi_1
X_15612_ _12665_ _12666_ VGND VGND VPWR VPWR _12668_ sky130_fd_sc_hd__xnor2_1
X_19380_ _06437_ _06438_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__nor2_1
X_16592_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[0\] _03920_
+ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__a21o_1
XFILLER_222_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28578_ clknet_leaf_169_clk _02376_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_234_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18331_ _05491_ _05494_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__or3_1
X_15543_ _12600_ _12599_ VGND VGND VPWR VPWR _12601_ sky130_fd_sc_hd__and2b_1
XFILLER_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27529_ clknet_leaf_240_clk _01327_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18262_ _05434_ _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__nand2_1
X_15474_ _12531_ _12532_ _12499_ _12501_ VGND VGND VPWR VPWR _12534_ sky130_fd_sc_hd__o211a_1
X_14425_ _11590_ _11607_ VGND VGND VPWR VPWR _11608_ sky130_fd_sc_hd__xor2_1
X_17213_ systolic_inst.B_outs\[10\]\[2\] _04474_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__and2_1
XFILLER_202_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18193_ net116 _05376_ _05377_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17144_ _04429_ _04430_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__nand2_1
XFILLER_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14356_ _11498_ _11500_ _11540_ VGND VGND VPWR VPWR _11541_ sky130_fd_sc_hd__o21ai_1
XFILLER_204_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13307_ A_in\[16\] deser_A.word_buffer\[16\] net93 VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__mux2_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17075_ _04362_ _04367_ _04371_ net60 VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__a31o_1
X_14287_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[7\] _11473_ net118
+ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__mux2_1
XFILLER_226_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16026_ net108 _13022_ _13023_ VGND VGND VPWR VPWR _13024_ sky130_fd_sc_hd__or3_1
X_13238_ deser_A.word_buffer\[76\] deser_A.serial_word\[76\] net127 VGND VGND VPWR
+ VPWR _00086_ sky130_fd_sc_hd__mux2_1
XFILLER_112_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13169_ deser_A.word_buffer\[7\] deser_A.serial_word\[7\] net127 VGND VGND VPWR VPWR
+ _00017_ sky130_fd_sc_hd__mux2_1
XFILLER_174_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17977_ _05094_ _05128_ _05130_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19716_ _06717_ _06718_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__or2_1
XFILLER_133_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16928_ _04243_ _04242_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__and2b_1
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19647_ systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[3\] VGND VGND VPWR
+ VPWR _06653_ sky130_fd_sc_hd__nand2_1
X_16859_ _04174_ _04175_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19578_ _06607_ _06608_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__nand2_1
XFILLER_20_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18529_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[6\]
+ systolic_inst.A_outs\[8\]\[7\] VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__nand4_1
XFILLER_209_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21540_ _08331_ _08351_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__nand2_1
XFILLER_181_1356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21471_ systolic_inst.A_outs\[3\]\[7\] systolic_inst.A_outs\[2\]\[7\] net122 VGND
+ VGND VPWR VPWR _01721_ sky130_fd_sc_hd__mux2_1
XFILLER_53_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23210_ _09861_ VGND VGND VPWR VPWR _09862_ sky130_fd_sc_hd__inv_2
XFILLER_147_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20422_ net120 _07356_ _07357_ _07358_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__a31o_1
XFILLER_119_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24190_ systolic_inst.A_shift\[24\]\[5\] net70 _10505_ systolic_inst.A_shift\[25\]\[5\]
+ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__a22o_1
XFILLER_222_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23141_ _09801_ _09802_ VGND VGND VPWR VPWR _09803_ sky130_fd_sc_hd__nand2_1
Xclkload140 clknet_leaf_255_clk VGND VGND VPWR VPWR clkload140/Y sky130_fd_sc_hd__inv_6
XFILLER_106_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20353_ _07286_ _07290_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_77_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload151 clknet_leaf_299_clk VGND VGND VPWR VPWR clkload151/X sky130_fd_sc_hd__clkbuf_8
XFILLER_179_1296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload162 clknet_leaf_223_clk VGND VGND VPWR VPWR clkload162/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload173 clknet_leaf_249_clk VGND VGND VPWR VPWR clkload173/Y sky130_fd_sc_hd__inv_6
Xclkload184 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload184/Y sky130_fd_sc_hd__clkinv_2
X_23072_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[1\]\[1\]
+ VGND VGND VPWR VPWR _09744_ sky130_fd_sc_hd__nand2_1
Xclkload195 clknet_leaf_54_clk VGND VGND VPWR VPWR clkload195/Y sky130_fd_sc_hd__clkinvlp_4
X_20284_ _07222_ _07223_ _07201_ _07204_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_129_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22023_ _08796_ _08798_ _08795_ VGND VGND VPWR VPWR _08801_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_129_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26900_ clknet_leaf_15_A_in_serial_clk _00698_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_27880_ clknet_leaf_37_clk _01678_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26831_ clknet_leaf_87_clk _00633_ net153 VGND VGND VPWR VPWR B_in\[103\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26762_ clknet_leaf_77_clk _00564_ net143 VGND VGND VPWR VPWR B_in\[34\] sky130_fd_sc_hd__dfrtp_1
X_29550_ clknet_leaf_229_clk _03345_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_86_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23974_ _10512_ systolic_inst.B_shift\[9\]\[6\] _11332_ VGND VGND VPWR VPWR _02008_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28501_ clknet_leaf_112_clk _02299_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_25713_ systolic_inst.acc_wires\[5\]\[29\] C_out\[189\] net46 VGND VGND VPWR VPWR
+ _03015_ sky130_fd_sc_hd__mux2_1
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_235_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22925_ _09561_ _09569_ _09568_ VGND VGND VPWR VPWR _09604_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_235_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26693_ clknet_leaf_1_B_in_serial_clk _00496_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29481_ clknet_leaf_271_clk _03279_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25644_ systolic_inst.acc_wires\[3\]\[24\] C_out\[120\] net50 VGND VGND VPWR VPWR
+ _02946_ sky130_fd_sc_hd__mux2_1
X_28432_ clknet_leaf_27_clk _02230_ VGND VGND VPWR VPWR systolic_inst.A_shift\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_232_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22856_ _09535_ _09536_ VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__or2_1
XFILLER_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21807_ _08544_ _08548_ _08577_ _08610_ _08576_ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__o311a_1
X_28363_ clknet_leaf_62_clk _02161_ VGND VGND VPWR VPWR systolic_inst.B_shift\[22\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25575_ systolic_inst.acc_wires\[1\]\[19\] C_out\[51\] net35 VGND VGND VPWR VPWR
+ _02877_ sky130_fd_sc_hd__mux2_1
XFILLER_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22787_ _09438_ _09468_ _09469_ VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__nand3_1
XFILLER_40_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27314_ clknet_leaf_290_clk _01112_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24526_ net114 ser_C.shift_reg\[91\] VGND VGND VPWR VPWR _10733_ sky130_fd_sc_hd__and2_1
XFILLER_197_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28294_ clknet_leaf_101_clk _02092_ VGND VGND VPWR VPWR systolic_inst.B_shift\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_21738_ _08542_ _08543_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__xor2_1
XFILLER_240_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27245_ clknet_leaf_274_clk _01043_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24457_ C_out\[55\] net100 net82 ser_C.shift_reg\[55\] _10698_ VGND VGND VPWR VPWR
+ _02305_ sky130_fd_sc_hd__a221o_1
X_21669_ _08475_ _08476_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__and2b_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14210_ _11378_ _11398_ VGND VGND VPWR VPWR _11399_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_193_Right_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23408_ systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[6\] VGND VGND VPWR
+ VPWR _10034_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15190_ _11712_ _12295_ _12297_ systolic_inst.acc_wires\[14\]\[6\] net107 VGND VGND
+ VPWR VPWR _01048_ sky130_fd_sc_hd__a32o_1
X_27176_ clknet_leaf_248_clk _00974_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24388_ net7 ser_C.shift_reg\[22\] VGND VGND VPWR VPWR _10664_ sky130_fd_sc_hd__and2_1
XFILLER_123_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26127_ deser_B.serial_word\[82\] deser_B.shift_reg\[82\] net56 VGND VGND VPWR VPWR
+ _03429_ sky130_fd_sc_hd__mux2_1
X_14141_ net107 systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[0\] _11334_
+ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23339_ systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[5\]
+ systolic_inst.B_outs\[0\]\[0\] VGND VGND VPWR VPWR _09967_ sky130_fd_sc_hd__a22o_1
XFILLER_10_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14072_ deser_B.shift_reg\[106\] deser_B.shift_reg\[107\] net126 VGND VGND VPWR VPWR
+ _00898_ sky130_fd_sc_hd__mux2_1
X_26058_ deser_B.serial_word\[13\] deser_B.shift_reg\[13\] net55 VGND VGND VPWR VPWR
+ _03360_ sky130_fd_sc_hd__mux2_1
XFILLER_180_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17900_ _05092_ _05094_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__nor2_1
X_25009_ C_out\[331\] net97 net80 ser_C.shift_reg\[331\] _10974_ VGND VGND VPWR VPWR
+ _02581_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_14_A_in_serial_clk clknet_2_3__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_14_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_79_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18880_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[8\]\[12\]
+ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__nand2_1
XFILLER_133_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17831_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[3\] _05028_ net116
+ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__mux2_1
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17762_ _04967_ _04969_ _04981_ _04982_ _04975_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__a311oi_4
XFILLER_187_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14974_ _12092_ _12093_ VGND VGND VPWR VPWR _12095_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19501_ _06541_ _06543_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__nand2_1
X_16713_ _04000_ _04033_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13925_ deser_A.serial_word\[86\] deser_A.shift_reg\[86\] net57 VGND VGND VPWR VPWR
+ _00751_ sky130_fd_sc_hd__mux2_1
XFILLER_208_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29679_ clknet_leaf_0_B_in_serial_clk _03474_ net134 VGND VGND VPWR VPWR deser_B.serial_word\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_17693_ _04924_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__inv_2
XFILLER_207_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19432_ net62 _06482_ _06484_ systolic_inst.acc_wires\[7\]\[4\] net105 VGND VGND
+ VPWR VPWR _01494_ sky130_fd_sc_hd__a32o_1
XFILLER_228_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13856_ deser_A.serial_word\[17\] deser_A.shift_reg\[17\] net58 VGND VGND VPWR VPWR
+ _00682_ sky130_fd_sc_hd__mux2_1
XFILLER_63_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16644_ _03964_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__xor2_1
XFILLER_90_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19363_ _06421_ _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__nor2_1
XFILLER_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13787_ B_in\[94\] deser_B.word_buffer\[94\] net89 VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__mux2_1
XFILLER_76_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16575_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.A_outs\[10\]\[0\] net118 VGND
+ VGND VPWR VPWR _01202_ sky130_fd_sc_hd__mux2_1
XFILLER_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18314_ _05479_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__nand2_1
X_15526_ _12582_ _12583_ VGND VGND VPWR VPWR _12584_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _06353_ _06354_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15457_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[4\] _12515_ _12516_
+ VGND VGND VPWR VPWR _12517_ sky130_fd_sc_hd__nand4_2
XFILLER_54_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18245_ _05414_ _05417_ _05420_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_152_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14408_ systolic_inst.B_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\] VGND VGND
+ VPWR VPWR _11591_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_152_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15388_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.A_outs\[13\]\[1\] systolic_inst.B_outs\[13\]\[2\]
+ systolic_inst.B_outs\[13\]\[3\] VGND VGND VPWR VPWR _12451_ sky130_fd_sc_hd__and4_1
X_18176_ _05290_ _05338_ _05337_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__o21ba_1
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17127_ net62 _04415_ _04416_ systolic_inst.acc_wires\[11\]\[23\] net105 VGND VGND
+ VPWR VPWR _01257_ sky130_fd_sc_hd__a32o_1
XFILLER_116_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14339_ systolic_inst.B_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[5\] systolic_inst.A_outs\[15\]\[6\]
+ systolic_inst.B_outs\[15\]\[3\] VGND VGND VPWR VPWR _11524_ sky130_fd_sc_hd__a22oi_1
XFILLER_237_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17058_ _04349_ _04350_ _04357_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a21o_1
XFILLER_104_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16009_ _13005_ _13006_ VGND VGND VPWR VPWR _13007_ sky130_fd_sc_hd__nand2_1
XFILLER_217_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20971_ systolic_inst.B_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[6\]
+ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__and3_1
X_22710_ _09393_ _09394_ _09384_ VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__a21o_1
XFILLER_54_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23690_ _10307_ _10302_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ _11258_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22641_ _09343_ _09345_ _09351_ VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__a21o_1
XFILLER_20_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25360_ net112 ser_C.shift_reg\[508\] VGND VGND VPWR VPWR _11150_ sky130_fd_sc_hd__and2_1
X_22572_ _09291_ _09292_ _09285_ _09290_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__o211ai_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24311_ systolic_inst.A_shift\[11\]\[3\] A_in\[43\] net59 VGND VGND VPWR VPWR _10629_
+ sky130_fd_sc_hd__mux2_1
XFILLER_221_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21523_ _08329_ _08335_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__nor2_1
XFILLER_107_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25291_ ser_C.parallel_data\[472\] net102 net74 ser_C.shift_reg\[472\] _11115_ VGND
+ VGND VPWR VPWR _02722_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27030_ clknet_leaf_12_B_in_serial_clk _00828_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24242_ _10606_ systolic_inst.A_shift\[18\]\[4\] net70 VGND VGND VPWR VPWR _02182_
+ sky130_fd_sc_hd__mux2_1
X_21454_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[30\]
+ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__nand2_1
XFILLER_147_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_228_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20405_ _07332_ _07341_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24173_ systolic_inst.A_shift\[26\]\[4\] net70 _10505_ systolic_inst.A_shift\[27\]\[4\]
+ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__a22o_1
XFILLER_108_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21385_ _08230_ _08229_ systolic_inst.acc_wires\[4\]\[19\] _11258_ VGND VGND VPWR
+ VPWR _01701_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23124_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[1\]\[9\]
+ VGND VGND VPWR VPWR _09788_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_224_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20336_ _07262_ _07273_ _07274_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__nand3_1
XFILLER_123_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28981_ clknet_leaf_59_clk _02779_ VGND VGND VPWR VPWR systolic_inst.A_shift\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27932_ clknet_leaf_180_clk _01730_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_23055_ _09729_ _09728_ VGND VGND VPWR VPWR _09730_ sky130_fd_sc_hd__nand2b_1
XFILLER_122_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20267_ net109 _07206_ _07207_ _07208_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__o31ai_1
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22006_ systolic_inst.acc_wires\[3\]\[16\] systolic_inst.acc_wires\[3\]\[17\] systolic_inst.acc_wires\[3\]\[18\]
+ systolic_inst.acc_wires\[3\]\[19\] systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__o41a_1
XFILLER_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20198_ _07156_ _07160_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__nor2_1
X_27863_ clknet_leaf_142_clk _01661_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_89_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29602_ clknet_leaf_20_B_in_serial_clk _03397_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_236_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26814_ clknet_leaf_68_clk _00616_ net135 VGND VGND VPWR VPWR B_in\[86\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27794_ clknet_leaf_45_clk _01592_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_186_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29533_ clknet_leaf_258_clk _03331_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[505\]
+ sky130_fd_sc_hd__dfrtp_1
X_26745_ clknet_leaf_51_clk _00547_ net144 VGND VGND VPWR VPWR B_in\[17\] sky130_fd_sc_hd__dfrtp_1
X_23957_ systolic_inst.B_shift\[11\]\[4\] _11332_ net83 systolic_inst.B_shift\[15\]\[4\]
+ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__a22o_1
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13710_ B_in\[17\] deser_B.word_buffer\[17\] net86 VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__mux2_1
X_22908_ _09515_ _09585_ VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__and2_1
XFILLER_56_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26676_ clknet_leaf_10_B_in_serial_clk _00479_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_14690_ systolic_inst.acc_wires\[15\]\[20\] systolic_inst.acc_wires\[15\]\[21\] systolic_inst.acc_wires\[15\]\[22\]
+ systolic_inst.acc_wires\[15\]\[23\] systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _11844_ sky130_fd_sc_hd__o41a_1
X_29464_ clknet_leaf_331_clk _03262_ net136 VGND VGND VPWR VPWR C_out\[436\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23888_ _10473_ _10474_ VGND VGND VPWR VPWR _10475_ sky130_fd_sc_hd__nand2_1
X_13641_ deser_B.word_buffer\[77\] deser_B.serial_word\[77\] net123 VGND VGND VPWR
+ VPWR _00478_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28415_ clknet_leaf_67_clk _02213_ VGND VGND VPWR VPWR systolic_inst.B_shift\[23\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25627_ systolic_inst.acc_wires\[3\]\[7\] C_out\[103\] net48 VGND VGND VPWR VPWR
+ _02929_ sky130_fd_sc_hd__mux2_1
X_22839_ _09513_ _09519_ VGND VGND VPWR VPWR _09520_ sky130_fd_sc_hd__xnor2_1
XFILLER_232_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29395_ clknet_leaf_237_clk _03193_ net145 VGND VGND VPWR VPWR C_out\[367\] sky130_fd_sc_hd__dfrtp_1
XFILLER_201_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16360_ _03658_ _03717_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__xnor2_1
X_25558_ systolic_inst.acc_wires\[1\]\[2\] C_out\[34\] net36 VGND VGND VPWR VPWR _02860_
+ sky130_fd_sc_hd__mux2_1
X_13572_ deser_B.word_buffer\[8\] deser_B.serial_word\[8\] net124 VGND VGND VPWR VPWR
+ _00409_ sky130_fd_sc_hd__mux2_1
X_28346_ clknet_leaf_343_clk _02144_ VGND VGND VPWR VPWR systolic_inst.A_shift\[25\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15311_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[24\]
+ VGND VGND VPWR VPWR _12401_ sky130_fd_sc_hd__and2_1
X_24509_ C_out\[81\] _11302_ net81 ser_C.shift_reg\[81\] _10724_ VGND VGND VPWR VPWR
+ _02331_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_213_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28277_ clknet_leaf_127_clk _02075_ VGND VGND VPWR VPWR systolic_inst.B_shift\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16291_ _03639_ _03641_ _03670_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nand3_1
XFILLER_73_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25489_ _00008_ _11223_ VGND VGND VPWR VPWR _11224_ sky130_fd_sc_hd__nor2_1
XFILLER_199_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15242_ _12340_ _12341_ VGND VGND VPWR VPWR _12342_ sky130_fd_sc_hd__and2_1
X_18030_ _05150_ _05219_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__and2_1
XFILLER_157_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27228_ clknet_leaf_276_clk _01026_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15173_ _12281_ _12282_ _12274_ _12278_ VGND VGND VPWR VPWR _12283_ sky130_fd_sc_hd__a211o_1
X_27159_ clknet_leaf_294_clk _00957_ net138 VGND VGND VPWR VPWR systolic_inst.B_outs\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_201_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14124_ systolic_inst.A_outs\[15\]\[0\] systolic_inst.A_outs\[14\]\[0\] net118 VGND
+ VGND VPWR VPWR _00946_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19981_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[13\] _06976_ net119
+ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__mux2_1
XFILLER_141_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14055_ deser_B.shift_reg\[89\] deser_B.shift_reg\[90\] deser_B.receiving VGND VGND
+ VPWR VPWR _00881_ sky130_fd_sc_hd__mux2_1
X_18932_ _06026_ _06030_ _06032_ net61 VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__a31o_1
XFILLER_140_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_951 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18863_ _05972_ _05973_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__nand2_1
XFILLER_95_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17814_ _05011_ _05012_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nand2_1
XFILLER_239_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18794_ _05914_ _05915_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_199_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17745_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[25\]
+ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__xor2_2
XFILLER_212_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14957_ _12076_ _12077_ VGND VGND VPWR VPWR _12078_ sky130_fd_sc_hd__nor2_1
XFILLER_236_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13908_ deser_A.serial_word\[69\] deser_A.shift_reg\[69\] net57 VGND VGND VPWR VPWR
+ _00734_ sky130_fd_sc_hd__mux2_1
XFILLER_235_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17676_ _04906_ _04909_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_158_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14888_ _11976_ _12010_ VGND VGND VPWR VPWR _12011_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_158_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19415_ _06468_ _06469_ _06461_ _06464_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__a211o_1
X_16627_ _03933_ _03949_ _03951_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__and3_1
XFILLER_223_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13839_ deser_A.serial_word\[0\] deser_A.shift_reg\[0\] net58 VGND VGND VPWR VPWR
+ _00665_ sky130_fd_sc_hd__mux2_1
XFILLER_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19346_ _06404_ _06405_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_154_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16558_ _03902_ _03904_ _03905_ net61 VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__a31o_1
XFILLER_91_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15509_ _12538_ _12566_ VGND VGND VPWR VPWR _12568_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_61_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19277_ net105 _06339_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__or2_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16489_ _03843_ _03845_ _03847_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_14_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18228_ net66 _05405_ _05407_ systolic_inst.acc_wires\[9\]\[5\] net107 VGND VGND
+ VPWR VPWR _01367_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_9_A_in_serial_clk clknet_2_2__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_9_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_113_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18159_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[14\] VGND
+ VGND VPWR VPWR _05346_ sky130_fd_sc_hd__and2_1
XFILLER_172_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21170_ systolic_inst.B_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[5\] VGND VGND VPWR
+ VPWR _08039_ sky130_fd_sc_hd__or2_1
XFILLER_137_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20121_ _07082_ _07089_ _07095_ _07088_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__a211o_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20052_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[6\]\[6\]
+ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__or2_1
XFILLER_86_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24860_ net110 ser_C.shift_reg\[258\] VGND VGND VPWR VPWR _10900_ sky130_fd_sc_hd__and2_1
XFILLER_86_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23811_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[18\]
+ VGND VGND VPWR VPWR _10410_ sky130_fd_sc_hd__or2_1
XFILLER_2_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24791_ C_out\[222\] net99 net79 ser_C.shift_reg\[222\] _10865_ VGND VGND VPWR VPWR
+ _02472_ sky130_fd_sc_hd__a221o_1
XFILLER_6_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26530_ clknet_leaf_5_A_in_serial_clk _00333_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_214_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23742_ _10347_ _10348_ _10346_ VGND VGND VPWR VPWR _10351_ sky130_fd_sc_hd__a21bo_1
XFILLER_148_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ _07826_ _07827_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_217_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_217_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26461_ clknet_leaf_1_A_in_serial_clk _00268_ net132 VGND VGND VPWR VPWR deser_A.bit_idx\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_23673_ _10266_ _10272_ _10291_ VGND VGND VPWR VPWR _10292_ sky130_fd_sc_hd__o21ai_1
X_20885_ _07742_ _07760_ _07761_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__or3_1
X_28200_ clknet_leaf_129_clk _01998_ VGND VGND VPWR VPWR systolic_inst.B_shift\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_25412_ _11175_ systolic_inst.A_shift\[1\]\[5\] net71 VGND VGND VPWR VPWR _02783_
+ sky130_fd_sc_hd__mux2_1
X_22624_ _09296_ _09297_ _09317_ _09336_ VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__a211o_1
X_29180_ clknet_leaf_135_clk _02978_ net142 VGND VGND VPWR VPWR C_out\[152\] sky130_fd_sc_hd__dfrtp_1
X_26392_ clknet_leaf_16_clk _00199_ net132 VGND VGND VPWR VPWR A_in\[60\] sky130_fd_sc_hd__dfrtp_1
X_28131_ clknet_leaf_129_clk _01929_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_23_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25343_ ser_C.parallel_data\[498\] net102 net77 ser_C.shift_reg\[498\] _11141_ VGND
+ VGND VPWR VPWR _02748_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_12_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22555_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[2\]\[12\]
+ _09276_ _09278_ VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__a211o_1
XFILLER_139_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28062_ clknet_leaf_121_clk _01860_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_21506_ _08312_ _08318_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25274_ net111 ser_C.shift_reg\[465\] VGND VGND VPWR VPWR _11107_ sky130_fd_sc_hd__and2_1
X_22486_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[2\]\[3\]
+ VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__or2_1
XFILLER_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27013_ clknet_leaf_21_B_in_serial_clk _00811_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24225_ systolic_inst.A_shift\[20\]\[4\] A_in\[76\] net59 VGND VGND VPWR VPWR _10598_
+ sky130_fd_sc_hd__mux2_1
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21437_ _08273_ _08274_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24156_ _10579_ systolic_inst.A_shift\[27\]\[1\] net70 VGND VGND VPWR VPWR _02123_
+ sky130_fd_sc_hd__mux2_1
XFILLER_162_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21368_ _11713_ _08216_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__nor2_1
XFILLER_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23107_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[1\]\[6\]
+ VGND VGND VPWR VPWR _09774_ sky130_fd_sc_hd__or2_1
X_20319_ _07256_ _07257_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__or2_1
X_28964_ clknet_leaf_79_clk _02762_ VGND VGND VPWR VPWR systolic_inst.B_shift\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24087_ systolic_inst.B_shift\[2\]\[6\] _11332_ net83 systolic_inst.B_shift\[6\]\[6\]
+ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_57_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21299_ _08149_ _08153_ _08155_ _08156_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__o211ai_2
XFILLER_107_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23038_ net109 systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[14\] VGND
+ VGND VPWR VPWR _09713_ sky130_fd_sc_hd__and2_1
XFILLER_153_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27915_ clknet_leaf_135_clk _01713_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28895_ clknet_leaf_285_clk _02693_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[443\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27846_ clknet_leaf_179_clk _01644_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_15860_ _12892_ _12893_ VGND VGND VPWR VPWR _12894_ sky130_fd_sc_hd__and2_1
XFILLER_77_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_202_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_202_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14811_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[4\]
+ systolic_inst.A_outs\[14\]\[5\] VGND VGND VPWR VPWR _11936_ sky130_fd_sc_hd__and4_1
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27777_ clknet_leaf_176_clk _01575_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15791_ _12832_ _12833_ _12834_ VGND VGND VPWR VPWR _12835_ sky130_fd_sc_hd__a21o_1
XFILLER_79_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24989_ C_out\[321\] net102 net74 ser_C.shift_reg\[321\] _10964_ VGND VGND VPWR VPWR
+ _02571_ sky130_fd_sc_hd__a221o_1
XFILLER_229_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29516_ clknet_leaf_255_clk _03314_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[488\]
+ sky130_fd_sc_hd__dfrtp_1
X_17530_ _04714_ _04751_ _04750_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_194_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26728_ clknet_leaf_73_clk _00530_ net144 VGND VGND VPWR VPWR B_in\[0\] sky130_fd_sc_hd__dfrtp_1
X_14742_ systolic_inst.A_outs\[14\]\[2\] systolic_inst.A_outs\[13\]\[2\] net120 VGND
+ VGND VPWR VPWR _01012_ sky130_fd_sc_hd__mux2_1
XFILLER_233_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_194_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14673_ _11820_ _11826_ _11827_ net61 VGND VGND VPWR VPWR _11830_ sky130_fd_sc_hd__a31o_1
X_29447_ clknet_leaf_300_clk _03245_ net139 VGND VGND VPWR VPWR C_out\[419\] sky130_fd_sc_hd__dfrtp_1
X_17461_ systolic_inst.B_outs\[10\]\[5\] systolic_inst.A_outs\[10\]\[6\] VGND VGND
+ VPWR VPWR _04715_ sky130_fd_sc_hd__nand2_1
XFILLER_233_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26659_ clknet_leaf_2_B_in_serial_clk _00462_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[61\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_192_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_192_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19200_ _06264_ _06234_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__nand2b_1
XFILLER_44_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13624_ deser_B.word_buffer\[60\] deser_B.serial_word\[60\] net123 VGND VGND VPWR
+ VPWR _00461_ sky130_fd_sc_hd__mux2_1
X_16412_ _03780_ _03781_ _03775_ _03778_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__a211o_1
XFILLER_60_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29378_ clknet_leaf_244_clk _03176_ net145 VGND VGND VPWR VPWR C_out\[350\] sky130_fd_sc_hd__dfrtp_1
X_17392_ systolic_inst.A_outs\[10\]\[4\] systolic_inst.B_outs\[10\]\[5\] VGND VGND
+ VPWR VPWR _04648_ sky130_fd_sc_hd__nand2_1
XFILLER_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19131_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[6\] _06197_ net119
+ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16343_ _03720_ _03721_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__nor2_1
XFILLER_41_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28329_ clknet_leaf_2_clk _02127_ VGND VGND VPWR VPWR systolic_inst.A_shift\[27\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13555_ deser_A.shift_reg\[119\] deser_A.shift_reg\[120\] net130 VGND VGND VPWR VPWR
+ _00392_ sky130_fd_sc_hd__mux2_1
XFILLER_201_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19062_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[3\]
+ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__and3_1
X_16274_ _03654_ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__xnor2_1
X_13486_ deser_A.shift_reg\[50\] deser_A.shift_reg\[51\] net130 VGND VGND VPWR VPWR
+ _00323_ sky130_fd_sc_hd__mux2_1
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15225_ _12298_ _12301_ _12310_ _12326_ VGND VGND VPWR VPWR _12327_ sky130_fd_sc_hd__a211o_1
X_18013_ _05166_ _05168_ _05204_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__a21o_1
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15156_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[14\]\[2\]
+ VGND VGND VPWR VPWR _12268_ sky130_fd_sc_hd__and2_1
XFILLER_236_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14107_ systolic_inst.A_shift\[12\]\[7\] net71 _11333_ A_in\[63\] VGND VGND VPWR
+ VPWR _00929_ sky130_fd_sc_hd__a22o_1
XFILLER_236_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19964_ _06895_ _06959_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__nand2_1
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15087_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[12\] _12204_ net118
+ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__mux2_1
XFILLER_234_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14038_ deser_B.shift_reg\[72\] deser_B.shift_reg\[73\] deser_B.receiving VGND VGND
+ VPWR VPWR _00864_ sky130_fd_sc_hd__mux2_1
X_18915_ _06014_ _06017_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__or2_1
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19895_ systolic_inst.B_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\] VGND VGND VPWR
+ VPWR _06893_ sky130_fd_sc_hd__or2_1
XFILLER_136_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18846_ _05952_ _05954_ _05958_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__a21o_1
XFILLER_228_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18777_ _05871_ _05873_ _05898_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__and3_1
X_15989_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _12989_ sky130_fd_sc_hd__and2_1
XFILLER_36_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17728_ _04951_ _04952_ _04953_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_102_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_B_in_serial_clk clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_16_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_36_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17659_ _04892_ _04893_ _04894_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_183_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_183_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20670_ _07587_ _07588_ _07586_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__a21bo_1
XFILLER_211_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19329_ _06345_ _06361_ _06359_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__o21a_1
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22340_ _09081_ _09082_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__nand2_1
XFILLER_31_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22271_ _08978_ _08979_ _08977_ VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24010_ systolic_inst.B_shift\[7\]\[1\] net70 net83 systolic_inst.B_shift\[11\]\[1\]
+ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__a22o_1
XFILLER_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21222_ _11271_ systolic_inst.A_outs\[4\]\[7\] _07850_ _08062_ VGND VGND VPWR VPWR
+ _08089_ sky130_fd_sc_hd__o211a_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21153_ _08021_ _08022_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__nor2_1
XFILLER_219_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20104_ net60 _07083_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__nor2_1
XFILLER_160_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21084_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\] systolic_inst.A_outs\[4\]\[6\]
+ systolic_inst.A_outs\[4\]\[7\] VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__and4_1
XFILLER_115_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25961_ systolic_inst.acc_wires\[13\]\[21\] C_out\[437\] net20 VGND VGND VPWR VPWR
+ _03263_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27700_ clknet_leaf_198_clk _01498_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_20035_ _07024_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24912_ net110 ser_C.shift_reg\[284\] VGND VGND VPWR VPWR _10926_ sky130_fd_sc_hd__and2_1
X_28680_ clknet_leaf_195_clk _02478_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25892_ systolic_inst.acc_wires\[11\]\[16\] C_out\[368\] net40 VGND VGND VPWR VPWR
+ _03194_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_219_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27631_ clknet_leaf_324_clk _01429_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24843_ C_out\[248\] net98 net78 ser_C.shift_reg\[248\] _10891_ VGND VGND VPWR VPWR
+ _02498_ sky130_fd_sc_hd__a221o_1
XFILLER_27_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24774_ net113 ser_C.shift_reg\[215\] VGND VGND VPWR VPWR _10857_ sky130_fd_sc_hd__and2_1
X_27562_ clknet_leaf_306_clk _01360_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_21986_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[16\]
+ _08766_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__a21oi_1
X_29301_ clknet_leaf_312_clk _03099_ net141 VGND VGND VPWR VPWR C_out\[273\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23725_ _10334_ _10335_ _10336_ VGND VGND VPWR VPWR _10337_ sky130_fd_sc_hd__a21o_1
XFILLER_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26513_ clknet_leaf_11_A_in_serial_clk _00316_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_20937_ systolic_inst.B_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[5\] systolic_inst.B_outs\[4\]\[5\]
+ systolic_inst.A_outs\[4\]\[1\] VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_174_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_174_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27493_ clknet_leaf_227_clk _01291_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_226_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29232_ clknet_leaf_204_clk _03030_ net147 VGND VGND VPWR VPWR C_out\[204\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23656_ _10224_ _10227_ _10274_ _10275_ VGND VGND VPWR VPWR _10276_ sky130_fd_sc_hd__a211oi_2
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26444_ clknet_leaf_347_clk _00251_ net132 VGND VGND VPWR VPWR A_in\[112\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20868_ _07744_ _07745_ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__nand2b_1
XFILLER_186_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22607_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[20\]
+ _09321_ VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_46_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26375_ clknet_leaf_28_clk _00182_ net133 VGND VGND VPWR VPWR A_in\[43\] sky130_fd_sc_hd__dfrtp_1
X_29163_ clknet_leaf_40_clk _02961_ net142 VGND VGND VPWR VPWR C_out\[135\] sky130_fd_sc_hd__dfrtp_1
XFILLER_161_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23587_ _10191_ _10207_ VGND VGND VPWR VPWR _10209_ sky130_fd_sc_hd__and2_1
XFILLER_139_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20799_ _07694_ _07698_ _07695_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__a21bo_1
XFILLER_70_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28114_ clknet_leaf_47_clk _01912_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_10_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25326_ net112 ser_C.shift_reg\[491\] VGND VGND VPWR VPWR _11133_ sky130_fd_sc_hd__and2_1
X_13340_ A_in\[49\] deser_A.word_buffer\[49\] net92 VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__mux2_1
X_22538_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[2\]\[11\]
+ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__nor2_1
XFILLER_210_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29094_ clknet_leaf_112_clk _02892_ net150 VGND VGND VPWR VPWR C_out\[66\] sky130_fd_sc_hd__dfrtp_1
XFILLER_154_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28045_ clknet_leaf_128_clk _01843_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_25257_ ser_C.parallel_data\[455\] net102 net74 ser_C.shift_reg\[455\] _11098_ VGND
+ VGND VPWR VPWR _02705_ sky130_fd_sc_hd__a221o_1
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13271_ deser_A.word_buffer\[109\] deser_A.serial_word\[109\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__mux2_1
X_22469_ net122 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[2\]\[0\]
+ VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__a21oi_1
XFILLER_202_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15010_ _12072_ _12129_ VGND VGND VPWR VPWR _12130_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_187_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24208_ _10589_ systolic_inst.A_shift\[20\]\[3\] net71 VGND VGND VPWR VPWR _02165_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25188_ net111 ser_C.shift_reg\[422\] VGND VGND VPWR VPWR _11064_ sky130_fd_sc_hd__and2_1
XFILLER_237_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24139_ systolic_inst.A_shift\[29\]\[1\] A_in\[105\] net59 VGND VGND VPWR VPWR _10571_
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_183_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_63_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_204_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_204_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28947_ clknet_leaf_258_clk _02745_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[495\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16961_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[14\] _04275_ net119
+ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__mux2_1
XFILLER_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18700_ _05825_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__inv_2
XFILLER_237_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15912_ _12917_ _12937_ VGND VGND VPWR VPWR _12938_ sky130_fd_sc_hd__nor2_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19680_ _06651_ _06671_ _06673_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_196_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28878_ clknet_leaf_289_clk _02676_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[426\]
+ sky130_fd_sc_hd__dfrtp_1
X_16892_ _04169_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18631_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__inv_2
X_27829_ clknet_leaf_141_clk _01627_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15843_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[13\]\[14\]
+ VGND VGND VPWR VPWR _12879_ sky130_fd_sc_hd__or2_1
XFILLER_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18562_ _05628_ _05663_ _05662_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__a21bo_1
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15774_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[13\]\[4\]
+ VGND VGND VPWR VPWR _12820_ sky130_fd_sc_hd__nand2_1
XFILLER_64_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1096 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17513_ _04765_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__inv_2
X_14725_ _11866_ _11869_ _11868_ VGND VGND VPWR VPWR _11874_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_165_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_165_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18493_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[5\] _05623_
+ _05624_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17444_ _04697_ _04698_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__nand2_1
X_14656_ net107 systolic_inst.acc_wires\[15\]\[18\] net69 _11815_ VGND VGND VPWR VPWR
+ _00996_ sky130_fd_sc_hd__a22o_1
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13607_ deser_B.word_buffer\[43\] deser_B.serial_word\[43\] net124 VGND VGND VPWR
+ VPWR _00444_ sky130_fd_sc_hd__mux2_1
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17375_ _04630_ _04631_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__nor2_1
XFILLER_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14587_ _11751_ _11754_ VGND VGND VPWR VPWR _11756_ sky130_fd_sc_hd__nand2_1
XFILLER_229_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19114_ systolic_inst.A_outs\[7\]\[1\] systolic_inst.B_outs\[7\]\[6\] VGND VGND VPWR
+ VPWR _06181_ sky130_fd_sc_hd__nand2_1
XFILLER_159_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16326_ _03703_ _03704_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__and2b_1
XFILLER_185_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13538_ deser_A.shift_reg\[102\] deser_A.shift_reg\[103\] net129 VGND VGND VPWR VPWR
+ _00375_ sky130_fd_sc_hd__mux2_1
XFILLER_199_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19045_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[2\]
+ systolic_inst.A_outs\[7\]\[3\] VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__nand4_2
X_16257_ _03638_ _03637_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__nand2b_1
X_13469_ deser_A.shift_reg\[33\] deser_A.shift_reg\[34\] deser_A.receiving VGND VGND
+ VPWR VPWR _00306_ sky130_fd_sc_hd__mux2_1
XFILLER_199_1085 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15208_ net61 _12312_ VGND VGND VPWR VPWR _12313_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16188_ _03569_ _03570_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15139_ _12030_ _12173_ _12245_ _12243_ VGND VGND VPWR VPWR _12254_ sky130_fd_sc_hd__a31o_1
XFILLER_153_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19947_ _06942_ _06943_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__or2_1
XFILLER_87_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19878_ _06876_ _06875_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_3_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18829_ net63 _05943_ _05945_ systolic_inst.acc_wires\[8\]\[4\] net108 VGND VGND
+ VPWR VPWR _01430_ sky130_fd_sc_hd__a32o_1
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21840_ _08556_ _08642_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_90_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21771_ _08538_ _08540_ _08574_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_156_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_156_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_224_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23510_ _10089_ _10092_ _10132_ _10133_ VGND VGND VPWR VPWR _10134_ sky130_fd_sc_hd__a211o_2
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20722_ _07628_ _07632_ _07634_ _07635_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__a211o_1
X_24490_ net112 ser_C.shift_reg\[73\] VGND VGND VPWR VPWR _10715_ sky130_fd_sc_hd__and2_1
XFILLER_145_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23441_ systolic_inst.A_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[5\] _10025_ VGND
+ VGND VPWR VPWR _10066_ sky130_fd_sc_hd__and3_1
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20653_ _07574_ _07575_ _07576_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__a21o_1
XFILLER_51_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26160_ deser_B.serial_word\[115\] deser_B.shift_reg\[115\] net56 VGND VGND VPWR
+ VPWR _03462_ sky130_fd_sc_hd__mux2_1
XFILLER_137_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23372_ systolic_inst.A_outs\[0\]\[2\] systolic_inst.B_outs\[0\]\[3\] systolic_inst.A_outs\[0\]\[3\]
+ systolic_inst.B_outs\[0\]\[4\] VGND VGND VPWR VPWR _09999_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_134_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20584_ _07514_ _07515_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_134_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25111_ C_out\[382\] net97 net77 ser_C.shift_reg\[382\] _11025_ VGND VGND VPWR VPWR
+ _02632_ sky130_fd_sc_hd__a221o_1
X_22323_ _09064_ _09065_ VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26091_ deser_B.serial_word\[46\] deser_B.shift_reg\[46\] net55 VGND VGND VPWR VPWR
+ _03393_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25042_ net113 ser_C.shift_reg\[349\] VGND VGND VPWR VPWR _10991_ sky130_fd_sc_hd__and2_1
XFILLER_219_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22254_ _08995_ _08998_ VGND VGND VPWR VPWR _08999_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21205_ _07991_ _08072_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__nand2_1
XFILLER_219_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22185_ _08925_ _08926_ _08930_ VGND VGND VPWR VPWR _08932_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_240_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_240_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28801_ clknet_leaf_240_clk _02599_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[349\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_160_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21136_ _08004_ _08005_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__nor2_1
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26993_ clknet_leaf_0_A_in_serial_clk _00791_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28732_ clknet_leaf_302_clk _02530_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[280\]
+ sky130_fd_sc_hd__dfrtp_1
X_21067_ _07922_ _07938_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__nor2_1
X_25944_ systolic_inst.acc_wires\[13\]\[4\] C_out\[420\] net27 VGND VGND VPWR VPWR
+ _03246_ sky130_fd_sc_hd__mux2_1
XFILLER_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20018_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[6\]\[1\]
+ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__or2_1
XFILLER_86_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28663_ clknet_leaf_176_clk _02461_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[211\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_Left_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25875_ systolic_inst.acc_wires\[10\]\[31\] C_out\[351\] net41 VGND VGND VPWR VPWR
+ _03177_ sky130_fd_sc_hd__mux2_1
XFILLER_104_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27614_ clknet_leaf_321_clk _01412_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_238_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24826_ net113 ser_C.shift_reg\[241\] VGND VGND VPWR VPWR _10883_ sky130_fd_sc_hd__and2_1
XFILLER_62_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28594_ clknet_leaf_43_clk _02392_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[142\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_238_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27545_ clknet_leaf_34_clk _01343_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_21969_ _08748_ _08751_ _08754_ VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__a21oi_1
X_24757_ C_out\[205\] net99 net79 ser_C.shift_reg\[205\] _10848_ VGND VGND VPWR VPWR
+ _02455_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_147_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_147_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_48_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14510_ _11620_ _11689_ VGND VGND VPWR VPWR _11690_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23708_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[0\]\[3\]
+ VGND VGND VPWR VPWR _10322_ sky130_fd_sc_hd__nand2_1
X_15490_ systolic_inst.A_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[4\]
+ systolic_inst.B_outs\[13\]\[3\] VGND VGND VPWR VPWR _12549_ sky130_fd_sc_hd__a22oi_1
XFILLER_214_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24688_ net112 ser_C.shift_reg\[172\] VGND VGND VPWR VPWR _10814_ sky130_fd_sc_hd__and2_1
X_27476_ clknet_leaf_306_clk _01274_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29215_ clknet_leaf_180_clk _03013_ net148 VGND VGND VPWR VPWR C_out\[187\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23639_ _10257_ _10258_ VGND VGND VPWR VPWR _10259_ sky130_fd_sc_hd__nor2_1
XFILLER_120_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14441_ systolic_inst.B_outs\[15\]\[6\] systolic_inst.A_outs\[15\]\[6\] _11273_ systolic_inst.A_outs\[15\]\[5\]
+ VGND VGND VPWR VPWR _11623_ sky130_fd_sc_hd__o2bb2a_1
X_26427_ clknet_leaf_4_clk _00234_ net133 VGND VGND VPWR VPWR A_in\[95\] sky130_fd_sc_hd__dfrtp_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29146_ clknet_leaf_175_clk _02944_ net150 VGND VGND VPWR VPWR C_out\[118\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17160_ net105 systolic_inst.acc_wires\[11\]\[28\] net62 _04444_ VGND VGND VPWR VPWR
+ _01262_ sky130_fd_sc_hd__a22o_1
X_14372_ _11554_ _11555_ VGND VGND VPWR VPWR _11556_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_189_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26358_ clknet_leaf_65_clk _00165_ net134 VGND VGND VPWR VPWR A_in\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1056 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13323_ A_in\[32\] deser_A.word_buffer\[32\] net93 VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__mux2_1
X_16111_ _13099_ _03496_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__nor2_1
XFILLER_127_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25309_ ser_C.parallel_data\[481\] net102 net74 ser_C.shift_reg\[481\] _11124_ VGND
+ VGND VPWR VPWR _02731_ sky130_fd_sc_hd__a221o_1
XFILLER_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29077_ clknet_leaf_155_clk _02875_ net150 VGND VGND VPWR VPWR C_out\[49\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26289_ clknet_leaf_26_A_in_serial_clk _00097_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_17091_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[18\]
+ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_185_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28028_ clknet_leaf_162_clk _01826_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_196_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16042_ _13037_ _13038_ VGND VGND VPWR VPWR _13039_ sky130_fd_sc_hd__and2b_1
X_13254_ deser_A.word_buffer\[92\] deser_A.serial_word\[92\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__mux2_1
XFILLER_170_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13185_ deser_A.word_buffer\[23\] deser_A.serial_word\[23\] net128 VGND VGND VPWR
+ VPWR _00033_ sky130_fd_sc_hd__mux2_1
X_19801_ _06792_ _06800_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_144_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17993_ net116 _05183_ _05184_ _05185_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__a31o_1
XFILLER_46_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19732_ _06689_ _06691_ _06733_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__and3_1
X_16944_ _04257_ _04258_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__nand2_1
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19663_ _06667_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__inv_2
XFILLER_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16875_ _04155_ _04161_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__or3_1
XFILLER_238_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18614_ systolic_inst.A_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[6\] _11259_ systolic_inst.A_outs\[8\]\[2\]
+ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__o2bb2a_1
X_15826_ net108 systolic_inst.acc_wires\[13\]\[11\] net67 _12864_ VGND VGND VPWR VPWR
+ _01117_ sky130_fd_sc_hd__a22o_1
X_19594_ net106 systolic_inst.acc_wires\[7\]\[28\] net62 _06622_ VGND VGND VPWR VPWR
+ _01518_ sky130_fd_sc_hd__a22o_1
XFILLER_37_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18545_ _05639_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_138_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15757_ _12805_ VGND VGND VPWR VPWR _12806_ sky130_fd_sc_hd__inv_2
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14708_ _11857_ _11859_ VGND VGND VPWR VPWR _11860_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18476_ systolic_inst.A_outs\[8\]\[2\] systolic_inst.B_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\]
+ systolic_inst.A_outs\[8\]\[1\] VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_174_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ _12672_ _12678_ _12708_ _12707_ VGND VGND VPWR VPWR _12742_ sky130_fd_sc_hd__a31o_1
XFILLER_33_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17427_ _04680_ _04681_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_99_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14639_ _11799_ _11800_ VGND VGND VPWR VPWR _11801_ sky130_fd_sc_hd__and2_1
XFILLER_53_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17358_ _04613_ _04614_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__nor2_1
XFILLER_179_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16309_ systolic_inst.B_outs\[12\]\[6\] systolic_inst.A_outs\[12\]\[7\] VGND VGND
+ VPWR VPWR _03689_ sky130_fd_sc_hd__nand2_1
Xclkload300 clknet_leaf_180_clk VGND VGND VPWR VPWR clkload300/Y sky130_fd_sc_hd__inv_8
XFILLER_147_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload311 clknet_leaf_151_clk VGND VGND VPWR VPWR clkload311/Y sky130_fd_sc_hd__inv_8
XFILLER_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17289_ _04519_ _04546_ _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_310_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_310_clk
+ sky130_fd_sc_hd__clkbuf_8
Xclkload322 clknet_leaf_157_clk VGND VGND VPWR VPWR clkload322/Y sky130_fd_sc_hd__clkinv_4
XFILLER_88_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload333 clknet_leaf_161_clk VGND VGND VPWR VPWR clkload333/X sky130_fd_sc_hd__clkbuf_8
Xclkload30 clknet_leaf_335_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__clkinv_2
X_19028_ net105 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[0\] _06100_
+ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__a21o_1
Xclkload41 clknet_leaf_341_clk VGND VGND VPWR VPWR clkload41/Y sky130_fd_sc_hd__inv_6
Xclkload344 clknet_leaf_29_A_in_serial_clk VGND VGND VPWR VPWR clkload344/Y sky130_fd_sc_hd__inv_8
XFILLER_146_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload52 clknet_leaf_302_clk VGND VGND VPWR VPWR clkload52/Y sky130_fd_sc_hd__inv_6
Xclkload355 clknet_leaf_6_A_in_serial_clk VGND VGND VPWR VPWR clkload355/Y sky130_fd_sc_hd__bufinv_16
Xclkload366 clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR clkload366/Y sky130_fd_sc_hd__inv_6
XFILLER_155_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload63 clknet_leaf_4_clk VGND VGND VPWR VPWR clkload63/Y sky130_fd_sc_hd__clkinv_4
XFILLER_86_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload377 clknet_leaf_32_B_in_serial_clk VGND VGND VPWR VPWR clkload377/X sky130_fd_sc_hd__clkbuf_8
Xclkload74 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload74/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload388 clknet_leaf_8_B_in_serial_clk VGND VGND VPWR VPWR clkload388/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_90_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload85 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload85/Y sky130_fd_sc_hd__clkinv_2
Xclkload96 clknet_leaf_217_clk VGND VGND VPWR VPWR clkload96/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_90_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23990_ _10520_ systolic_inst.B_shift\[8\]\[6\] net72 VGND VGND VPWR VPWR _02016_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22941_ net122 _09619_ VGND VGND VPWR VPWR _09620_ sky130_fd_sc_hd__nand2_1
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22872_ _09513_ _09519_ _09518_ VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__a21o_1
X_25660_ systolic_inst.acc_wires\[4\]\[8\] C_out\[136\] net29 VGND VGND VPWR VPWR
+ _02962_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21823_ _08625_ _08626_ VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_30_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24611_ C_out\[132\] net103 net75 ser_C.shift_reg\[132\] _10775_ VGND VGND VPWR VPWR
+ _02382_ sky130_fd_sc_hd__a221o_1
X_25591_ systolic_inst.acc_wires\[2\]\[3\] C_out\[67\] net34 VGND VGND VPWR VPWR _02893_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_129_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_233_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24542_ net113 ser_C.shift_reg\[99\] VGND VGND VPWR VPWR _10741_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27330_ clknet_leaf_287_clk _01128_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_21754_ _08558_ _08559_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__nor2_1
XFILLER_52_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_233_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20705_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[5\]\[13\]
+ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__xor2_1
X_24473_ C_out\[63\] net100 net82 ser_C.shift_reg\[63\] _10706_ VGND VGND VPWR VPWR
+ _02313_ sky130_fd_sc_hd__a221o_1
XFILLER_180_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27261_ clknet_leaf_271_clk _01059_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_43_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21685_ _08491_ _08492_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_43_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29000_ clknet_leaf_92_clk _02798_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23424_ _10048_ _10049_ VGND VGND VPWR VPWR _10050_ sky130_fd_sc_hd__nand2b_1
XFILLER_138_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26212_ clknet_leaf_13_A_in_serial_clk _00020_ net144 VGND VGND VPWR VPWR deser_A.word_buffer\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_184_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20636_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[5\]\[3\]
+ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__nand2_1
X_27192_ clknet_leaf_255_clk _00990_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload2 clknet_5_2__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_12
XFILLER_177_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26143_ deser_B.serial_word\[98\] deser_B.shift_reg\[98\] _00001_ VGND VGND VPWR
+ VPWR _03445_ sky130_fd_sc_hd__mux2_1
X_23355_ _09955_ _09957_ VGND VGND VPWR VPWR _09983_ sky130_fd_sc_hd__nand2b_1
XFILLER_164_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20567_ _07467_ _07470_ _07498_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__o21ai_1
XFILLER_137_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_A_in_serial_clk clknet_2_1__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_22_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_301_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_301_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_221_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22306_ _09049_ VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__inv_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26074_ deser_B.serial_word\[29\] deser_B.shift_reg\[29\] net56 VGND VGND VPWR VPWR
+ _03376_ sky130_fd_sc_hd__mux2_1
XFILLER_192_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23286_ _11258_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[0\] _09918_
+ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__a21o_1
X_20498_ _07430_ _07431_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__or2_1
XFILLER_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25025_ C_out\[339\] net97 net77 ser_C.shift_reg\[339\] _10982_ VGND VGND VPWR VPWR
+ _02589_ sky130_fd_sc_hd__a221o_1
XFILLER_30_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22237_ systolic_inst.B_outs\[2\]\[7\] _08948_ _08949_ VGND VGND VPWR VPWR _08982_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_180_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22168_ systolic_inst.A_outs\[2\]\[4\] _08878_ _08896_ _08895_ _08892_ VGND VGND
+ VPWR VPWR _08915_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_37_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21119_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[7\] _07960_ _07884_
+ systolic_inst.A_outs\[4\]\[5\] VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__a32o_1
XFILLER_232_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22099_ _08850_ _08848_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[1\]
+ net109 VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_182_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14990_ systolic_inst.A_outs\[14\]\[6\] _12109_ _12108_ VGND VGND VPWR VPWR _12110_
+ sky130_fd_sc_hd__a21bo_1
X_26976_ clknet_leaf_28_A_in_serial_clk _00774_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_28715_ clknet_leaf_314_clk _02513_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[263\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25927_ systolic_inst.acc_wires\[12\]\[19\] C_out\[403\] net17 VGND VGND VPWR VPWR
+ _03229_ sky130_fd_sc_hd__mux2_1
X_13941_ deser_A.serial_word\[102\] deser_A.shift_reg\[102\] net57 VGND VGND VPWR
+ VPWR _00767_ sky130_fd_sc_hd__mux2_1
XFILLER_232_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29695_ clknet_leaf_11_clk _03490_ VGND VGND VPWR VPWR systolic_inst.A_shift\[30\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28646_ clknet_leaf_202_clk _02444_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[194\]
+ sky130_fd_sc_hd__dfrtp_1
X_16660_ _03942_ _03959_ _03958_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_178_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13872_ deser_A.serial_word\[33\] deser_A.shift_reg\[33\] net58 VGND VGND VPWR VPWR
+ _00698_ sky130_fd_sc_hd__mux2_1
X_25858_ systolic_inst.acc_wires\[10\]\[14\] C_out\[334\] net12 VGND VGND VPWR VPWR
+ _03160_ sky130_fd_sc_hd__mux2_1
XFILLER_207_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15611_ _12666_ _12665_ VGND VGND VPWR VPWR _12667_ sky130_fd_sc_hd__nand2b_1
X_24809_ C_out\[231\] net99 net79 ser_C.shift_reg\[231\] _10874_ VGND VGND VPWR VPWR
+ _02481_ sky130_fd_sc_hd__a221o_1
X_28577_ clknet_leaf_172_clk _02375_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[125\]
+ sky130_fd_sc_hd__dfrtp_1
X_16591_ net118 systolic_inst.B_outs\[11\]\[0\] systolic_inst.A_outs\[11\]\[0\] VGND
+ VGND VPWR VPWR _03920_ sky130_fd_sc_hd__and3_1
X_25789_ systolic_inst.acc_wires\[8\]\[9\] C_out\[265\] net22 VGND VGND VPWR VPWR
+ _03091_ sky130_fd_sc_hd__mux2_1
XFILLER_90_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18330_ systolic_inst.acc_wires\[9\]\[16\] systolic_inst.acc_wires\[9\]\[17\] systolic_inst.acc_wires\[9\]\[18\]
+ systolic_inst.acc_wires\[9\]\[19\] systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__o41a_1
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15542_ _12546_ _12561_ _12560_ VGND VGND VPWR VPWR _12600_ sky130_fd_sc_hd__o21a_1
XFILLER_76_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27528_ clknet_leaf_240_clk _01326_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18261_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[9\]\[11\]
+ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__nand2_1
X_27459_ clknet_leaf_237_clk _01257_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_15473_ _12499_ _12501_ _12531_ _12532_ VGND VGND VPWR VPWR _12533_ sky130_fd_sc_hd__a211oi_1
X_17212_ systolic_inst.A_outs\[10\]\[0\] systolic_inst.A_outs\[10\]\[1\] systolic_inst.B_outs\[10\]\[3\]
+ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__and3_1
X_14424_ _11604_ _11605_ VGND VGND VPWR VPWR _11607_ sky130_fd_sc_hd__xor2_1
XFILLER_198_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18192_ net116 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[9\]\[0\]
+ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__a21oi_1
XFILLER_126_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29129_ clknet_leaf_171_clk _02927_ net148 VGND VGND VPWR VPWR C_out\[101\] sky130_fd_sc_hd__dfrtp_1
XFILLER_155_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17143_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[26\]
+ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__nand2_1
X_14355_ _11523_ _11539_ VGND VGND VPWR VPWR _11540_ sky130_fd_sc_hd__xor2_1
XFILLER_156_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13306_ A_in\[15\] deser_A.word_buffer\[15\] net93 VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__mux2_1
XFILLER_156_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14286_ _11434_ _11471_ _11472_ VGND VGND VPWR VPWR _11473_ sky130_fd_sc_hd__o21ba_1
X_17074_ _04362_ _04367_ _04371_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16025_ _13002_ _13019_ _13021_ VGND VGND VPWR VPWR _13023_ sky130_fd_sc_hd__and3_1
X_13237_ deser_A.word_buffer\[75\] deser_A.serial_word\[75\] net127 VGND VGND VPWR
+ VPWR _00085_ sky130_fd_sc_hd__mux2_1
XFILLER_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13168_ deser_A.word_buffer\[6\] deser_A.serial_word\[6\] net127 VGND VGND VPWR VPWR
+ _00016_ sky130_fd_sc_hd__mux2_1
XFILLER_135_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17976_ _05159_ _05167_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__xnor2_1
XFILLER_242_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19715_ _06687_ _06716_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__nor2_1
XFILLER_211_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16927_ _04199_ _04212_ _04210_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__o21a_1
XFILLER_111_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19646_ _06650_ _06651_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__or2_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16858_ _04175_ _04174_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__nand2b_1
XFILLER_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15809_ _12845_ _12847_ VGND VGND VPWR VPWR _12850_ sky130_fd_sc_hd__nand2_1
X_19577_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[26\]
+ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__nand2_1
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16789_ _04106_ _04107_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18528_ systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[6\] systolic_inst.A_outs\[8\]\[7\]
+ systolic_inst.B_outs\[8\]\[0\] VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__a22o_1
XFILLER_222_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18459_ _05572_ _05589_ _05590_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__or3_1
XFILLER_194_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21470_ systolic_inst.A_outs\[3\]\[6\] systolic_inst.A_outs\[2\]\[6\] net122 VGND
+ VGND VPWR VPWR _01720_ sky130_fd_sc_hd__mux2_1
XFILLER_193_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20421_ net109 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[8\] VGND
+ VGND VPWR VPWR _07358_ sky130_fd_sc_hd__and2_1
XFILLER_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23140_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[1\]\[11\]
+ VGND VGND VPWR VPWR _09802_ sky130_fd_sc_hd__nand2_1
XFILLER_134_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20352_ _07288_ _07289_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__and2b_1
Xclkload130 clknet_leaf_265_clk VGND VGND VPWR VPWR clkload130/Y sky130_fd_sc_hd__bufinv_16
XFILLER_88_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload141 clknet_leaf_256_clk VGND VGND VPWR VPWR clkload141/X sky130_fd_sc_hd__clkbuf_8
XFILLER_128_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload152 clknet_leaf_305_clk VGND VGND VPWR VPWR clkload152/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload163 clknet_leaf_224_clk VGND VGND VPWR VPWR clkload163/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23071_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[1\]\[1\]
+ VGND VGND VPWR VPWR _09743_ sky130_fd_sc_hd__and2_1
XFILLER_150_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload174 clknet_leaf_195_clk VGND VGND VPWR VPWR clkload174/Y sky130_fd_sc_hd__bufinv_16
X_20283_ _07201_ _07204_ _07222_ _07223_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__a211o_1
Xclkload185 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload185/Y sky130_fd_sc_hd__inv_8
XFILLER_115_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload196 clknet_leaf_55_clk VGND VGND VPWR VPWR clkload196/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_129_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22022_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[23\]
+ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__xor2_1
XFILLER_161_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_222_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26830_ clknet_leaf_87_clk _00632_ net153 VGND VGND VPWR VPWR B_in\[102\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_222_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26761_ clknet_leaf_77_clk _00563_ net143 VGND VGND VPWR VPWR B_in\[33\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23973_ systolic_inst.B_shift\[13\]\[6\] B_in\[46\] _00008_ VGND VGND VPWR VPWR _10512_
+ sky130_fd_sc_hd__mux2_1
XFILLER_99_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28500_ clknet_leaf_112_clk _02298_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_25712_ systolic_inst.acc_wires\[5\]\[28\] C_out\[188\] net46 VGND VGND VPWR VPWR
+ _03014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_235_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22924_ _09601_ _09602_ VGND VGND VPWR VPWR _09603_ sky130_fd_sc_hd__nand2_1
X_29480_ clknet_leaf_271_clk _03278_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_235_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26692_ clknet_leaf_1_B_in_serial_clk _00495_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28431_ clknet_leaf_26_clk _02229_ VGND VGND VPWR VPWR systolic_inst.A_shift\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25643_ systolic_inst.acc_wires\[3\]\[23\] C_out\[119\] net50 VGND VGND VPWR VPWR
+ _02945_ sky130_fd_sc_hd__mux2_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22855_ systolic_inst.B_outs\[1\]\[7\] _09429_ _09461_ _09497_ VGND VGND VPWR VPWR
+ _09536_ sky130_fd_sc_hd__o31a_1
XFILLER_231_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21806_ _08544_ _08548_ _08577_ _08576_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__o31a_1
X_28362_ clknet_leaf_68_clk _02160_ VGND VGND VPWR VPWR systolic_inst.B_shift\[22\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25574_ systolic_inst.acc_wires\[1\]\[18\] C_out\[50\] net35 VGND VGND VPWR VPWR
+ _02876_ sky130_fd_sc_hd__mux2_1
X_22786_ _09466_ _09467_ _09456_ VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__a21o_1
XFILLER_231_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27313_ clknet_leaf_293_clk _01111_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24525_ C_out\[89\] net100 net82 ser_C.shift_reg\[89\] _10732_ VGND VGND VPWR VPWR
+ _02339_ sky130_fd_sc_hd__a221o_1
X_21737_ _08542_ _08543_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__nor2_1
XFILLER_227_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28293_ clknet_leaf_99_clk _02091_ VGND VGND VPWR VPWR systolic_inst.B_shift\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27244_ clknet_leaf_274_clk _01042_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24456_ net114 ser_C.shift_reg\[56\] VGND VGND VPWR VPWR _10698_ sky130_fd_sc_hd__and2_1
X_21668_ _08476_ _08475_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__and2b_1
XFILLER_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23407_ _09991_ _10031_ VGND VGND VPWR VPWR _10033_ sky130_fd_sc_hd__xnor2_1
X_20619_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[5\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__a21o_1
X_24387_ C_out\[20\] net104 _10643_ ser_C.shift_reg\[20\] _10663_ VGND VGND VPWR VPWR
+ _02270_ sky130_fd_sc_hd__a221o_1
X_27175_ clknet_leaf_255_clk _00973_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_21599_ _08404_ _08408_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__nor2_1
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14140_ net118 systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[0\] VGND
+ VGND VPWR VPWR _11334_ sky130_fd_sc_hd__and3_1
X_26126_ deser_B.serial_word\[81\] deser_B.shift_reg\[81\] net55 VGND VGND VPWR VPWR
+ _03428_ sky130_fd_sc_hd__mux2_1
X_23338_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[5\]
+ systolic_inst.A_outs\[0\]\[5\] VGND VGND VPWR VPWR _09966_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_10_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14071_ deser_B.shift_reg\[105\] deser_B.shift_reg\[106\] net126 VGND VGND VPWR VPWR
+ _00897_ sky130_fd_sc_hd__mux2_1
X_23269_ _09910_ _09911_ VGND VGND VPWR VPWR _09912_ sky130_fd_sc_hd__nand2_1
X_26057_ deser_B.serial_word\[12\] deser_B.shift_reg\[12\] net55 VGND VGND VPWR VPWR
+ _03359_ sky130_fd_sc_hd__mux2_1
XFILLER_153_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25008_ net111 ser_C.shift_reg\[332\] VGND VGND VPWR VPWR _10974_ sky130_fd_sc_hd__and2_1
XFILLER_239_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17830_ _05025_ _05026_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__xnor2_1
XFILLER_239_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_210_Right_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17761_ systolic_inst.acc_wires\[10\]\[26\] systolic_inst.acc_wires\[10\]\[27\] systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__o21a_1
X_14973_ _12093_ _12092_ VGND VGND VPWR VPWR _12094_ sky130_fd_sc_hd__nand2b_1
XFILLER_48_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26959_ clknet_leaf_2_A_in_serial_clk _00757_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19500_ _06528_ _06536_ _06542_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__o21ai_1
XFILLER_43_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16712_ systolic_inst.A_outs\[11\]\[1\] systolic_inst.B_outs\[11\]\[6\] _04033_ VGND
+ VGND VPWR VPWR _04034_ sky130_fd_sc_hd__and3_1
X_13924_ deser_A.serial_word\[85\] deser_A.shift_reg\[85\] net57 VGND VGND VPWR VPWR
+ _00750_ sky130_fd_sc_hd__mux2_1
X_29678_ clknet_leaf_33_B_in_serial_clk _03473_ net134 VGND VGND VPWR VPWR deser_B.serial_word\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_17692_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[17\]
+ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__xor2_2
XFILLER_212_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19431_ _06483_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__inv_2
XFILLER_63_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28629_ clknet_leaf_207_clk _02427_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[177\]
+ sky130_fd_sc_hd__dfrtp_1
X_16643_ _03965_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__nor2_1
XFILLER_223_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13855_ deser_A.serial_word\[16\] deser_A.shift_reg\[16\] net58 VGND VGND VPWR VPWR
+ _00681_ sky130_fd_sc_hd__mux2_1
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19362_ _06419_ _06420_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__and2b_1
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16574_ net108 systolic_inst.acc_wires\[12\]\[31\] net67 _03919_ VGND VGND VPWR VPWR
+ _01201_ sky130_fd_sc_hd__a22o_1
XFILLER_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13786_ B_in\[93\] deser_B.word_buffer\[93\] net89 VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__mux2_1
XFILLER_204_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18313_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[18\]
+ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__nand2_1
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15525_ systolic_inst.B_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[5\]
+ systolic_inst.B_outs\[13\]\[3\] VGND VGND VPWR VPWR _12583_ sky130_fd_sc_hd__a22oi_1
XFILLER_163_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19293_ _06354_ _06353_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__nand2b_1
XFILLER_43_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18244_ _05414_ _05417_ _05420_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__nand3_1
XFILLER_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15456_ systolic_inst.B_outs\[13\]\[3\] systolic_inst.A_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\]
+ systolic_inst.A_outs\[13\]\[2\] VGND VGND VPWR VPWR _12516_ sky130_fd_sc_hd__a22o_1
XFILLER_204_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _11588_ _11589_ VGND VGND VPWR VPWR _11590_ sky130_fd_sc_hd__or2_1
XFILLER_89_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18175_ _05290_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__xnor2_1
XFILLER_191_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15387_ systolic_inst.A_outs\[13\]\[1\] systolic_inst.B_outs\[13\]\[2\] systolic_inst.B_outs\[13\]\[3\]
+ systolic_inst.A_outs\[13\]\[0\] VGND VGND VPWR VPWR _12450_ sky130_fd_sc_hd__a22oi_1
XFILLER_204_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17126_ _04407_ _04411_ _04414_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__a21o_1
XFILLER_15_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14338_ _11521_ _11522_ VGND VGND VPWR VPWR _11523_ sky130_fd_sc_hd__or2_1
XFILLER_171_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17057_ _04351_ _04355_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_165_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14269_ _11452_ _11455_ VGND VGND VPWR VPWR _11456_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_111_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16008_ systolic_inst.A_outs\[12\]\[1\] systolic_inst.B_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\]
+ systolic_inst.A_outs\[12\]\[0\] VGND VGND VPWR VPWR _13006_ sky130_fd_sc_hd__a22o_1
XFILLER_125_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17959_ _05151_ _05148_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__and2b_1
XFILLER_22_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20970_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[5\] VGND VGND VPWR
+ VPWR _07844_ sky130_fd_sc_hd__nand2_1
XFILLER_226_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19629_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[0\] _06637_
+ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__a21o_1
XFILLER_241_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22640_ systolic_inst.acc_wires\[2\]\[24\] systolic_inst.acc_wires\[2\]\[25\] systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__o21a_1
XFILLER_202_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_230_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22571_ _09285_ _09290_ _09291_ _09292_ VGND VGND VPWR VPWR _09293_ sky130_fd_sc_hd__a211o_1
XFILLER_146_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_118_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21522_ _08314_ _08333_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24310_ _10628_ systolic_inst.A_shift\[10\]\[2\] net70 VGND VGND VPWR VPWR _02228_
+ sky130_fd_sc_hd__mux2_1
XFILLER_210_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25290_ net111 ser_C.shift_reg\[473\] VGND VGND VPWR VPWR _11115_ sky130_fd_sc_hd__and2_1
XFILLER_221_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24241_ systolic_inst.A_shift\[19\]\[4\] A_in\[68\] net59 VGND VGND VPWR VPWR _10606_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21453_ _08278_ _08281_ _08284_ _08287_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__o31a_1
XFILLER_222_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20404_ _07337_ _07339_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_21_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24172_ systolic_inst.A_shift\[26\]\[3\] net70 _10505_ systolic_inst.A_shift\[27\]\[3\]
+ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__a22o_1
X_21384_ _08222_ _08226_ _08228_ _11713_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__a31o_1
XFILLER_107_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23123_ _09787_ _09786_ systolic_inst.acc_wires\[1\]\[8\] net109 VGND VGND VPWR VPWR
+ _01882_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_224_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20335_ _07271_ _07272_ _07241_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_224_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28980_ clknet_leaf_24_clk _02778_ VGND VGND VPWR VPWR systolic_inst.A_shift\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_224_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23054_ _09654_ _09703_ _09702_ VGND VGND VPWR VPWR _09729_ sky130_fd_sc_hd__o21ba_1
X_27931_ clknet_leaf_136_clk _01729_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_20266_ net109 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[3\] VGND
+ VGND VPWR VPWR _07208_ sky130_fd_sc_hd__nand2_1
XFILLER_192_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22005_ _08759_ _08763_ _08785_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27862_ clknet_leaf_215_clk _01660_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_20197_ net106 systolic_inst.acc_wires\[6\]\[27\] net62 _07162_ VGND VGND VPWR VPWR
+ _01581_ sky130_fd_sc_hd__a22o_1
XFILLER_62_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29601_ clknet_leaf_18_B_in_serial_clk _03396_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_26813_ clknet_leaf_55_clk _00615_ net144 VGND VGND VPWR VPWR B_in\[85\] sky130_fd_sc_hd__dfrtp_1
XFILLER_153_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27793_ clknet_leaf_42_clk _01591_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_5_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29532_ clknet_leaf_259_clk _03330_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[504\]
+ sky130_fd_sc_hd__dfrtp_1
X_26744_ clknet_leaf_125_clk _00546_ net144 VGND VGND VPWR VPWR B_in\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_229_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23956_ systolic_inst.B_shift\[11\]\[3\] net71 net83 systolic_inst.B_shift\[15\]\[3\]
+ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__a22o_1
XFILLER_57_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22907_ _09515_ _09585_ VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__nor2_1
X_29463_ clknet_leaf_331_clk _03261_ net136 VGND VGND VPWR VPWR C_out\[435\] sky130_fd_sc_hd__dfrtp_1
X_26675_ clknet_leaf_9_B_in_serial_clk _00478_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23887_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[30\]
+ VGND VGND VPWR VPWR _10474_ sky130_fd_sc_hd__or2_1
XFILLER_44_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28414_ clknet_leaf_63_clk _02212_ VGND VGND VPWR VPWR systolic_inst.B_shift\[23\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13640_ deser_B.word_buffer\[76\] deser_B.serial_word\[76\] net123 VGND VGND VPWR
+ VPWR _00477_ sky130_fd_sc_hd__mux2_1
X_25626_ systolic_inst.acc_wires\[3\]\[6\] C_out\[102\] net48 VGND VGND VPWR VPWR
+ _02928_ sky130_fd_sc_hd__mux2_1
X_22838_ _09514_ _09517_ VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__xnor2_1
X_29394_ clknet_leaf_235_clk _03192_ net145 VGND VGND VPWR VPWR C_out\[366\] sky130_fd_sc_hd__dfrtp_1
XFILLER_112_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28345_ clknet_leaf_343_clk _02143_ VGND VGND VPWR VPWR systolic_inst.A_shift\[25\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_25557_ systolic_inst.acc_wires\[1\]\[1\] C_out\[33\] net36 VGND VGND VPWR VPWR _02859_
+ sky130_fd_sc_hd__mux2_1
X_13571_ deser_B.word_buffer\[7\] deser_B.serial_word\[7\] net124 VGND VGND VPWR VPWR
+ _00408_ sky130_fd_sc_hd__mux2_1
XFILLER_188_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22769_ _09450_ _09451_ VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__or2_1
XFILLER_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_160_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15310_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[24\]
+ VGND VGND VPWR VPWR _12400_ sky130_fd_sc_hd__nor2_1
XFILLER_40_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24508_ net112 ser_C.shift_reg\[82\] VGND VGND VPWR VPWR _10724_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_213_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28276_ clknet_leaf_123_clk _02074_ VGND VGND VPWR VPWR systolic_inst.B_shift\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16290_ _03639_ _03641_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__a21o_1
X_25488_ systolic_inst.cycle_cnt\[18\] _11220_ VGND VGND VPWR VPWR _11223_ sky130_fd_sc_hd__and2_1
XFILLER_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15241_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[14\]\[14\]
+ VGND VGND VPWR VPWR _12341_ sky130_fd_sc_hd__nand2_1
XFILLER_36_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27227_ clknet_leaf_326_clk _01025_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_24439_ C_out\[46\] _11302_ net81 ser_C.shift_reg\[46\] _10689_ VGND VGND VPWR VPWR
+ _02296_ sky130_fd_sc_hd__a221o_1
XFILLER_201_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15172_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[14\]\[4\]
+ VGND VGND VPWR VPWR _12282_ sky130_fd_sc_hd__or2_1
X_27158_ clknet_leaf_296_clk _00956_ net138 VGND VGND VPWR VPWR systolic_inst.B_outs\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_67_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26109_ deser_B.serial_word\[64\] deser_B.shift_reg\[64\] net56 VGND VGND VPWR VPWR
+ _03411_ sky130_fd_sc_hd__mux2_1
X_14123_ systolic_inst.A_shift\[21\]\[7\] net71 _11333_ A_in\[95\] VGND VGND VPWR
+ VPWR _00945_ sky130_fd_sc_hd__a22o_1
XFILLER_236_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19980_ _06974_ _06975_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27089_ clknet_leaf_1_B_in_serial_clk _00887_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_125_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18931_ _06026_ _06030_ _06032_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__a21oi_1
X_14054_ deser_B.shift_reg\[88\] deser_B.shift_reg\[89\] net125 VGND VGND VPWR VPWR
+ _00880_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18862_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[8\]\[10\]
+ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_160_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17813_ systolic_inst.A_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[2\] VGND VGND VPWR
+ VPWR _05012_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_24_B_in_serial_clk clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_24_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_121_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18793_ _05833_ _05896_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17744_ _04968_ _04967_ systolic_inst.acc_wires\[10\]\[24\] net105 VGND VGND VPWR
+ VPWR _01322_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_208_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14956_ systolic_inst.B_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[5\]
+ systolic_inst.A_outs\[14\]\[6\] VGND VGND VPWR VPWR _12077_ sky130_fd_sc_hd__and4_1
XFILLER_36_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13907_ deser_A.serial_word\[68\] deser_A.shift_reg\[68\] net57 VGND VGND VPWR VPWR
+ _00733_ sky130_fd_sc_hd__mux2_1
X_17675_ _04906_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__nand2_1
X_14887_ _12006_ _12009_ VGND VGND VPWR VPWR _12010_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_158_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19414_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[7\]\[2\]
+ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__or2_1
XFILLER_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16626_ systolic_inst.A_outs\[11\]\[4\] _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__nand2_1
X_13838_ _00001_ _11321_ _11329_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_158_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap90 _00005_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_6
XFILLER_189_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19345_ systolic_inst.A_outs\[7\]\[6\] _11261_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_100_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16557_ _03902_ _03904_ _03905_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13769_ B_in\[76\] deser_B.word_buffer\[76\] net90 VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__mux2_1
XFILLER_189_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_42_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15508_ _12538_ _12566_ VGND VGND VPWR VPWR _12567_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_61_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19276_ _06299_ _06337_ _06336_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__a21oi_2
XFILLER_203_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16488_ _03843_ _03845_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_61_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18227_ _05406_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__inv_2
X_15439_ _12475_ _12498_ VGND VGND VPWR VPWR _12500_ sky130_fd_sc_hd__xor2_1
XFILLER_54_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18158_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[13\] _05344_
+ _05345_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__a22o_1
XFILLER_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17109_ net62 _04400_ _04401_ systolic_inst.acc_wires\[11\]\[20\] net105 VGND VGND
+ VPWR VPWR _01254_ sky130_fd_sc_hd__a32o_1
XFILLER_190_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18089_ _05276_ _05277_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__and2b_1
XFILLER_102_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20120_ _07097_ _07096_ systolic_inst.acc_wires\[6\]\[15\] net106 VGND VGND VPWR
+ VPWR _01569_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20051_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[6\]\[6\]
+ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__nand2_1
XFILLER_219_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23810_ _11258_ systolic_inst.acc_wires\[0\]\[17\] net64 _10409_ VGND VGND VPWR VPWR
+ _01947_ sky130_fd_sc_hd__a22o_1
XFILLER_113_1251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24790_ net113 ser_C.shift_reg\[223\] VGND VGND VPWR VPWR _10865_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23741_ net63 _10349_ _10350_ systolic_inst.acc_wires\[0\]\[7\] _11258_ VGND VGND
+ VPWR VPWR _01937_ sky130_fd_sc_hd__a32o_1
XFILLER_113_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20953_ _07826_ _07827_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__and2_1
XFILLER_226_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_217_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_217_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26460_ clknet_leaf_1_A_in_serial_clk _00267_ net132 VGND VGND VPWR VPWR deser_A.bit_idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23672_ _10286_ _10290_ VGND VGND VPWR VPWR _10291_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20884_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[4\] _07757_ _07759_
+ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__a22oi_1
Xclkbuf_2_2__f_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_2_2__leaf_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_148_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25411_ systolic_inst.A_shift\[2\]\[5\] A_in\[13\] net59 VGND VGND VPWR VPWR _11175_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22623_ _09316_ _09322_ _09327_ _09333_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__nand4_1
XFILLER_228_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26391_ clknet_leaf_16_clk _00198_ net132 VGND VGND VPWR VPWR A_in\[59\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_33_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
X_28130_ clknet_leaf_100_clk _01928_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22554_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[2\]\[13\]
+ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__xor2_1
X_25342_ net112 ser_C.shift_reg\[499\] VGND VGND VPWR VPWR _11141_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_23_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21505_ _08312_ _08318_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__or2_1
X_28061_ clknet_leaf_121_clk _01859_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22485_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[2\]\[3\]
+ VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__nand2_1
X_25273_ ser_C.parallel_data\[463\] net102 net74 ser_C.shift_reg\[463\] _11106_ VGND
+ VGND VPWR VPWR _02713_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_101_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27012_ clknet_leaf_21_B_in_serial_clk _00810_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_108_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21436_ _08267_ _08271_ _08268_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__a21bo_1
X_24224_ _10597_ systolic_inst.A_shift\[19\]\[3\] net70 VGND VGND VPWR VPWR _02173_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24155_ systolic_inst.A_shift\[28\]\[1\] A_in\[97\] net59 VGND VGND VPWR VPWR _10579_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21367_ _08211_ _08214_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__nor2_1
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23106_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[1\]\[6\]
+ VGND VGND VPWR VPWR _09773_ sky130_fd_sc_hd__nand2_1
X_20318_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[5\]
+ systolic_inst.A_outs\[5\]\[6\] VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__and4_1
X_24086_ systolic_inst.B_shift\[2\]\[5\] _11332_ net83 systolic_inst.B_shift\[6\]\[5\]
+ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__a22o_1
X_28963_ clknet_leaf_246_clk _02761_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[511\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21298_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[4\]\[7\]
+ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__or2_1
XFILLER_150_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23037_ net122 _09710_ _09711_ _09712_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__a31o_1
X_27914_ clknet_leaf_134_clk _01712_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_20249_ _07189_ _07190_ _07185_ VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__or3b_1
XFILLER_66_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28894_ clknet_leaf_286_clk _02692_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27845_ clknet_leaf_181_clk _01643_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_110_Left_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_202_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[5\]
+ systolic_inst.B_outs\[14\]\[0\] VGND VGND VPWR VPWR _11935_ sky130_fd_sc_hd__a22oi_1
XFILLER_92_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_202_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27776_ clknet_leaf_177_clk _01574_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
X_15790_ _12827_ _12828_ _12826_ VGND VGND VPWR VPWR _12834_ sky130_fd_sc_hd__a21bo_1
X_24988_ net111 ser_C.shift_reg\[322\] VGND VGND VPWR VPWR _10964_ sky130_fd_sc_hd__and2_1
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29515_ clknet_leaf_254_clk _03313_ net140 VGND VGND VPWR VPWR ser_C.parallel_data\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26727_ clknet_leaf_7_B_in_serial_clk _00529_ net5 VGND VGND VPWR VPWR deser_B.serial_toggle
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14741_ systolic_inst.A_outs\[14\]\[1\] systolic_inst.A_outs\[13\]\[1\] net120 VGND
+ VGND VPWR VPWR _01011_ sky130_fd_sc_hd__mux2_1
XFILLER_229_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23939_ _10498_ systolic_inst.B_shift\[10\]\[1\] _11332_ VGND VGND VPWR VPWR _01987_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_194_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_194_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29446_ clknet_leaf_300_clk _03244_ net139 VGND VGND VPWR VPWR C_out\[418\] sky130_fd_sc_hd__dfrtp_1
X_17460_ _04643_ _04713_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__xnor2_4
XFILLER_229_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26658_ clknet_leaf_30_B_in_serial_clk _00461_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_14672_ _11820_ _11826_ _11827_ VGND VGND VPWR VPWR _11829_ sky130_fd_sc_hd__a21oi_1
XFILLER_233_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16411_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[12\]\[7\]
+ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__or2_1
X_25609_ systolic_inst.acc_wires\[2\]\[21\] C_out\[85\] net52 VGND VGND VPWR VPWR
+ _02911_ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_13623_ deser_B.word_buffer\[59\] deser_B.serial_word\[59\] net124 VGND VGND VPWR
+ VPWR _00460_ sky130_fd_sc_hd__mux2_1
XFILLER_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29377_ clknet_leaf_244_clk _03175_ net145 VGND VGND VPWR VPWR C_out\[349\] sky130_fd_sc_hd__dfrtp_1
X_17391_ _04643_ _04646_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__xnor2_1
XFILLER_242_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26589_ clknet_leaf_30_A_in_serial_clk _00392_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[119\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_24_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_13_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19130_ _06166_ _06196_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__xnor2_1
X_16342_ _03694_ _03697_ _03719_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__and3_1
X_28328_ clknet_leaf_0_clk _02126_ VGND VGND VPWR VPWR systolic_inst.A_shift\[27\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13554_ deser_A.shift_reg\[118\] deser_A.shift_reg\[119\] net130 VGND VGND VPWR VPWR
+ _00391_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19061_ systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[3\] systolic_inst.A_outs\[7\]\[4\]
+ systolic_inst.B_outs\[7\]\[0\] VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__a22o_1
X_28259_ clknet_leaf_98_clk _02057_ VGND VGND VPWR VPWR systolic_inst.B_shift\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16273_ _03620_ _03624_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__and2_1
XFILLER_199_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13485_ deser_A.shift_reg\[49\] deser_A.shift_reg\[50\] net130 VGND VGND VPWR VPWR
+ _00322_ sky130_fd_sc_hd__mux2_1
XFILLER_201_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18012_ _05195_ _05203_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__xnor2_1
X_15224_ _12316_ _12321_ _12322_ VGND VGND VPWR VPWR _12326_ sky130_fd_sc_hd__nand3_1
XFILLER_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15155_ _11712_ _12266_ _12267_ systolic_inst.acc_wires\[14\]\[1\] net107 VGND VGND
+ VPWR VPWR _01043_ sky130_fd_sc_hd__a32o_1
XFILLER_236_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14106_ systolic_inst.A_shift\[12\]\[6\] net71 _11333_ A_in\[62\] VGND VGND VPWR
+ VPWR _00928_ sky130_fd_sc_hd__a22o_1
XFILLER_181_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19963_ _06956_ _06957_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__xnor2_1
X_15086_ _12201_ _12202_ VGND VGND VPWR VPWR _12204_ sky130_fd_sc_hd__xor2_1
XFILLER_99_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14037_ deser_B.shift_reg\[71\] deser_B.shift_reg\[72\] net126 VGND VGND VPWR VPWR
+ _00863_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18914_ _06014_ _06017_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__nor2_1
X_19894_ _06890_ _06891_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__nand2_1
XFILLER_80_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18845_ _05952_ _05954_ _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__nand3_1
XFILLER_45_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18776_ _05871_ _05873_ _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__a21oi_1
XFILLER_227_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15988_ systolic_inst.A_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[2\] _12986_ VGND
+ VGND VPWR VPWR _12988_ sky130_fd_sc_hd__a21o_1
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17727_ _04952_ _04953_ _04951_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__o21ai_1
X_14939_ _12059_ _12060_ VGND VGND VPWR VPWR _12061_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_102_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17658_ _04892_ _04893_ _04894_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__and3_1
XFILLER_235_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16609_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[2\]
+ systolic_inst.A_outs\[11\]\[3\] VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__nand4_2
XFILLER_56_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17589_ _04832_ _04833_ _04834_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__and3_1
XFILLER_91_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_17_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19328_ _06376_ _06388_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19259_ _06312_ _06320_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__or2_1
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22270_ _09013_ _09014_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__xor2_1
XFILLER_178_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21221_ _11258_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[14\] VGND
+ VGND VPWR VPWR _08088_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_132_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21152_ _07976_ _07979_ _08019_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_93_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20103_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[6\]\[12\]
+ _07079_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_242_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21083_ systolic_inst.B_outs\[4\]\[4\] systolic_inst.A_outs\[4\]\[6\] systolic_inst.A_outs\[4\]\[7\]
+ systolic_inst.B_outs\[4\]\[3\] VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__a22o_1
X_25960_ systolic_inst.acc_wires\[13\]\[20\] C_out\[436\] net20 VGND VGND VPWR VPWR
+ _03262_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20034_ _07020_ _07021_ _07022_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__and3_1
X_24911_ C_out\[282\] net103 net75 ser_C.shift_reg\[282\] _10925_ VGND VGND VPWR VPWR
+ _02532_ sky130_fd_sc_hd__a221o_1
XFILLER_113_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25891_ systolic_inst.acc_wires\[11\]\[15\] C_out\[367\] net40 VGND VGND VPWR VPWR
+ _03193_ sky130_fd_sc_hd__mux2_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_219_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_219_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27630_ clknet_leaf_323_clk _01428_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24842_ net113 ser_C.shift_reg\[249\] VGND VGND VPWR VPWR _10891_ sky130_fd_sc_hd__and2_1
XFILLER_150_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27561_ clknet_leaf_305_clk _01359_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_24773_ C_out\[213\] net98 net78 ser_C.shift_reg\[213\] _10856_ VGND VGND VPWR VPWR
+ _02463_ sky130_fd_sc_hd__a221o_1
XFILLER_113_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21985_ _08768_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__inv_2
XFILLER_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29300_ clknet_leaf_312_clk _03098_ net142 VGND VGND VPWR VPWR C_out\[272\] sky130_fd_sc_hd__dfrtp_1
X_26512_ clknet_leaf_11_A_in_serial_clk _00315_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_23724_ _10329_ _10330_ _10328_ VGND VGND VPWR VPWR _10336_ sky130_fd_sc_hd__a21bo_1
X_27492_ clknet_leaf_227_clk _01290_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_20936_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[5\]
+ systolic_inst.B_outs\[4\]\[5\] VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__nand4_1
XFILLER_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29231_ clknet_leaf_204_clk _03029_ net147 VGND VGND VPWR VPWR C_out\[203\] sky130_fd_sc_hd__dfrtp_1
X_26443_ clknet_leaf_347_clk _00250_ net132 VGND VGND VPWR VPWR A_in\[111\] sky130_fd_sc_hd__dfrtp_1
X_23655_ _10238_ _10241_ _10273_ VGND VGND VPWR VPWR _10275_ sky130_fd_sc_hd__and3_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20867_ _07742_ _07743_ _07731_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__a21o_1
XFILLER_242_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22606_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[21\]
+ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__xor2_1
XFILLER_70_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29162_ clknet_leaf_309_clk _02960_ net142 VGND VGND VPWR VPWR C_out\[134\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26374_ clknet_leaf_23_clk _00181_ net133 VGND VGND VPWR VPWR A_in\[42\] sky130_fd_sc_hd__dfrtp_1
XFILLER_224_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20798_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[27\]
+ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__xnor2_1
X_23586_ _10191_ _10207_ VGND VGND VPWR VPWR _10208_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28113_ clknet_leaf_47_clk _01911_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_25325_ ser_C.parallel_data\[489\] net97 net77 ser_C.shift_reg\[489\] _11132_ VGND
+ VGND VPWR VPWR _02739_ sky130_fd_sc_hd__a221o_1
X_29093_ clknet_leaf_112_clk _02891_ net150 VGND VGND VPWR VPWR C_out\[65\] sky130_fd_sc_hd__dfrtp_1
X_22537_ net109 systolic_inst.acc_wires\[2\]\[10\] net65 _09263_ VGND VGND VPWR VPWR
+ _01820_ sky130_fd_sc_hd__a22o_1
XFILLER_195_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28044_ clknet_leaf_127_clk _01842_ net144 VGND VGND VPWR VPWR systolic_inst.A_outs\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_139_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25256_ net111 ser_C.shift_reg\[456\] VGND VGND VPWR VPWR _11098_ sky130_fd_sc_hd__and2_1
X_13270_ deser_A.word_buffer\[108\] deser_A.serial_word\[108\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__mux2_1
XFILLER_108_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22468_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[2\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__a21o_1
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24207_ systolic_inst.A_shift\[21\]\[3\] A_in\[83\] net59 VGND VGND VPWR VPWR _10589_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_187_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21419_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[24\]
+ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__and2_1
X_22399_ _09126_ _09139_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__xnor2_1
X_25187_ C_out\[420\] net102 net74 ser_C.shift_reg\[420\] _11063_ VGND VGND VPWR VPWR
+ _02670_ sky130_fd_sc_hd__a221o_1
XFILLER_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_208_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24138_ _10570_ systolic_inst.A_shift\[28\]\[0\] net70 VGND VGND VPWR VPWR _02114_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16960_ _04271_ _04273_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_204_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24069_ systolic_inst.B_shift\[19\]\[6\] B_in\[30\] net59 VGND VGND VPWR VPWR _10552_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28946_ clknet_leaf_258_clk _02744_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[494\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_133_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15911_ systolic_inst.acc_wires\[13\]\[20\] systolic_inst.acc_wires\[13\]\[21\] systolic_inst.acc_wires\[13\]\[22\]
+ systolic_inst.acc_wires\[13\]\[23\] systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12937_ sky130_fd_sc_hd__o41a_1
XFILLER_77_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28877_ clknet_leaf_290_clk _02675_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[425\]
+ sky130_fd_sc_hd__dfrtp_1
X_16891_ _04205_ _04206_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__xnor2_1
XFILLER_237_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_188_Right_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18630_ _05719_ _05721_ _05756_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__and3_1
X_27828_ clknet_leaf_140_clk _01626_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15842_ _12874_ _12876_ _12878_ systolic_inst.acc_wires\[13\]\[13\] net108 VGND VGND
+ VPWR VPWR _01119_ sky130_fd_sc_hd__a32o_1
XFILLER_237_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18561_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[7\] _05690_ net115
+ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__mux2_1
X_27759_ clknet_leaf_211_clk _01557_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15773_ net66 _12817_ _12819_ systolic_inst.acc_wires\[13\]\[3\] net107 VGND VGND
+ VPWR VPWR _01109_ sky130_fd_sc_hd__a32o_1
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17512_ _04763_ _04764_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__or2_1
XFILLER_206_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14724_ _11872_ VGND VGND VPWR VPWR _11873_ sky130_fd_sc_hd__inv_2
XFILLER_217_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18492_ _05621_ _05622_ net115 VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__o21a_1
XFILLER_220_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29429_ clknet_leaf_344_clk _03227_ net131 VGND VGND VPWR VPWR C_out\[401\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17443_ _04640_ _04696_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__or2_1
X_14655_ _11812_ _11814_ VGND VGND VPWR VPWR _11815_ sky130_fd_sc_hd__xor2_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13606_ deser_B.word_buffer\[42\] deser_B.serial_word\[42\] net123 VGND VGND VPWR
+ VPWR _00443_ sky130_fd_sc_hd__mux2_1
XFILLER_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17374_ _04590_ _04592_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__nor2_1
X_14586_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[15\]\[8\]
+ _11752_ _11754_ VGND VGND VPWR VPWR _11755_ sky130_fd_sc_hd__a211o_1
X_19113_ systolic_inst.A_outs\[7\]\[1\] systolic_inst.B_outs\[7\]\[5\] systolic_inst.B_outs\[7\]\[6\]
+ systolic_inst.A_outs\[7\]\[0\] VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__a22oi_1
XFILLER_9_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16325_ _03704_ _03703_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__and2b_1
XFILLER_229_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13537_ deser_A.shift_reg\[101\] deser_A.shift_reg\[102\] net129 VGND VGND VPWR VPWR
+ _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_173_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19044_ _06112_ _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__nor2_1
XFILLER_118_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16256_ _03597_ _03599_ _03598_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__o21ba_1
X_13468_ deser_A.shift_reg\[32\] deser_A.shift_reg\[33\] deser_A.receiving VGND VGND
+ VPWR VPWR _00305_ sky130_fd_sc_hd__mux2_1
XFILLER_199_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15207_ _12305_ _12308_ VGND VGND VPWR VPWR _12312_ sky130_fd_sc_hd__and2_1
XFILLER_173_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16187_ _03570_ _03569_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__nand2b_1
X_13399_ A_in\[108\] deser_A.word_buffer\[108\] _00003_ VGND VGND VPWR VPWR _00247_
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15138_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[14\] _12251_
+ _12253_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__a22o_1
XFILLER_173_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_206_Left_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19946_ _06854_ _06912_ _06911_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__a21oi_1
X_15069_ _12146_ _12186_ VGND VGND VPWR VPWR _12187_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_4_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19877_ _06824_ _06841_ _06839_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__o21a_1
XFILLER_96_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18828_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__inv_2
XFILLER_3_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18759_ _05881_ _05882_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__nor2_1
XFILLER_224_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21770_ _08575_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__inv_2
XFILLER_36_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20721_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[15\]
+ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__and2_1
XFILLER_93_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_215_Left_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_A_in_serial_clk clknet_2_0__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_30_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_212_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23440_ _10034_ _10036_ _10035_ VGND VGND VPWR VPWR _10065_ sky130_fd_sc_hd__o21ba_1
X_20652_ _07569_ _07570_ _07568_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__a21bo_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23371_ systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[6\] VGND VGND VPWR
+ VPWR _09998_ sky130_fd_sc_hd__nand2_1
XFILLER_143_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20583_ _07481_ _07483_ _07513_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__or3_1
XFILLER_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_18__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_18__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_108_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25110_ net112 ser_C.shift_reg\[383\] VGND VGND VPWR VPWR _11025_ sky130_fd_sc_hd__and2_1
XFILLER_191_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22322_ systolic_inst.A_outs\[2\]\[4\] systolic_inst.B_outs\[2\]\[6\] _11265_ systolic_inst.A_outs\[2\]\[3\]
+ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_95_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26090_ deser_B.serial_word\[45\] deser_B.shift_reg\[45\] net55 VGND VGND VPWR VPWR
+ _03392_ sky130_fd_sc_hd__mux2_1
XFILLER_137_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22253_ _08996_ _08997_ VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__nor2_1
XFILLER_152_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25041_ C_out\[347\] net97 net77 ser_C.shift_reg\[347\] _10990_ VGND VGND VPWR VPWR
+ _02597_ sky130_fd_sc_hd__a221o_1
XFILLER_219_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21204_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[7\] _08039_ _07884_
+ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__a31o_1
XFILLER_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_224_Left_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22184_ _08925_ _08926_ _08930_ VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_240_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_240_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21135_ systolic_inst.A_outs\[4\]\[5\] systolic_inst.B_outs\[4\]\[6\] _08003_ VGND
+ VGND VPWR VPWR _08005_ sky130_fd_sc_hd__a21oi_1
X_28800_ clknet_leaf_240_clk _02598_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[348\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_219_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26992_ clknet_leaf_0_A_in_serial_clk _00790_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28731_ clknet_leaf_291_clk _02529_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[279\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_115_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21066_ _07935_ _07936_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__xor2_1
X_25943_ systolic_inst.acc_wires\[13\]\[3\] C_out\[419\] net14 VGND VGND VPWR VPWR
+ _03245_ sky130_fd_sc_hd__mux2_1
XFILLER_59_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20017_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[6\]\[1\]
+ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__nand2_1
XFILLER_115_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28662_ clknet_leaf_177_clk _02460_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[210\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25874_ systolic_inst.acc_wires\[10\]\[30\] C_out\[350\] net41 VGND VGND VPWR VPWR
+ _03176_ sky130_fd_sc_hd__mux2_1
XFILLER_100_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27613_ clknet_leaf_321_clk _01411_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24825_ C_out\[239\] net99 net79 ser_C.shift_reg\[239\] _10882_ VGND VGND VPWR VPWR
+ _02489_ sky130_fd_sc_hd__a221o_1
XFILLER_98_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28593_ clknet_leaf_42_clk _02391_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[141\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_238_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_233_Left_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27544_ clknet_leaf_34_clk _01342_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_24756_ net113 ser_C.shift_reg\[206\] VGND VGND VPWR VPWR _10848_ sky130_fd_sc_hd__and2_1
X_21968_ _08752_ _08753_ VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23707_ net63 _10319_ _10321_ systolic_inst.acc_wires\[0\]\[2\] _11258_ VGND VGND
+ VPWR VPWR _01932_ sky130_fd_sc_hd__a32o_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20919_ systolic_inst.B_outs\[4\]\[3\] _07729_ _07769_ _07767_ VGND VGND VPWR VPWR
+ _07795_ sky130_fd_sc_hd__a31o_1
X_27475_ clknet_leaf_220_clk _01273_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_24687_ C_out\[170\] net104 net76 ser_C.shift_reg\[170\] _10813_ VGND VGND VPWR VPWR
+ _02420_ sky130_fd_sc_hd__a221o_1
XFILLER_226_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21899_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[3\]\[5\]
+ VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__nand2_1
X_29214_ clknet_leaf_179_clk _03012_ net148 VGND VGND VPWR VPWR C_out\[186\] sky130_fd_sc_hd__dfrtp_1
XFILLER_120_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26426_ clknet_leaf_8_clk _00233_ net134 VGND VGND VPWR VPWR A_in\[94\] sky130_fd_sc_hd__dfrtp_1
X_14440_ _11619_ _11621_ VGND VGND VPWR VPWR _11622_ sky130_fd_sc_hd__nand2_2
X_23638_ _11269_ systolic_inst.B_outs\[0\]\[7\] _10120_ VGND VGND VPWR VPWR _10258_
+ sky130_fd_sc_hd__and3_1
XFILLER_126_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29145_ clknet_leaf_165_clk _02943_ net150 VGND VGND VPWR VPWR C_out\[117\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26357_ clknet_leaf_65_clk _00164_ net134 VGND VGND VPWR VPWR A_in\[25\] sky130_fd_sc_hd__dfrtp_1
X_14371_ _11518_ _11553_ VGND VGND VPWR VPWR _11555_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_189_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23569_ _10145_ _10190_ VGND VGND VPWR VPWR _10191_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16110_ _13070_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13322_ A_in\[31\] deser_A.word_buffer\[31\] net92 VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__mux2_1
X_25308_ net111 ser_C.shift_reg\[482\] VGND VGND VPWR VPWR _11124_ sky130_fd_sc_hd__and2_1
X_29076_ clknet_leaf_112_clk _02874_ net150 VGND VGND VPWR VPWR C_out\[48\] sky130_fd_sc_hd__dfrtp_1
XFILLER_128_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17090_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[18\]
+ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__or2_1
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26288_ clknet_leaf_27_A_in_serial_clk _00096_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_196_1226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_185_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28027_ clknet_leaf_161_clk _01825_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_16041_ systolic_inst.A_outs\[12\]\[2\] systolic_inst.B_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\]
+ systolic_inst.A_outs\[12\]\[1\] VGND VGND VPWR VPWR _13038_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_242_Left_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25239_ ser_C.parallel_data\[446\] net102 net74 ser_C.shift_reg\[446\] _11089_ VGND
+ VGND VPWR VPWR _02696_ sky130_fd_sc_hd__a221o_1
X_13253_ deser_A.word_buffer\[91\] deser_A.serial_word\[91\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13184_ deser_A.word_buffer\[22\] deser_A.serial_word\[22\] net128 VGND VGND VPWR
+ VPWR _00032_ sky130_fd_sc_hd__mux2_1
XFILLER_123_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19800_ _06792_ _06800_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_144_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17992_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[8\] VGND
+ VGND VPWR VPWR _05185_ sky130_fd_sc_hd__and2_1
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19731_ _06689_ _06691_ _06733_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__a21oi_1
X_16943_ _04169_ _04256_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__nand2_1
X_28929_ clknet_leaf_266_clk _02727_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[477\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19662_ _06663_ _06666_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16874_ _04190_ _04191_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__nor2_1
XFILLER_77_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15825_ _12862_ _12863_ VGND VGND VPWR VPWR _12864_ sky130_fd_sc_hd__xnor2_1
X_18613_ systolic_inst.A_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[6\]
+ systolic_inst.B_outs\[8\]\[7\] VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__and4b_1
X_19593_ _06618_ _06621_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__xor2_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15756_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[13\]\[0\]
+ _12803_ _12804_ VGND VGND VPWR VPWR _12805_ sky130_fd_sc_hd__and4_1
X_18544_ _05670_ _05673_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _11850_ _11852_ _11858_ VGND VGND VPWR VPWR _11859_ sky130_fd_sc_hd__a21o_1
X_18475_ systolic_inst.A_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[2\] systolic_inst.B_outs\[8\]\[3\]
+ systolic_inst.B_outs\[8\]\[4\] VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_174_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ _12738_ _12740_ VGND VGND VPWR VPWR _12741_ sky130_fd_sc_hd__nand2_1
XFILLER_209_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17426_ systolic_inst.A_outs\[10\]\[4\] systolic_inst.B_outs\[10\]\[6\] _11275_ systolic_inst.A_outs\[10\]\[3\]
+ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_99_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14638_ _11787_ _11794_ _11795_ VGND VGND VPWR VPWR _11800_ sky130_fd_sc_hd__o21ba_1
XFILLER_61_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17357_ systolic_inst.A_outs\[10\]\[2\] systolic_inst.B_outs\[10\]\[6\] _11275_ systolic_inst.A_outs\[10\]\[1\]
+ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_202_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14569_ _11734_ _11735_ _11733_ VGND VGND VPWR VPWR _11741_ sky130_fd_sc_hd__a21bo_1
XFILLER_147_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16308_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[12\] _03688_ net115
+ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__mux2_1
XFILLER_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload301 clknet_leaf_182_clk VGND VGND VPWR VPWR clkload301/Y sky130_fd_sc_hd__inv_8
X_17288_ _04540_ _04541_ _04545_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__a21o_1
Xclkload312 clknet_leaf_152_clk VGND VGND VPWR VPWR clkload312/Y sky130_fd_sc_hd__inv_6
XFILLER_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload20 clknet_5_24__leaf_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__inv_8
XFILLER_146_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload323 clknet_leaf_158_clk VGND VGND VPWR VPWR clkload323/Y sky130_fd_sc_hd__inv_6
X_19027_ net119 systolic_inst.B_outs\[7\]\[0\] systolic_inst.A_outs\[7\]\[0\] VGND
+ VGND VPWR VPWR _06100_ sky130_fd_sc_hd__and3_1
Xclkload334 clknet_leaf_162_clk VGND VGND VPWR VPWR clkload334/Y sky130_fd_sc_hd__clkinvlp_4
X_16239_ _03551_ _03585_ _03582_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__a21oi_1
Xclkload31 clknet_leaf_336_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__inv_8
XPHY_EDGE_ROW_224_Right_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload42 clknet_leaf_346_clk VGND VGND VPWR VPWR clkload42/X sky130_fd_sc_hd__clkbuf_8
Xclkload345 clknet_leaf_30_A_in_serial_clk VGND VGND VPWR VPWR clkload345/X sky130_fd_sc_hd__clkbuf_8
Xclkload356 clknet_leaf_7_A_in_serial_clk VGND VGND VPWR VPWR clkload356/Y sky130_fd_sc_hd__clkinv_4
Xclkload53 clknet_leaf_313_clk VGND VGND VPWR VPWR clkload53/Y sky130_fd_sc_hd__inv_8
Xclkload367 clknet_2_2__leaf_B_in_serial_clk VGND VGND VPWR VPWR clkload367/Y sky130_fd_sc_hd__inv_8
XFILLER_155_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload64 clknet_leaf_7_clk VGND VGND VPWR VPWR clkload64/Y sky130_fd_sc_hd__clkinv_8
XFILLER_103_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload378 clknet_leaf_33_B_in_serial_clk VGND VGND VPWR VPWR clkload378/Y sky130_fd_sc_hd__inv_6
XFILLER_86_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload75 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload75/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_90_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload389 clknet_leaf_9_B_in_serial_clk VGND VGND VPWR VPWR clkload389/Y sky130_fd_sc_hd__bufinv_16
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload86 clknet_leaf_303_clk VGND VGND VPWR VPWR clkload86/Y sky130_fd_sc_hd__inv_8
XFILLER_173_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload97 clknet_leaf_218_clk VGND VGND VPWR VPWR clkload97/Y sky130_fd_sc_hd__clkinv_2
XFILLER_216_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19929_ systolic_inst.A_outs\[6\]\[5\] systolic_inst.B_outs\[6\]\[6\] systolic_inst.A_outs\[6\]\[6\]
+ systolic_inst.B_outs\[6\]\[7\] VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__and4b_1
XFILLER_64_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22940_ _09580_ _09617_ _09616_ VGND VGND VPWR VPWR _09619_ sky130_fd_sc_hd__a21o_1
XFILLER_60_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22871_ net122 _09549_ _09550_ _09551_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__a31o_1
XFILLER_23_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24610_ net110 ser_C.shift_reg\[133\] VGND VGND VPWR VPWR _10775_ sky130_fd_sc_hd__and2_1
X_21822_ _08556_ _08595_ _08594_ VGND VGND VPWR VPWR _08626_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_84_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25590_ systolic_inst.acc_wires\[2\]\[2\] C_out\[66\] net34 VGND VGND VPWR VPWR _02892_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_233_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24541_ C_out\[97\] net99 net79 ser_C.shift_reg\[97\] _10740_ VGND VGND VPWR VPWR
+ _02347_ sky130_fd_sc_hd__a221o_1
XFILLER_197_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_233_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21753_ systolic_inst.A_outs\[3\]\[5\] systolic_inst.B_outs\[3\]\[6\] _11274_ systolic_inst.A_outs\[3\]\[4\]
+ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_233_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20704_ net109 systolic_inst.acc_wires\[5\]\[12\] net64 _07620_ VGND VGND VPWR VPWR
+ _01630_ sky130_fd_sc_hd__a22o_1
XFILLER_24_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27260_ clknet_leaf_270_clk _01058_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_43_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24472_ net114 ser_C.shift_reg\[64\] VGND VGND VPWR VPWR _10706_ sky130_fd_sc_hd__and2_1
XFILLER_211_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21684_ systolic_inst.A_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[6\] _11274_ systolic_inst.A_outs\[3\]\[2\]
+ VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_43_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26211_ clknet_leaf_13_A_in_serial_clk _00019_ net144 VGND VGND VPWR VPWR deser_A.word_buffer\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23423_ _10002_ _10007_ _10005_ VGND VGND VPWR VPWR _10049_ sky130_fd_sc_hd__a21bo_1
XFILLER_138_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20635_ net63 _07559_ _07561_ systolic_inst.acc_wires\[5\]\[2\] net107 VGND VGND
+ VPWR VPWR _01620_ sky130_fd_sc_hd__a32o_1
XFILLER_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27191_ clknet_leaf_247_clk _00989_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload3 clknet_5_3__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_6
Xwire118 net120 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_12
XFILLER_221_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26142_ deser_B.serial_word\[97\] deser_B.shift_reg\[97\] _00001_ VGND VGND VPWR
+ VPWR _03444_ sky130_fd_sc_hd__mux2_1
XFILLER_177_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23354_ _09970_ _09981_ VGND VGND VPWR VPWR _09982_ sky130_fd_sc_hd__xor2_1
X_20566_ _07469_ _07496_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22305_ _09010_ _09012_ _09046_ VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26073_ deser_B.serial_word\[28\] deser_B.shift_reg\[28\] net56 VGND VGND VPWR VPWR
+ _03375_ sky130_fd_sc_hd__mux2_1
XFILLER_153_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23285_ net121 systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[0\] VGND
+ VGND VPWR VPWR _09918_ sky130_fd_sc_hd__and3_1
X_20497_ _07322_ _07429_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__and2_1
XFILLER_180_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25024_ net112 ser_C.shift_reg\[340\] VGND VGND VPWR VPWR _10982_ sky130_fd_sc_hd__and2_1
XFILLER_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22236_ _08918_ _08953_ _08952_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_180_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22167_ net109 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[5\] _08913_
+ _08914_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_7_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21118_ _07953_ _07954_ _07956_ _07958_ _07917_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__a32o_1
X_22098_ net122 _08849_ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__nand2_1
X_26975_ clknet_leaf_28_A_in_serial_clk _00773_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21049_ _07877_ _07919_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__or2_1
X_25926_ systolic_inst.acc_wires\[12\]\[18\] C_out\[402\] net17 VGND VGND VPWR VPWR
+ _03228_ sky130_fd_sc_hd__mux2_1
X_13940_ deser_A.serial_word\[101\] deser_A.shift_reg\[101\] net57 VGND VGND VPWR
+ VPWR _00766_ sky130_fd_sc_hd__mux2_1
X_28714_ clknet_leaf_325_clk _02512_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[262\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29694_ clknet_leaf_9_clk _03489_ VGND VGND VPWR VPWR systolic_inst.A_shift\[30\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28645_ clknet_leaf_208_clk _02443_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13871_ deser_A.serial_word\[32\] deser_A.shift_reg\[32\] net58 VGND VGND VPWR VPWR
+ _00697_ sky130_fd_sc_hd__mux2_1
XFILLER_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25857_ systolic_inst.acc_wires\[10\]\[13\] C_out\[333\] net12 VGND VGND VPWR VPWR
+ _03159_ sky130_fd_sc_hd__mux2_1
X_15610_ _12615_ _12632_ _12631_ VGND VGND VPWR VPWR _12666_ sky130_fd_sc_hd__o21ba_1
XFILLER_75_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xload_slew59 _00008_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_16
X_24808_ net113 ser_C.shift_reg\[232\] VGND VGND VPWR VPWR _10874_ sky130_fd_sc_hd__and2_1
XFILLER_74_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28576_ clknet_leaf_172_clk _02374_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_16590_ systolic_inst.B_outs\[10\]\[7\] systolic_inst.B_outs\[6\]\[7\] net120 VGND
+ VGND VPWR VPWR _01217_ sky130_fd_sc_hd__mux2_1
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25788_ systolic_inst.acc_wires\[8\]\[8\] C_out\[264\] net22 VGND VGND VPWR VPWR
+ _03090_ sky130_fd_sc_hd__mux2_1
X_15541_ _12581_ _12598_ VGND VGND VPWR VPWR _12599_ sky130_fd_sc_hd__xor2_1
X_27527_ clknet_leaf_236_clk _01325_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_231_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24739_ C_out\[196\] net97 net77 ser_C.shift_reg\[196\] _10839_ VGND VGND VPWR VPWR
+ _02446_ sky130_fd_sc_hd__a221o_1
XFILLER_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18260_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[9\]\[11\]
+ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__or2_1
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27458_ clknet_leaf_237_clk _01256_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_15472_ _12529_ _12530_ _12507_ VGND VGND VPWR VPWR _12532_ sky130_fd_sc_hd__o21a_1
XFILLER_43_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17211_ systolic_inst.A_outs\[10\]\[1\] systolic_inst.B_outs\[10\]\[2\] systolic_inst.B_outs\[10\]\[3\]
+ systolic_inst.A_outs\[10\]\[0\] VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__a22oi_2
X_14423_ _11604_ _11605_ VGND VGND VPWR VPWR _11606_ sky130_fd_sc_hd__nand2b_1
X_26409_ clknet_leaf_4_clk _00216_ net131 VGND VGND VPWR VPWR A_in\[77\] sky130_fd_sc_hd__dfrtp_1
X_18191_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[9\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__a21o_1
X_27389_ clknet_leaf_337_clk _01187_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29128_ clknet_leaf_171_clk _02926_ net148 VGND VGND VPWR VPWR C_out\[100\] sky130_fd_sc_hd__dfrtp_1
X_17142_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[26\]
+ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__or2_1
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14354_ _11537_ _11538_ VGND VGND VPWR VPWR _11539_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13305_ A_in\[14\] deser_A.word_buffer\[14\] net93 VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__mux2_1
X_29059_ clknet_leaf_107_clk _02857_ net151 VGND VGND VPWR VPWR C_out\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17073_ _04369_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__or2_1
XFILLER_183_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14285_ _11435_ _11468_ _11434_ VGND VGND VPWR VPWR _11472_ sky130_fd_sc_hd__a21boi_1
XFILLER_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16024_ _13019_ _13021_ _13002_ VGND VGND VPWR VPWR _13022_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13236_ deser_A.word_buffer\[74\] deser_A.serial_word\[74\] net127 VGND VGND VPWR
+ VPWR _00084_ sky130_fd_sc_hd__mux2_1
XFILLER_152_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13167_ deser_A.word_buffer\[5\] deser_A.serial_word\[5\] net127 VGND VGND VPWR VPWR
+ _00015_ sky130_fd_sc_hd__mux2_1
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17975_ _05159_ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_163_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19714_ _06687_ _06716_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__and2_1
XFILLER_133_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16926_ _04200_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19645_ systolic_inst.A_outs\[6\]\[0\] systolic_inst.A_outs\[6\]\[1\] systolic_inst.B_outs\[6\]\[2\]
+ systolic_inst.B_outs\[6\]\[3\] VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__and4_1
X_16857_ _04135_ _04137_ _04136_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__o21ba_1
XFILLER_93_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15808_ _12844_ _12847_ VGND VGND VPWR VPWR _12849_ sky130_fd_sc_hd__nand2_1
X_19576_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[26\]
+ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__or2_1
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16788_ _04107_ _04106_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__nand2b_1
XFILLER_34_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15739_ _12744_ _12768_ _12790_ VGND VGND VPWR VPWR _12791_ sky130_fd_sc_hd__a21o_1
X_18527_ _05633_ _05635_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__nand2_1
XFILLER_94_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18458_ _05572_ _05589_ _05590_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__nor3_1
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17409_ _04627_ _04629_ _04664_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__a21o_1
X_18389_ _05542_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20420_ _07354_ _07355_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_116_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1058 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20351_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[5\] systolic_inst.A_outs\[5\]\[6\]
+ systolic_inst.B_outs\[5\]\[1\] VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload120 clknet_leaf_293_clk VGND VGND VPWR VPWR clkload120/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_295_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_295_clk
+ sky130_fd_sc_hd__clkbuf_8
Xclkload131 clknet_leaf_266_clk VGND VGND VPWR VPWR clkload131/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload142 clknet_leaf_257_clk VGND VGND VPWR VPWR clkload142/Y sky130_fd_sc_hd__inv_6
Xclkload153 clknet_leaf_201_clk VGND VGND VPWR VPWR clkload153/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_77_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23070_ net122 _09741_ _09742_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__a21oi_1
Xclkload164 clknet_leaf_225_clk VGND VGND VPWR VPWR clkload164/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_77_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20282_ _07219_ _07221_ _07213_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__a21oi_1
Xclkload175 clknet_leaf_196_clk VGND VGND VPWR VPWR clkload175/Y sky130_fd_sc_hd__clkinv_2
Xclkload186 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload186/X sky130_fd_sc_hd__clkbuf_8
XFILLER_192_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22021_ net106 systolic_inst.acc_wires\[3\]\[22\] net65 _08799_ VGND VGND VPWR VPWR
+ _01768_ sky130_fd_sc_hd__a22o_1
Xclkload197 clknet_leaf_61_clk VGND VGND VPWR VPWR clkload197/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_129_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_222_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26760_ clknet_leaf_76_clk _00562_ net144 VGND VGND VPWR VPWR B_in\[32\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23972_ _10511_ systolic_inst.B_shift\[9\]\[5\] _11332_ VGND VGND VPWR VPWR _02007_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25711_ systolic_inst.acc_wires\[5\]\[27\] C_out\[187\] net48 VGND VGND VPWR VPWR
+ _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_57_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22923_ _09592_ _09600_ VGND VGND VPWR VPWR _09602_ sky130_fd_sc_hd__or2_1
XFILLER_151_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_235_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26691_ clknet_leaf_33_B_in_serial_clk _00494_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_235_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_235_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28430_ clknet_leaf_25_clk _02228_ VGND VGND VPWR VPWR systolic_inst.A_shift\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25642_ systolic_inst.acc_wires\[3\]\[22\] C_out\[118\] net50 VGND VGND VPWR VPWR
+ _02944_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22854_ _09525_ _09534_ VGND VGND VPWR VPWR _09535_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21805_ _08609_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__inv_2
X_28361_ clknet_leaf_75_clk _02159_ VGND VGND VPWR VPWR systolic_inst.B_shift\[22\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25573_ systolic_inst.acc_wires\[1\]\[17\] C_out\[49\] net34 VGND VGND VPWR VPWR
+ _02875_ sky130_fd_sc_hd__mux2_1
XFILLER_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22785_ _09456_ _09466_ _09467_ VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__nand3_1
X_27312_ clknet_leaf_293_clk _01110_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24524_ net114 ser_C.shift_reg\[90\] VGND VGND VPWR VPWR _10732_ sky130_fd_sc_hd__and2_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28292_ clknet_leaf_99_clk _02090_ VGND VGND VPWR VPWR systolic_inst.B_shift\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_21736_ _08480_ _08505_ _08504_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__a21boi_1
XFILLER_223_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27243_ clknet_leaf_279_clk _01041_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24455_ C_out\[54\] net100 net82 ser_C.shift_reg\[54\] _10697_ VGND VGND VPWR VPWR
+ _02304_ sky130_fd_sc_hd__a221o_1
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21667_ _08435_ _08437_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__and2_1
XFILLER_177_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_A_in_serial_clk clknet_2_2__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_4_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_23406_ _09991_ _10031_ VGND VGND VPWR VPWR _10032_ sky130_fd_sc_hd__nand2_1
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20618_ systolic_inst.ce_local _07540_ _07547_ _07541_ VGND VGND VPWR VPWR _01617_
+ sky130_fd_sc_hd__a31o_1
X_27174_ clknet_leaf_248_clk _00972_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24386_ net7 ser_C.shift_reg\[21\] VGND VGND VPWR VPWR _10663_ sky130_fd_sc_hd__and2_1
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21598_ _11274_ _08407_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26125_ deser_B.serial_word\[80\] deser_B.shift_reg\[80\] net55 VGND VGND VPWR VPWR
+ _03427_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_286_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_286_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_193_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23337_ _09939_ _09941_ _09959_ _09960_ VGND VGND VPWR VPWR _09965_ sky130_fd_sc_hd__a211o_1
X_20549_ _07479_ _07480_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14070_ deser_B.shift_reg\[104\] deser_B.shift_reg\[105\] net126 VGND VGND VPWR VPWR
+ _00896_ sky130_fd_sc_hd__mux2_1
X_26056_ deser_B.serial_word\[11\] deser_B.shift_reg\[11\] net55 VGND VGND VPWR VPWR
+ _03358_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_32_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_32_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_23268_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[30\]
+ VGND VGND VPWR VPWR _09911_ sky130_fd_sc_hd__or2_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25007_ C_out\[330\] net97 net80 ser_C.shift_reg\[330\] _10973_ VGND VGND VPWR VPWR
+ _02580_ sky130_fd_sc_hd__a221o_1
XFILLER_238_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22219_ _08929_ _08964_ VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__xnor2_1
X_23199_ net109 systolic_inst.acc_wires\[1\]\[19\] net65 _09852_ VGND VGND VPWR VPWR
+ _01893_ sky130_fd_sc_hd__a22o_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14972_ _12050_ _12051_ _12053_ VGND VGND VPWR VPWR _12093_ sky130_fd_sc_hd__o21a_1
XFILLER_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17760_ _04974_ _04978_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__nor2_1
X_26958_ clknet_leaf_2_A_in_serial_clk _00756_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13923_ deser_A.serial_word\[84\] deser_A.shift_reg\[84\] net57 VGND VGND VPWR VPWR
+ _00749_ sky130_fd_sc_hd__mux2_1
X_16711_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[7\] VGND VGND
+ VPWR VPWR _04033_ sky130_fd_sc_hd__and2b_1
X_17691_ net105 systolic_inst.acc_wires\[10\]\[16\] _04921_ _04923_ VGND VGND VPWR
+ VPWR _01314_ sky130_fd_sc_hd__a22o_1
X_25909_ systolic_inst.acc_wires\[12\]\[1\] C_out\[385\] net20 VGND VGND VPWR VPWR
+ _03211_ sky130_fd_sc_hd__mux2_1
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29677_ clknet_leaf_32_B_in_serial_clk _03472_ net134 VGND VGND VPWR VPWR deser_B.serial_word\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26889_ clknet_leaf_6_A_in_serial_clk _00687_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_210_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_210_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_35_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19430_ _06473_ _06477_ _06480_ _06481_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__o211a_1
X_16642_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[4\]
+ systolic_inst.A_outs\[11\]\[5\] VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__and4_1
X_28628_ clknet_leaf_206_clk _02426_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[176\]
+ sky130_fd_sc_hd__dfrtp_1
X_13854_ deser_A.serial_word\[15\] deser_A.shift_reg\[15\] net58 VGND VGND VPWR VPWR
+ _00680_ sky130_fd_sc_hd__mux2_1
XFILLER_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19361_ _06420_ _06419_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__and2b_1
X_16573_ _03917_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__xnor2_1
X_28559_ clknet_leaf_169_clk _02357_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_13785_ B_in\[92\] deser_B.word_buffer\[92\] net89 VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__mux2_1
XFILLER_188_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18312_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[18\]
+ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__or2_1
X_15524_ systolic_inst.B_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[4\]
+ systolic_inst.A_outs\[13\]\[5\] VGND VGND VPWR VPWR _12582_ sky130_fd_sc_hd__and4_1
XFILLER_206_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19292_ _06313_ _06315_ _06314_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__o21ba_1
XFILLER_76_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18243_ _05418_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__nand2_1
XFILLER_203_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15455_ systolic_inst.A_outs\[13\]\[2\] systolic_inst.B_outs\[13\]\[3\] systolic_inst.A_outs\[13\]\[3\]
+ systolic_inst.B_outs\[13\]\[4\] VGND VGND VPWR VPWR _12515_ sky130_fd_sc_hd__nand4_2
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14406_ _11518_ _11587_ VGND VGND VPWR VPWR _11589_ sky130_fd_sc_hd__and2_1
XFILLER_15_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18174_ _05359_ _05360_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_152_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15386_ net116 _12448_ _12449_ _12442_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__a31o_1
XFILLER_89_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17125_ _04407_ _04411_ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_277_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_277_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_237_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14337_ _11478_ _11520_ VGND VGND VPWR VPWR _11522_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_169_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17056_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[11\]\[12\]
+ _04353_ _04355_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__a211o_1
X_14268_ _11416_ _11453_ VGND VGND VPWR VPWR _11455_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_111_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16007_ systolic_inst.A_outs\[12\]\[0\] systolic_inst.A_outs\[12\]\[1\] systolic_inst.B_outs\[12\]\[3\]
+ systolic_inst.B_outs\[12\]\[4\] VGND VGND VPWR VPWR _13005_ sky130_fd_sc_hd__nand4_1
X_13219_ deser_A.word_buffer\[57\] deser_A.serial_word\[57\] net128 VGND VGND VPWR
+ VPWR _00067_ sky130_fd_sc_hd__mux2_1
XFILLER_174_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14199_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[3\]
+ systolic_inst.B_outs\[15\]\[4\] VGND VGND VPWR VPWR _11388_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_72_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17958_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] _05150_ VGND
+ VGND VPWR VPWR _05151_ sky130_fd_sc_hd__a21o_1
XFILLER_97_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16909_ _04223_ _04225_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_109_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17889_ _05053_ _05083_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__and2_1
XFILLER_81_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_201_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_201_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19628_ net119 systolic_inst.B_outs\[6\]\[0\] systolic_inst.A_outs\[6\]\[0\] VGND
+ VGND VPWR VPWR _06637_ sky130_fd_sc_hd__and3_1
XFILLER_54_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19559_ _06585_ _06589_ _06592_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_230_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22570_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[15\]
+ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__and2_1
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21521_ _08314_ _08333_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__nor2_1
XFILLER_142_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24240_ _10605_ systolic_inst.A_shift\[18\]\[3\] net70 VGND VGND VPWR VPWR _02181_
+ sky130_fd_sc_hd__mux2_1
X_21452_ systolic_inst.acc_wires\[4\]\[28\] systolic_inst.acc_wires\[4\]\[29\] systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__o21ai_1
XFILLER_119_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_268_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_268_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_228_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20403_ systolic_inst.B_outs\[5\]\[7\] _07337_ _07338_ VGND VGND VPWR VPWR _07340_
+ sky130_fd_sc_hd__and3_1
XFILLER_181_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21383_ _08222_ _08226_ _08228_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_21_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24171_ systolic_inst.A_shift\[26\]\[2\] net70 _10505_ systolic_inst.A_shift\[27\]\[2\]
+ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_165_Left_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23122_ _09784_ _09785_ net64 VGND VGND VPWR VPWR _09787_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_224_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20334_ _07241_ _07271_ _07272_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__nand3_1
XFILLER_107_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23053_ _09654_ _09727_ VGND VGND VPWR VPWR _09728_ sky130_fd_sc_hd__xnor2_1
X_27930_ clknet_leaf_134_clk _01728_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_20265_ _07192_ _07194_ _07205_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__a21oi_1
XFILLER_157_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22004_ _08765_ _08769_ _08774_ _08779_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__or4_1
XFILLER_192_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27861_ clknet_leaf_141_clk _01659_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20196_ _07160_ _07161_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29600_ clknet_leaf_18_B_in_serial_clk _03395_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_26812_ clknet_leaf_75_clk _00614_ net144 VGND VGND VPWR VPWR B_in\[84\] sky130_fd_sc_hd__dfrtp_1
XFILLER_131_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27792_ clknet_leaf_41_clk _01590_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26743_ clknet_leaf_97_clk _00545_ net153 VGND VGND VPWR VPWR B_in\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29531_ clknet_leaf_259_clk _03329_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23955_ systolic_inst.B_shift\[11\]\[2\] net70 net83 systolic_inst.B_shift\[15\]\[2\]
+ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_174_Left_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22906_ _09557_ _09558_ _09559_ VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__o21ba_1
X_29462_ clknet_leaf_331_clk _03260_ net136 VGND VGND VPWR VPWR C_out\[434\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26674_ clknet_leaf_13_B_in_serial_clk _00477_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_23886_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[30\]
+ VGND VGND VPWR VPWR _10473_ sky130_fd_sc_hd__nand2_1
XFILLER_45_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_B_in_serial_clk clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_11_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_25625_ systolic_inst.acc_wires\[3\]\[5\] C_out\[101\] net48 VGND VGND VPWR VPWR
+ _02927_ sky130_fd_sc_hd__mux2_1
X_28413_ clknet_leaf_60_clk _02211_ VGND VGND VPWR VPWR systolic_inst.B_shift\[23\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_22837_ _09517_ _09514_ VGND VGND VPWR VPWR _09518_ sky130_fd_sc_hd__and2b_1
X_29393_ clknet_leaf_235_clk _03191_ net145 VGND VGND VPWR VPWR C_out\[365\] sky130_fd_sc_hd__dfrtp_1
XFILLER_147_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28344_ clknet_leaf_343_clk _02142_ VGND VGND VPWR VPWR systolic_inst.A_shift\[25\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_25556_ systolic_inst.acc_wires\[1\]\[0\] C_out\[32\] net54 VGND VGND VPWR VPWR _02858_
+ sky130_fd_sc_hd__mux2_1
X_13570_ deser_B.word_buffer\[6\] deser_B.serial_word\[6\] net124 VGND VGND VPWR VPWR
+ _00407_ sky130_fd_sc_hd__mux2_1
XFILLER_241_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22768_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[5\]
+ systolic_inst.A_outs\[1\]\[6\] VGND VGND VPWR VPWR _09451_ sky130_fd_sc_hd__and4_1
XFILLER_201_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24507_ C_out\[80\] net100 net80 ser_C.shift_reg\[80\] _10723_ VGND VGND VPWR VPWR
+ _02330_ sky130_fd_sc_hd__a221o_1
XFILLER_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_213_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21719_ _08522_ _08525_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__xnor2_1
X_28275_ clknet_leaf_130_clk _02073_ VGND VGND VPWR VPWR systolic_inst.B_shift\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25487_ systolic_inst.cycle_cnt\[17\] systolic_inst.cycle_cnt\[16\] _11306_ _11215_
+ systolic_inst.cycle_cnt\[18\] VGND VGND VPWR VPWR _11222_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_213_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22699_ _09383_ _09384_ _09379_ VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__or3b_1
XFILLER_197_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15240_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[14\]\[14\]
+ VGND VGND VPWR VPWR _12340_ sky130_fd_sc_hd__or2_1
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27226_ clknet_leaf_326_clk _01024_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_24438_ net114 ser_C.shift_reg\[47\] VGND VGND VPWR VPWR _10689_ sky130_fd_sc_hd__and2_1
XFILLER_200_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_183_Left_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_259_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_259_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15171_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[14\]\[4\]
+ VGND VGND VPWR VPWR _12281_ sky130_fd_sc_hd__nand2_1
X_27157_ clknet_leaf_294_clk _00955_ net138 VGND VGND VPWR VPWR systolic_inst.B_outs\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_24369_ C_out\[11\] net104 _10643_ ser_C.shift_reg\[11\] _10654_ VGND VGND VPWR VPWR
+ _02261_ sky130_fd_sc_hd__a221o_1
XFILLER_181_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26108_ deser_B.serial_word\[63\] deser_B.shift_reg\[63\] net56 VGND VGND VPWR VPWR
+ _03410_ sky130_fd_sc_hd__mux2_1
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14122_ systolic_inst.A_shift\[21\]\[6\] net71 _11333_ A_in\[94\] VGND VGND VPWR
+ VPWR _00944_ sky130_fd_sc_hd__a22o_1
XFILLER_4_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27088_ clknet_leaf_0_B_in_serial_clk _00886_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_193_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14053_ deser_B.shift_reg\[87\] deser_B.shift_reg\[88\] net125 VGND VGND VPWR VPWR
+ _00879_ sky130_fd_sc_hd__mux2_1
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18930_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[19\]
+ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__xnor2_1
X_26039_ systolic_inst.B_outs\[15\]\[3\] systolic_inst.B_outs\[11\]\[3\] net118 VGND
+ VGND VPWR VPWR _03341_ sky130_fd_sc_hd__mux2_1
XFILLER_234_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18861_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[8\]\[10\]
+ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_160_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17812_ _05003_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__xnor2_1
X_18792_ _05833_ _05834_ _05901_ _05899_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__a31o_1
XFILLER_239_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_192_Left_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14955_ systolic_inst.B_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[5\] systolic_inst.A_outs\[14\]\[6\]
+ systolic_inst.B_outs\[14\]\[3\] VGND VGND VPWR VPWR _12076_ sky130_fd_sc_hd__a22oi_1
X_17743_ _04961_ _04963_ _04966_ net60 VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__a31o_1
XFILLER_212_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13906_ deser_A.serial_word\[67\] deser_A.shift_reg\[67\] net57 VGND VGND VPWR VPWR
+ _00732_ sky130_fd_sc_hd__mux2_1
XFILLER_208_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14886_ _11975_ _12007_ VGND VGND VPWR VPWR _12009_ sky130_fd_sc_hd__xnor2_1
X_17674_ _04901_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__nand2_1
XFILLER_208_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19413_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[7\]\[2\]
+ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__nand2_1
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13837_ deser_B.bit_idx\[5\] _11327_ deser_B.bit_idx\[6\] VGND VGND VPWR VPWR _11329_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_158_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16625_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[3\]
+ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__and3_1
XFILLER_63_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap91 net92 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_12
XFILLER_189_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19344_ systolic_inst.B_outs\[7\]\[6\] systolic_inst.A_outs\[7\]\[7\] VGND VGND VPWR
+ VPWR _06404_ sky130_fd_sc_hd__nand2_1
X_16556_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[28\]
+ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__xnor2_1
X_13768_ B_in\[75\] deser_B.word_buffer\[75\] net90 VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__mux2_1
XFILLER_188_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15507_ _12563_ _12564_ VGND VGND VPWR VPWR _12566_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19275_ _06299_ _06336_ _06337_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__and3_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_16487_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[17\]
+ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_61_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13699_ B_in\[6\] deser_B.word_buffer\[6\] net84 VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__mux2_1
XFILLER_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15438_ _12475_ _12498_ VGND VGND VPWR VPWR _12499_ sky130_fd_sc_hd__nand2_1
X_18226_ _05396_ _05400_ _05403_ _05404_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__o211a_1
XFILLER_176_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15369_ systolic_inst.B_outs\[12\]\[5\] systolic_inst.B_outs\[8\]\[5\] net115 VGND
+ VGND VPWR VPWR _01087_ sky130_fd_sc_hd__mux2_1
X_18157_ _05313_ _05317_ _05343_ net116 VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__o31a_1
XFILLER_144_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17108_ _04398_ _04399_ _04396_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__o21ai_2
X_18088_ _05277_ _05276_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__and2b_1
XFILLER_172_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_886 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17039_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[11\]\[11\]
+ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__nor2_1
XFILLER_116_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20050_ net66 _07035_ _07037_ systolic_inst.acc_wires\[6\]\[5\] net106 VGND VGND
+ VPWR VPWR _01559_ sky130_fd_sc_hd__a32o_1
XFILLER_139_1090 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23740_ _10346_ _10347_ _10348_ VGND VGND VPWR VPWR _10350_ sky130_fd_sc_hd__nand3_1
XFILLER_2_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20952_ _07788_ _07789_ _07790_ _07793_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__a31o_1
XFILLER_242_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_217_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23671_ _10261_ _10288_ _10289_ VGND VGND VPWR VPWR _10290_ sky130_fd_sc_hd__a21oi_2
XFILLER_14_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20883_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[4\] _07757_ _07759_
+ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__and4_1
XFILLER_35_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25410_ _11174_ systolic_inst.A_shift\[1\]\[4\] net70 VGND VGND VPWR VPWR _02782_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22622_ _09335_ _09334_ systolic_inst.acc_wires\[2\]\[23\] net109 VGND VGND VPWR
+ VPWR _01833_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_27_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26390_ clknet_leaf_17_clk _00197_ net132 VGND VGND VPWR VPWR A_in\[58\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25341_ ser_C.parallel_data\[497\] net97 net77 ser_C.shift_reg\[497\] _11140_ VGND
+ VGND VPWR VPWR _02747_ sky130_fd_sc_hd__a221o_1
XFILLER_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22553_ net109 systolic_inst.acc_wires\[2\]\[12\] net65 _09277_ VGND VGND VPWR VPWR
+ _01822_ sky130_fd_sc_hd__a22o_1
XFILLER_22_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28060_ clknet_leaf_101_clk _01858_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_21504_ _08316_ _08317_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__nand2_1
X_25272_ net111 ser_C.shift_reg\[464\] VGND VGND VPWR VPWR _11106_ sky130_fd_sc_hd__and2_1
XFILLER_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22484_ net65 _09216_ _09218_ systolic_inst.acc_wires\[2\]\[2\] net109 VGND VGND
+ VPWR VPWR _01812_ sky130_fd_sc_hd__a32o_1
X_27011_ clknet_leaf_21_B_in_serial_clk _00809_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_194_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24223_ systolic_inst.A_shift\[20\]\[3\] A_in\[75\] net59 VGND VGND VPWR VPWR _10597_
+ sky130_fd_sc_hd__mux2_1
X_21435_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[27\]
+ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__xnor2_1
XFILLER_213_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24154_ _10578_ systolic_inst.A_shift\[27\]\[0\] net70 VGND VGND VPWR VPWR _02122_
+ sky130_fd_sc_hd__mux2_1
X_21366_ _08211_ _08214_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23105_ net64 _09770_ _09772_ systolic_inst.acc_wires\[1\]\[5\] _11258_ VGND VGND
+ VPWR VPWR _01879_ sky130_fd_sc_hd__a32o_1
XFILLER_150_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20317_ systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[5\] systolic_inst.A_outs\[5\]\[6\]
+ systolic_inst.B_outs\[5\]\[0\] VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__a22oi_1
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24085_ systolic_inst.B_shift\[2\]\[4\] _11332_ net83 systolic_inst.B_shift\[6\]\[4\]
+ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__a22o_1
X_28962_ clknet_leaf_246_clk _02760_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[510\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21297_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[4\]\[7\]
+ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23036_ net109 systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[13\] VGND
+ VGND VPWR VPWR _09712_ sky130_fd_sc_hd__and2_1
X_27913_ clknet_leaf_135_clk _01711_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_20248_ _07189_ _07190_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__or2_1
X_28893_ clknet_leaf_286_clk _02691_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[441\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20179_ _07142_ _07144_ _07147_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__and3_1
X_27844_ clknet_leaf_181_clk _01642_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_191_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_202_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_202_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27775_ clknet_leaf_177_clk _01573_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_24987_ C_out\[320\] net102 net74 ser_C.shift_reg\[320\] _10963_ VGND VGND VPWR VPWR
+ _02570_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_198_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29514_ clknet_leaf_260_clk _03312_ net140 VGND VGND VPWR VPWR ser_C.parallel_data\[486\]
+ sky130_fd_sc_hd__dfrtp_1
X_14740_ systolic_inst.A_outs\[14\]\[0\] systolic_inst.A_outs\[13\]\[0\] net116 VGND
+ VGND VPWR VPWR _01010_ sky130_fd_sc_hd__mux2_1
X_23938_ systolic_inst.B_shift\[14\]\[1\] B_in\[17\] net59 VGND VGND VPWR VPWR _10498_
+ sky130_fd_sc_hd__mux2_1
X_26726_ clknet_leaf_3_B_in_serial_clk _00006_ net144 VGND VGND VPWR VPWR deser_B.receiving
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_85_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_194_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_194_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26657_ clknet_leaf_24_B_in_serial_clk _00460_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_14671_ _11827_ VGND VGND VPWR VPWR _11828_ sky130_fd_sc_hd__inv_2
XFILLER_45_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29445_ clknet_leaf_300_clk _03243_ net141 VGND VGND VPWR VPWR C_out\[417\] sky130_fd_sc_hd__dfrtp_1
X_23869_ _10457_ _10458_ VGND VGND VPWR VPWR _10459_ sky130_fd_sc_hd__xnor2_1
XFILLER_229_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16410_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[12\]\[7\]
+ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__nand2_1
XFILLER_232_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25608_ systolic_inst.acc_wires\[2\]\[20\] C_out\[84\] net52 VGND VGND VPWR VPWR
+ _02910_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13622_ deser_B.word_buffer\[58\] deser_B.serial_word\[58\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__mux2_1
XFILLER_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17390_ _04644_ _04645_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__nor2_1
X_26588_ clknet_leaf_0_A_in_serial_clk _00391_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_29376_ clknet_leaf_240_clk _03174_ net145 VGND VGND VPWR VPWR C_out\[348\] sky130_fd_sc_hd__dfrtp_1
X_16341_ _03694_ _03697_ _03719_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__a21oi_1
X_25539_ systolic_inst.acc_wires\[0\]\[15\] C_out\[15\] net54 VGND VGND VPWR VPWR
+ _02841_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28327_ clknet_leaf_343_clk _02125_ VGND VGND VPWR VPWR systolic_inst.A_shift\[27\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13553_ deser_A.shift_reg\[117\] deser_A.shift_reg\[118\] net130 VGND VGND VPWR VPWR
+ _00390_ sky130_fd_sc_hd__mux2_1
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19060_ _06125_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__xnor2_1
X_28258_ clknet_leaf_98_clk _02056_ VGND VGND VPWR VPWR systolic_inst.B_shift\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16272_ _03651_ _03652_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13484_ deser_A.shift_reg\[48\] deser_A.shift_reg\[49\] net130 VGND VGND VPWR VPWR
+ _00321_ sky130_fd_sc_hd__mux2_1
XFILLER_173_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15223_ net107 systolic_inst.acc_wires\[14\]\[11\] _11712_ _12325_ VGND VGND VPWR
+ VPWR _01053_ sky130_fd_sc_hd__a22o_1
X_27209_ clknet_leaf_256_clk _01007_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_18011_ _05200_ _05201_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28189_ clknet_leaf_125_clk _01987_ VGND VGND VPWR VPWR systolic_inst.B_shift\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15154_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[14\]\[0\]
+ _12263_ _12264_ VGND VGND VPWR VPWR _12267_ sky130_fd_sc_hd__a22o_1
XFILLER_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14105_ systolic_inst.A_shift\[12\]\[5\] net72 _11333_ A_in\[61\] VGND VGND VPWR
+ VPWR _00927_ sky130_fd_sc_hd__a22o_1
XFILLER_236_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19962_ _06957_ _06956_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__nand2b_1
X_15085_ _12134_ _12138_ _12168_ _12201_ _12166_ VGND VGND VPWR VPWR _12203_ sky130_fd_sc_hd__o311a_1
X_14036_ deser_B.shift_reg\[70\] deser_B.shift_reg\[71\] net126 VGND VGND VPWR VPWR
+ _00862_ sky130_fd_sc_hd__mux2_1
XFILLER_180_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18913_ _06014_ _06017_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19893_ _06783_ _06889_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__nand2_1
XFILLER_45_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_B_in_serial_clk clknet_2_2__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_6_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_110_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18844_ _05956_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__nand2_1
XFILLER_68_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18775_ _05896_ _05897_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__nand2_1
X_15987_ systolic_inst.A_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[2\] _12986_ VGND
+ VGND VPWR VPWR _12987_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17726_ _04944_ _04945_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__nor2_1
XFILLER_94_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14938_ _12019_ _12021_ VGND VGND VPWR VPWR _12060_ sky130_fd_sc_hd__and2_1
XFILLER_242_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17657_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[10\]\[12\]
+ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14869_ _11969_ _11971_ _11970_ VGND VGND VPWR VPWR _11992_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_63_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16608_ _03932_ _03933_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__nor2_1
X_17588_ _04832_ _04833_ _04834_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__a21o_1
XFILLER_91_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19327_ _06386_ _06387_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__nand2_1
XFILLER_204_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16539_ net108 systolic_inst.acc_wires\[12\]\[25\] net67 _03890_ VGND VGND VPWR VPWR
+ _01195_ sky130_fd_sc_hd__a22o_1
XFILLER_91_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19258_ _06312_ _06320_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__nand2_1
XFILLER_176_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18209_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[9\]\[3\]
+ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__nand2_1
X_19189_ _06253_ _06252_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__nand2b_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21220_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[13\] _08087_ net117
+ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21151_ _08020_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20102_ _07073_ _07074_ _07081_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__a21o_1
XFILLER_137_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21082_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[7\] _07924_ _07884_
+ systolic_inst.A_outs\[4\]\[4\] VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_242_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20033_ _07020_ _07021_ _07022_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__a21o_1
XFILLER_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24910_ net110 ser_C.shift_reg\[283\] VGND VGND VPWR VPWR _10925_ sky130_fd_sc_hd__and2_1
XFILLER_99_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25890_ systolic_inst.acc_wires\[11\]\[14\] C_out\[366\] net40 VGND VGND VPWR VPWR
+ _03192_ sky130_fd_sc_hd__mux2_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_219_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24841_ C_out\[247\] net98 net78 ser_C.shift_reg\[247\] _10890_ VGND VGND VPWR VPWR
+ _02497_ sky130_fd_sc_hd__a221o_1
XFILLER_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_219_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27560_ clknet_leaf_305_clk _01358_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24772_ net113 ser_C.shift_reg\[214\] VGND VGND VPWR VPWR _10856_ sky130_fd_sc_hd__and2_1
XFILLER_6_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21984_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[17\]
+ VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__xor2_2
XFILLER_2_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26511_ clknet_leaf_11_A_in_serial_clk _00314_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_199_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23723_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[0\]\[5\]
+ VGND VGND VPWR VPWR _10335_ sky130_fd_sc_hd__or2_1
XFILLER_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27491_ clknet_leaf_227_clk _01289_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_20935_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[4\] VGND VGND VPWR
+ VPWR _07810_ sky130_fd_sc_hd__nand2_1
XFILLER_57_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29230_ clknet_leaf_203_clk _03028_ net147 VGND VGND VPWR VPWR C_out\[202\] sky130_fd_sc_hd__dfrtp_1
XFILLER_148_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26442_ clknet_leaf_347_clk _00249_ net132 VGND VGND VPWR VPWR A_in\[110\] sky130_fd_sc_hd__dfrtp_1
XFILLER_187_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23654_ _10238_ _10241_ _10273_ VGND VGND VPWR VPWR _10274_ sky130_fd_sc_hd__a21oi_1
XFILLER_214_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20866_ _07731_ _07742_ _07743_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_238_Right_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22605_ net65 _09320_ _09321_ systolic_inst.acc_wires\[2\]\[20\] net109 VGND VGND
+ VPWR VPWR _01830_ sky130_fd_sc_hd__a32o_1
X_29161_ clknet_leaf_309_clk _02959_ net142 VGND VGND VPWR VPWR C_out\[133\] sky130_fd_sc_hd__dfrtp_1
X_26373_ clknet_leaf_24_clk _00180_ net143 VGND VGND VPWR VPWR A_in\[41\] sky130_fd_sc_hd__dfrtp_1
X_23585_ _10205_ _10206_ VGND VGND VPWR VPWR _10207_ sky130_fd_sc_hd__or2_1
XFILLER_35_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20797_ net106 systolic_inst.acc_wires\[5\]\[26\] net68 _07699_ VGND VGND VPWR VPWR
+ _01644_ sky130_fd_sc_hd__a22o_1
XFILLER_168_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28112_ clknet_leaf_47_clk _01910_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_46_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25324_ net112 ser_C.shift_reg\[490\] VGND VGND VPWR VPWR _11132_ sky130_fd_sc_hd__and2_1
X_29092_ clknet_leaf_155_clk _02890_ net150 VGND VGND VPWR VPWR C_out\[64\] sky130_fd_sc_hd__dfrtp_1
X_22536_ _09260_ _09262_ VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__xor2_1
XFILLER_22_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28043_ clknet_leaf_166_clk _01841_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25255_ ser_C.parallel_data\[454\] net102 net74 ser_C.shift_reg\[454\] _11097_ VGND
+ VGND VPWR VPWR _02704_ sky130_fd_sc_hd__a221o_1
XFILLER_202_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22467_ _09204_ _09203_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ net106 VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_167_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24206_ _10588_ systolic_inst.A_shift\[20\]\[2\] net71 VGND VGND VPWR VPWR _02164_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_187_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21418_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[24\]
+ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__nor2_1
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25186_ net111 ser_C.shift_reg\[421\] VGND VGND VPWR VPWR _11063_ sky130_fd_sc_hd__and2_1
XFILLER_204_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22398_ _09137_ _09138_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__nand2_1
XFILLER_159_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_208_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24137_ systolic_inst.A_shift\[29\]\[0\] A_in\[104\] net59 VGND VGND VPWR VPWR _10570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21349_ _08188_ _08193_ _08192_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__o21a_1
XFILLER_11_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24068_ _10551_ systolic_inst.B_shift\[15\]\[5\] net71 VGND VGND VPWR VPWR _02063_
+ sky130_fd_sc_hd__mux2_1
X_28945_ clknet_leaf_257_clk _02743_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[493\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_204_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23019_ _09627_ _09693_ VGND VGND VPWR VPWR _09695_ sky130_fd_sc_hd__or2_1
X_15910_ _12892_ _12893_ _12915_ _12935_ VGND VGND VPWR VPWR _12936_ sky130_fd_sc_hd__a211o_1
XFILLER_133_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28876_ clknet_leaf_285_clk _02674_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[424\]
+ sky130_fd_sc_hd__dfrtp_1
X_16890_ _04206_ _04205_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__nand2b_1
XFILLER_104_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27827_ clknet_leaf_140_clk _01625_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15841_ net61 _12877_ VGND VGND VPWR VPWR _12878_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18560_ _05688_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__xor2_1
XFILLER_224_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27758_ clknet_leaf_209_clk _01556_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_15772_ _12818_ VGND VGND VPWR VPWR _12819_ sky130_fd_sc_hd__inv_2
XFILLER_79_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17511_ _04761_ _04762_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__and2_1
X_26709_ clknet_leaf_10_B_in_serial_clk _00512_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_14723_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[29\]
+ VGND VGND VPWR VPWR _11872_ sky130_fd_sc_hd__xor2_1
XFILLER_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18491_ _05621_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__nand2_1
XFILLER_73_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27689_ clknet_leaf_191_clk _01487_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14654_ _11804_ _11806_ _11813_ VGND VGND VPWR VPWR _11814_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29428_ clknet_leaf_344_clk _03226_ net131 VGND VGND VPWR VPWR C_out\[400\] sky130_fd_sc_hd__dfrtp_1
X_17442_ _04640_ _04696_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__nand2_1
XFILLER_232_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13605_ deser_B.word_buffer\[41\] deser_B.serial_word\[41\] net123 VGND VGND VPWR
+ VPWR _00442_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_205_Right_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14585_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[15\]\[9\]
+ VGND VGND VPWR VPWR _11754_ sky130_fd_sc_hd__xor2_1
X_17373_ _04598_ _04628_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__xor2_1
X_29359_ clknet_leaf_231_clk _03157_ net140 VGND VGND VPWR VPWR C_out\[331\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19112_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[4\] _06176_ _06177_
+ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__a22o_1
XFILLER_186_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16324_ _03660_ _03673_ _03671_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__o21a_1
X_13536_ deser_A.shift_reg\[100\] deser_A.shift_reg\[101\] net129 VGND VGND VPWR VPWR
+ _00373_ sky130_fd_sc_hd__mux2_1
XFILLER_242_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19043_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.A_outs\[7\]\[1\] systolic_inst.B_outs\[7\]\[2\]
+ systolic_inst.B_outs\[7\]\[3\] VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__and4_1
X_16255_ _03633_ _03636_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13467_ deser_A.shift_reg\[31\] deser_A.shift_reg\[32\] deser_A.receiving VGND VGND
+ VPWR VPWR _00304_ sky130_fd_sc_hd__mux2_1
XFILLER_51_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15206_ _12302_ _12310_ VGND VGND VPWR VPWR _12311_ sky130_fd_sc_hd__or2_1
XFILLER_103_1251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16186_ _03527_ _03529_ _03528_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_149_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13398_ A_in\[107\] deser_A.word_buffer\[107\] _00003_ VGND VGND VPWR VPWR _00246_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15137_ net107 _12252_ VGND VGND VPWR VPWR _12253_ sky130_fd_sc_hd__nor2_1
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19945_ _06890_ _06940_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__xor2_1
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15068_ _12183_ _12184_ VGND VGND VPWR VPWR _12186_ sky130_fd_sc_hd__xnor2_1
XFILLER_218_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14019_ deser_B.shift_reg\[53\] deser_B.shift_reg\[54\] net125 VGND VGND VPWR VPWR
+ _00845_ sky130_fd_sc_hd__mux2_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19876_ _06856_ _06874_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__xor2_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18827_ _05934_ _05938_ _05941_ _05942_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__o211a_1
XFILLER_67_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18758_ _05879_ _05880_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__and2b_1
XFILLER_209_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17709_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[20\]
+ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__nand2_1
XFILLER_110_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18689_ _05806_ _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__nand2_1
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20720_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[15\]
+ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__nor2_1
XFILLER_212_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20651_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[5\]\[5\]
+ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__or2_1
XFILLER_32_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23370_ _09995_ _09996_ VGND VGND VPWR VPWR _09997_ sky130_fd_sc_hd__nand2_1
XFILLER_108_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20582_ _07481_ _07483_ _07513_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_134_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22321_ systolic_inst.A_outs\[2\]\[3\] systolic_inst.A_outs\[2\]\[4\] systolic_inst.B_outs\[2\]\[6\]
+ systolic_inst.B_outs\[2\]\[7\] VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__and4b_1
XFILLER_177_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25040_ net113 ser_C.shift_reg\[348\] VGND VGND VPWR VPWR _10990_ sky130_fd_sc_hd__and2_1
XFILLER_191_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22252_ systolic_inst.A_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[6\] _11265_ systolic_inst.A_outs\[2\]\[1\]
+ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_178_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21203_ _08069_ _08070_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__or2_1
X_22183_ _08927_ _08929_ VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__nor2_1
XFILLER_105_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_240_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21134_ systolic_inst.A_outs\[4\]\[5\] systolic_inst.B_outs\[4\]\[6\] _08003_ VGND
+ VGND VPWR VPWR _08004_ sky130_fd_sc_hd__and3_1
Xclkbuf_2_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_26991_ clknet_leaf_30_A_in_serial_clk _00789_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28730_ clknet_leaf_291_clk _02528_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[278\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21065_ _07935_ _07936_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__and2b_1
XFILLER_48_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25942_ systolic_inst.acc_wires\[13\]\[2\] C_out\[418\] net27 VGND VGND VPWR VPWR
+ _03244_ sky130_fd_sc_hd__mux2_1
XFILLER_235_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20016_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[6\]\[1\]
+ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__and2_1
XFILLER_47_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28661_ clknet_leaf_181_clk _02459_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[209\]
+ sky130_fd_sc_hd__dfrtp_1
X_25873_ systolic_inst.acc_wires\[10\]\[29\] C_out\[349\] net41 VGND VGND VPWR VPWR
+ _03175_ sky130_fd_sc_hd__mux2_1
XFILLER_115_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24824_ net113 ser_C.shift_reg\[240\] VGND VGND VPWR VPWR _10882_ sky130_fd_sc_hd__and2_1
X_27612_ clknet_leaf_321_clk _01410_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28592_ clknet_leaf_39_clk _02390_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[140\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_191_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24755_ C_out\[204\] net99 net79 ser_C.shift_reg\[204\] _10847_ VGND VGND VPWR VPWR
+ _02454_ sky130_fd_sc_hd__a221o_1
X_27543_ clknet_leaf_34_clk _01341_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_21967_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[15\]
+ VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__nand2_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23706_ _10320_ VGND VGND VPWR VPWR _10321_ sky130_fd_sc_hd__inv_2
XFILLER_226_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ _07791_ _07792_ _07754_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__a21oi_1
X_27474_ clknet_leaf_221_clk _01272_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_24686_ net112 ser_C.shift_reg\[171\] VGND VGND VPWR VPWR _10813_ sky130_fd_sc_hd__and2_1
XFILLER_242_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21898_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[3\]\[5\]
+ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__and2_1
XFILLER_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29213_ clknet_leaf_181_clk _03011_ net148 VGND VGND VPWR VPWR C_out\[185\] sky130_fd_sc_hd__dfrtp_1
X_23637_ _11269_ systolic_inst.B_outs\[0\]\[7\] _10120_ VGND VGND VPWR VPWR _10257_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_42_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26425_ clknet_leaf_8_clk _00232_ net134 VGND VGND VPWR VPWR A_in\[93\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20849_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[2\]
+ systolic_inst.A_outs\[4\]\[0\] VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__a22o_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29144_ clknet_leaf_165_clk _02942_ net150 VGND VGND VPWR VPWR C_out\[116\] sky130_fd_sc_hd__dfrtp_1
X_26356_ clknet_leaf_65_clk _00163_ net134 VGND VGND VPWR VPWR A_in\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14370_ _11518_ _11553_ VGND VGND VPWR VPWR _11554_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_189_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23568_ _10185_ _10188_ VGND VGND VPWR VPWR _10190_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_189_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_189_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25307_ ser_C.parallel_data\[480\] net102 net74 ser_C.shift_reg\[480\] _11123_ VGND
+ VGND VPWR VPWR _02730_ sky130_fd_sc_hd__a221o_1
X_13321_ A_in\[30\] deser_A.word_buffer\[30\] net91 VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__mux2_1
X_22519_ _09244_ _09245_ _09243_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__a21bo_1
XFILLER_6_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29075_ clknet_leaf_112_clk _02873_ net150 VGND VGND VPWR VPWR C_out\[47\] sky130_fd_sc_hd__dfrtp_1
XFILLER_196_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26287_ clknet_leaf_27_A_in_serial_clk _00095_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[85\]
+ sky130_fd_sc_hd__dfrtp_1
X_23499_ _10121_ _10122_ VGND VGND VPWR VPWR _10123_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_185_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ systolic_inst.A_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[2\] systolic_inst.B_outs\[12\]\[3\]
+ systolic_inst.B_outs\[12\]\[4\] VGND VGND VPWR VPWR _13037_ sky130_fd_sc_hd__and4_1
X_28026_ clknet_leaf_161_clk _01824_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_196_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25238_ net111 ser_C.shift_reg\[447\] VGND VGND VPWR VPWR _11089_ sky130_fd_sc_hd__and2_1
X_13252_ deser_A.word_buffer\[90\] deser_A.serial_word\[90\] net128 VGND VGND VPWR
+ VPWR _00100_ sky130_fd_sc_hd__mux2_1
XFILLER_108_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13183_ deser_A.word_buffer\[21\] deser_A.serial_word\[21\] net128 VGND VGND VPWR
+ VPWR _00031_ sky130_fd_sc_hd__mux2_1
X_25169_ C_out\[411\] net101 net73 ser_C.shift_reg\[411\] _11054_ VGND VGND VPWR VPWR
+ _02661_ sky130_fd_sc_hd__a221o_1
XFILLER_237_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17991_ _05141_ _05144_ _05182_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__or3_1
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19730_ _06702_ _06732_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__xnor2_1
X_28928_ clknet_leaf_266_clk _02726_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[476\]
+ sky130_fd_sc_hd__dfrtp_1
X_16942_ _04169_ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__or2_1
XFILLER_238_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19661_ _06664_ _06665_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__nand2_1
XFILLER_42_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28859_ clknet_leaf_335_clk _02657_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[407\]
+ sky130_fd_sc_hd__dfrtp_1
X_16873_ _04150_ _04152_ _04188_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18612_ systolic_inst.B_outs\[8\]\[5\] systolic_inst.A_outs\[8\]\[4\] VGND VGND VPWR
+ VPWR _05740_ sky130_fd_sc_hd__nand2_1
X_15824_ _12855_ _12857_ _12853_ VGND VGND VPWR VPWR _12863_ sky130_fd_sc_hd__a21bo_1
XFILLER_49_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19592_ _06619_ _06620_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__nand2_1
Xclkbuf_5_24__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_24__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18543_ _05638_ _05671_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15755_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[13\]\[1\]
+ VGND VGND VPWR VPWR _12804_ sky130_fd_sc_hd__or2_1
XFILLER_46_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14706_ systolic_inst.acc_wires\[15\]\[24\] systolic_inst.acc_wires\[15\]\[25\] systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _11858_ sky130_fd_sc_hd__o21a_1
XFILLER_221_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18474_ _05588_ _05605_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__xor2_1
XFILLER_178_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15686_ _12736_ _12737_ VGND VGND VPWR VPWR _12740_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_174_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ systolic_inst.A_outs\[10\]\[3\] systolic_inst.A_outs\[10\]\[4\] systolic_inst.B_outs\[10\]\[6\]
+ systolic_inst.B_outs\[10\]\[7\] VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_99_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14637_ _11783_ _11790_ _11796_ _11789_ VGND VGND VPWR VPWR _11799_ sky130_fd_sc_hd__a211o_1
XFILLER_53_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14568_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[15\]\[6\]
+ VGND VGND VPWR VPWR _11740_ sky130_fd_sc_hd__or2_1
XFILLER_53_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17356_ systolic_inst.A_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[2\] systolic_inst.B_outs\[10\]\[6\]
+ systolic_inst.B_outs\[10\]\[7\] VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__and4b_1
XFILLER_144_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16307_ _03686_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__nor2_1
XFILLER_53_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13519_ deser_A.shift_reg\[83\] deser_A.shift_reg\[84\] net129 VGND VGND VPWR VPWR
+ _00356_ sky130_fd_sc_hd__mux2_1
XFILLER_179_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14499_ _11676_ _11677_ _11678_ VGND VGND VPWR VPWR _11679_ sky130_fd_sc_hd__a21oi_1
X_17287_ _04540_ _04541_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__nand3_2
Xclkload302 clknet_leaf_186_clk VGND VGND VPWR VPWR clkload302/Y sky130_fd_sc_hd__clkinv_8
XFILLER_105_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload313 clknet_leaf_153_clk VGND VGND VPWR VPWR clkload313/Y sky130_fd_sc_hd__inv_6
XFILLER_173_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload10 clknet_5_11__leaf_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__inv_8
XFILLER_220_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload324 clknet_leaf_148_clk VGND VGND VPWR VPWR clkload324/Y sky130_fd_sc_hd__clkinv_4
Xclkload21 clknet_5_25__leaf_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__inv_12
X_19026_ systolic_inst.B_outs\[6\]\[7\] systolic_inst.B_outs\[2\]\[7\] net120 VGND
+ VGND VPWR VPWR _01473_ sky130_fd_sc_hd__mux2_1
Xclkload335 clknet_leaf_163_clk VGND VGND VPWR VPWR clkload335/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_174_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload32 clknet_leaf_337_clk VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__clkinv_4
X_16238_ _03617_ _03618_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__xnor2_1
Xclkload43 clknet_leaf_288_clk VGND VGND VPWR VPWR clkload43/X sky130_fd_sc_hd__clkbuf_8
Xclkload346 clknet_leaf_19_A_in_serial_clk VGND VGND VPWR VPWR clkload346/X sky130_fd_sc_hd__clkbuf_4
XFILLER_133_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload357 clknet_leaf_9_A_in_serial_clk VGND VGND VPWR VPWR clkload357/Y sky130_fd_sc_hd__inv_6
Xclkload54 clknet_leaf_314_clk VGND VGND VPWR VPWR clkload54/Y sky130_fd_sc_hd__inv_6
Xclkload368 clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR clkload368/Y sky130_fd_sc_hd__inv_6
Xclkload65 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload65/Y sky130_fd_sc_hd__inv_6
Xclkload379 clknet_leaf_20_B_in_serial_clk VGND VGND VPWR VPWR clkload379/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_115_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload76 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload76/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_90_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16169_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[8\] VGND
+ VGND VPWR VPWR _03554_ sky130_fd_sc_hd__and2_1
Xclkload87 clknet_leaf_310_clk VGND VGND VPWR VPWR clkload87/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_90_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload98 clknet_leaf_306_clk VGND VGND VPWR VPWR clkload98/Y sky130_fd_sc_hd__inv_8
XFILLER_170_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19928_ systolic_inst.B_outs\[6\]\[6\] systolic_inst.A_outs\[6\]\[6\] _11278_ systolic_inst.A_outs\[6\]\[5\]
+ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_151_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19859_ systolic_inst.B_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[7\]
+ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__and3_1
XFILLER_112_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22870_ net109 systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[8\] VGND
+ VGND VPWR VPWR _09551_ sky130_fd_sc_hd__and2_1
XFILLER_151_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21821_ _08623_ _08624_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__nand2_1
XFILLER_71_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24540_ net113 ser_C.shift_reg\[98\] VGND VGND VPWR VPWR _10740_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_233_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21752_ systolic_inst.A_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[5\] systolic_inst.B_outs\[3\]\[6\]
+ systolic_inst.B_outs\[3\]\[7\] VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__and4b_1
XFILLER_149_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_233_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_233_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20703_ _07618_ _07619_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__nor2_1
X_24471_ C_out\[62\] net100 net82 ser_C.shift_reg\[62\] _10705_ VGND VGND VPWR VPWR
+ _02312_ sky130_fd_sc_hd__a221o_1
XFILLER_184_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21683_ systolic_inst.A_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[6\]
+ systolic_inst.B_outs\[3\]\[7\] VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_43_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26210_ clknet_leaf_13_A_in_serial_clk _00018_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23422_ _10038_ _10045_ VGND VGND VPWR VPWR _10048_ sky130_fd_sc_hd__xor2_1
X_20634_ _07560_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__inv_2
X_27190_ clknet_leaf_247_clk _00988_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload4 clknet_5_4__leaf_clk VGND VGND VPWR VPWR clkload4/X sky130_fd_sc_hd__clkbuf_8
X_26141_ deser_B.serial_word\[96\] deser_B.shift_reg\[96\] net56 VGND VGND VPWR VPWR
+ _03443_ sky130_fd_sc_hd__mux2_1
XFILLER_138_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23353_ _09979_ _09980_ VGND VGND VPWR VPWR _09981_ sky130_fd_sc_hd__xor2_1
XFILLER_20_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20565_ _07469_ _07496_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__nand2b_1
XFILLER_50_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22304_ _09047_ VGND VGND VPWR VPWR _09048_ sky130_fd_sc_hd__inv_2
X_26072_ deser_B.serial_word\[27\] deser_B.shift_reg\[27\] net56 VGND VGND VPWR VPWR
+ _03374_ sky130_fd_sc_hd__mux2_1
X_23284_ systolic_inst.A_outs\[0\]\[7\] systolic_inst.A_shift\[0\]\[7\] net117 VGND
+ VGND VPWR VPWR _01913_ sky130_fd_sc_hd__mux2_1
X_20496_ _07322_ _07429_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__nor2_1
XFILLER_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25023_ C_out\[338\] net97 net77 ser_C.shift_reg\[338\] _10981_ VGND VGND VPWR VPWR
+ _02588_ sky130_fd_sc_hd__a221o_1
X_22235_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[7\] _08980_ net122
+ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__mux2_1
XFILLER_156_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22166_ _08911_ _08912_ net122 VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_7_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21117_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[10\] _07987_ net117
+ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__mux2_1
X_22097_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[1\]
+ systolic_inst.B_outs\[2\]\[0\] VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__a22o_1
X_26974_ clknet_leaf_24_A_in_serial_clk _00772_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_28713_ clknet_leaf_325_clk _02511_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[261\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_219_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21048_ _07877_ _07919_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__nand2_1
X_25925_ systolic_inst.acc_wires\[12\]\[17\] C_out\[401\] net18 VGND VGND VPWR VPWR
+ _03227_ sky130_fd_sc_hd__mux2_1
XFILLER_87_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29693_ clknet_leaf_8_clk _03488_ VGND VGND VPWR VPWR systolic_inst.A_shift\[30\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28644_ clknet_leaf_207_clk _02442_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[192\]
+ sky130_fd_sc_hd__dfrtp_1
X_13870_ deser_A.serial_word\[31\] deser_A.shift_reg\[31\] net58 VGND VGND VPWR VPWR
+ _00696_ sky130_fd_sc_hd__mux2_1
XFILLER_235_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25856_ systolic_inst.acc_wires\[10\]\[12\] C_out\[332\] net12 VGND VGND VPWR VPWR
+ _03158_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_178_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24807_ C_out\[230\] net99 net79 ser_C.shift_reg\[230\] _10873_ VGND VGND VPWR VPWR
+ _02480_ sky130_fd_sc_hd__a221o_1
XFILLER_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28575_ clknet_leaf_173_clk _02373_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_22999_ _09622_ _09674_ VGND VGND VPWR VPWR _09676_ sky130_fd_sc_hd__xor2_1
XFILLER_131_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25787_ systolic_inst.acc_wires\[8\]\[7\] C_out\[263\] net22 VGND VGND VPWR VPWR
+ _03089_ sky130_fd_sc_hd__mux2_1
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15540_ _12595_ _12596_ VGND VGND VPWR VPWR _12598_ sky130_fd_sc_hd__xor2_1
X_27526_ clknet_leaf_236_clk _01324_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_24738_ net112 ser_C.shift_reg\[197\] VGND VGND VPWR VPWR _10839_ sky130_fd_sc_hd__and2_1
XFILLER_167_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15471_ _12507_ _12529_ _12530_ VGND VGND VPWR VPWR _12531_ sky130_fd_sc_hd__nor3_1
XFILLER_70_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24669_ C_out\[161\] net103 net76 ser_C.shift_reg\[161\] _10804_ VGND VGND VPWR VPWR
+ _02411_ sky130_fd_sc_hd__a221o_1
X_27457_ clknet_leaf_238_clk _01255_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_230_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14422_ _11560_ _11568_ _11567_ VGND VGND VPWR VPWR _11605_ sky130_fd_sc_hd__a21bo_1
X_17210_ net107 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[2\] _04471_
+ _04472_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__a22o_1
XFILLER_202_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26408_ clknet_leaf_4_clk _00215_ net131 VGND VGND VPWR VPWR A_in\[76\] sky130_fd_sc_hd__dfrtp_1
X_18190_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] _05369_
+ _05375_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__a22o_1
XFILLER_156_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27388_ clknet_leaf_337_clk _01186_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_29127_ clknet_leaf_173_clk _02925_ net148 VGND VGND VPWR VPWR C_out\[99\] sky130_fd_sc_hd__dfrtp_1
X_17141_ net62 _04427_ _04428_ systolic_inst.acc_wires\[11\]\[25\] net105 VGND VGND
+ VPWR VPWR _01259_ sky130_fd_sc_hd__a32o_1
XFILLER_50_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14353_ _11486_ _11495_ _11494_ VGND VGND VPWR VPWR _11538_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26339_ clknet_leaf_59_clk _00146_ net137 VGND VGND VPWR VPWR A_in\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_195_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13304_ A_in\[13\] deser_A.word_buffer\[13\] net93 VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__mux2_1
XFILLER_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17072_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[15\]
+ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__and2_1
X_29058_ clknet_leaf_108_clk _02856_ net151 VGND VGND VPWR VPWR C_out\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_171_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14284_ _11469_ _11470_ VGND VGND VPWR VPWR _11471_ sky130_fd_sc_hd__nor2_1
XFILLER_156_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28009_ clknet_leaf_149_clk _01807_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_16023_ _12996_ _12999_ _13018_ VGND VGND VPWR VPWR _13021_ sky130_fd_sc_hd__nand3_1
X_13235_ deser_A.word_buffer\[73\] deser_A.serial_word\[73\] net127 VGND VGND VPWR
+ VPWR _00083_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13166_ deser_A.word_buffer\[4\] deser_A.serial_word\[4\] net127 VGND VGND VPWR VPWR
+ _00014_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17974_ _05164_ _05165_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19713_ _06712_ _06715_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__xor2_1
X_16925_ _04238_ _04239_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__xor2_1
XFILLER_46_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19644_ systolic_inst.A_outs\[6\]\[1\] systolic_inst.B_outs\[6\]\[2\] systolic_inst.B_outs\[6\]\[3\]
+ systolic_inst.A_outs\[6\]\[0\] VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__a22oi_1
XFILLER_20_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16856_ _04170_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_122_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15807_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[13\]\[8\]
+ _12845_ _12847_ VGND VGND VPWR VPWR _12848_ sky130_fd_sc_hd__a211o_1
XFILLER_19_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19575_ net62 _06605_ _06606_ systolic_inst.acc_wires\[7\]\[25\] net106 VGND VGND
+ VPWR VPWR _01515_ sky130_fd_sc_hd__a32o_1
XFILLER_20_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16787_ systolic_inst.A_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[5\] _04069_ _04068_
+ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__a31oi_1
X_13999_ deser_B.shift_reg\[33\] deser_B.shift_reg\[34\] deser_B.receiving VGND VGND
+ VPWR VPWR _00825_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18526_ _05603_ _05631_ _05630_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15738_ _12738_ _12766_ _12767_ VGND VGND VPWR VPWR _12790_ sky130_fd_sc_hd__o21ai_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18457_ _05586_ _05588_ _05569_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15669_ _12688_ _12690_ _12689_ VGND VGND VPWR VPWR _12723_ sky130_fd_sc_hd__o21ba_1
XFILLER_60_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17408_ _04638_ _04663_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__xnor2_1
X_18388_ _05536_ _05539_ _05538_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__o21a_1
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17339_ _04595_ _04596_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__xor2_1
XFILLER_88_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20350_ systolic_inst.B_outs\[5\]\[1\] systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[5\]
+ systolic_inst.A_outs\[5\]\[6\] VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_116_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload110 clknet_leaf_285_clk VGND VGND VPWR VPWR clkload110/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload121 clknet_leaf_294_clk VGND VGND VPWR VPWR clkload121/Y sky130_fd_sc_hd__clkinv_2
Xclkload132 clknet_leaf_267_clk VGND VGND VPWR VPWR clkload132/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_161_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload143 clknet_leaf_258_clk VGND VGND VPWR VPWR clkload143/X sky130_fd_sc_hd__clkbuf_8
XFILLER_220_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload154 clknet_leaf_202_clk VGND VGND VPWR VPWR clkload154/Y sky130_fd_sc_hd__clkinvlp_4
X_19009_ _06092_ _06096_ _06097_ net61 VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_77_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20281_ _07213_ _07219_ _07221_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__and3_1
Xclkload165 clknet_leaf_232_clk VGND VGND VPWR VPWR clkload165/Y sky130_fd_sc_hd__inv_8
XFILLER_31_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload176 clknet_leaf_197_clk VGND VGND VPWR VPWR clkload176/Y sky130_fd_sc_hd__inv_4
Xclkload187 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload187/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_226_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22020_ _08796_ _08798_ VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__xor2_1
Xclkload198 clknet_leaf_62_clk VGND VGND VPWR VPWR clkload198/Y sky130_fd_sc_hd__clkinv_4
XFILLER_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_222_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23971_ systolic_inst.B_shift\[13\]\[5\] B_in\[45\] _00008_ VGND VGND VPWR VPWR _10511_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_239_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25710_ systolic_inst.acc_wires\[5\]\[26\] C_out\[186\] net46 VGND VGND VPWR VPWR
+ _03012_ sky130_fd_sc_hd__mux2_1
X_22922_ _09592_ _09600_ VGND VGND VPWR VPWR _09601_ sky130_fd_sc_hd__nand2_1
XFILLER_25_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26690_ clknet_leaf_32_B_in_serial_clk _00493_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_235_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_235_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_235_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25641_ systolic_inst.acc_wires\[3\]\[21\] C_out\[117\] net50 VGND VGND VPWR VPWR
+ _02943_ sky130_fd_sc_hd__mux2_1
XFILLER_216_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22853_ _09530_ _09532_ VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__xor2_1
XFILLER_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21804_ _08607_ _08608_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__or2_1
X_25572_ systolic_inst.acc_wires\[1\]\[16\] C_out\[48\] net35 VGND VGND VPWR VPWR
+ _02874_ sky130_fd_sc_hd__mux2_1
X_28360_ clknet_leaf_75_clk _02158_ VGND VGND VPWR VPWR systolic_inst.B_shift\[22\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_22784_ _09464_ _09465_ _09435_ VGND VGND VPWR VPWR _09467_ sky130_fd_sc_hd__a21o_1
XFILLER_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24523_ C_out\[88\] net100 net82 ser_C.shift_reg\[88\] _10731_ VGND VGND VPWR VPWR
+ _02338_ sky130_fd_sc_hd__a221o_1
XFILLER_227_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27311_ clknet_leaf_292_clk _01109_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_21735_ _08540_ _08541_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__nand2_1
X_28291_ clknet_leaf_72_clk _02089_ VGND VGND VPWR VPWR systolic_inst.B_shift\[19\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24454_ net114 ser_C.shift_reg\[55\] VGND VGND VPWR VPWR _10697_ sky130_fd_sc_hd__and2_1
X_27242_ clknet_leaf_278_clk _01040_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_21666_ _08473_ _08474_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__nor2_1
XFILLER_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23405_ _10024_ _10029_ VGND VGND VPWR VPWR _10031_ sky130_fd_sc_hd__xor2_1
X_20617_ _07536_ _07537_ _07546_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__a21oi_1
X_27173_ clknet_leaf_254_clk _00971_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24385_ C_out\[19\] net104 _10643_ ser_C.shift_reg\[19\] _10662_ VGND VGND VPWR VPWR
+ _02269_ sky130_fd_sc_hd__a221o_1
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21597_ _08405_ _08406_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__nand2_1
X_26124_ deser_B.serial_word\[79\] deser_B.shift_reg\[79\] net55 VGND VGND VPWR VPWR
+ _03426_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23336_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[4\] _09964_ net121
+ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__mux2_1
X_20548_ _07480_ _07479_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__and2b_1
XFILLER_123_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26055_ deser_B.serial_word\[10\] deser_B.shift_reg\[10\] net55 VGND VGND VPWR VPWR
+ _03357_ sky130_fd_sc_hd__mux2_1
XFILLER_153_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23267_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[30\]
+ VGND VGND VPWR VPWR _09910_ sky130_fd_sc_hd__nand2_1
XFILLER_197_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20479_ _07411_ _07412_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__xor2_1
XFILLER_106_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25006_ net111 ser_C.shift_reg\[331\] VGND VGND VPWR VPWR _10973_ sky130_fd_sc_hd__and2_1
XFILLER_193_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22218_ _08960_ _08963_ VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23198_ _09850_ _09851_ VGND VGND VPWR VPWR _09852_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22149_ _08879_ _08896_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__xor2_1
XFILLER_239_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14971_ _12074_ _12091_ VGND VGND VPWR VPWR _12092_ sky130_fd_sc_hd__xor2_1
X_26957_ clknet_leaf_1_A_in_serial_clk _00755_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_16710_ systolic_inst.A_outs\[11\]\[2\] systolic_inst.B_outs\[11\]\[5\] VGND VGND
+ VPWR VPWR _04032_ sky130_fd_sc_hd__nand2_1
X_25908_ systolic_inst.acc_wires\[12\]\[0\] C_out\[384\] net20 VGND VGND VPWR VPWR
+ _03210_ sky130_fd_sc_hd__mux2_1
X_13922_ deser_A.serial_word\[83\] deser_A.shift_reg\[83\] net57 VGND VGND VPWR VPWR
+ _00748_ sky130_fd_sc_hd__mux2_1
X_29676_ clknet_leaf_32_B_in_serial_clk _03471_ net134 VGND VGND VPWR VPWR deser_B.serial_word\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_17690_ net60 _04922_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__nor2_1
XFILLER_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26888_ clknet_leaf_8_A_in_serial_clk _00686_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28627_ clknet_leaf_146_clk _02425_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[175\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16641_ systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[5\]
+ systolic_inst.B_outs\[11\]\[0\] VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__a22oi_1
XFILLER_235_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25839_ systolic_inst.acc_wires\[9\]\[27\] C_out\[315\] net13 VGND VGND VPWR VPWR
+ _03141_ sky130_fd_sc_hd__mux2_1
X_13853_ deser_A.serial_word\[14\] deser_A.shift_reg\[14\] net58 VGND VGND VPWR VPWR
+ _00679_ sky130_fd_sc_hd__mux2_1
XFILLER_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19360_ _06375_ _06388_ _06386_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__o21a_1
XFILLER_204_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28558_ clknet_leaf_168_clk _02356_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_16572_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[31\]
+ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13784_ B_in\[91\] deser_B.word_buffer\[91\] net89 VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__mux2_1
XFILLER_215_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18311_ net106 systolic_inst.acc_wires\[9\]\[17\] net66 _05478_ VGND VGND VPWR VPWR
+ _01379_ sky130_fd_sc_hd__a22o_1
XFILLER_43_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15523_ _12574_ _12580_ VGND VGND VPWR VPWR _12581_ sky130_fd_sc_hd__xnor2_1
X_27509_ clknet_leaf_230_clk _01307_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_204_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19291_ _06349_ _06352_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__xor2_1
XFILLER_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28489_ clknet_leaf_116_clk _02287_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[9\]\[8\]
+ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__nand2_1
X_15454_ _12485_ _12513_ VGND VGND VPWR VPWR _12514_ sky130_fd_sc_hd__xor2_1
XFILLER_175_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14405_ _11518_ _11587_ VGND VGND VPWR VPWR _11588_ sky130_fd_sc_hd__nor2_1
XFILLER_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18173_ _05357_ _05358_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__and2b_1
XFILLER_141_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15385_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[2\] _12447_ VGND
+ VGND VPWR VPWR _12449_ sky130_fd_sc_hd__a21o_1
XFILLER_15_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17124_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__inv_2
XFILLER_50_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14336_ _11478_ _11520_ VGND VGND VPWR VPWR _11521_ sky130_fd_sc_hd__and2_1
XFILLER_184_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14267_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[6\] _11453_ VGND
+ VGND VPWR VPWR _11454_ sky130_fd_sc_hd__and3_1
X_17055_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[11\]\[13\]
+ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_111_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16006_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[2\] VGND VGND
+ VPWR VPWR _13004_ sky130_fd_sc_hd__and2_1
X_13218_ deser_A.word_buffer\[56\] deser_A.serial_word\[56\] net128 VGND VGND VPWR
+ VPWR _00066_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14198_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[5\] VGND VGND
+ VPWR VPWR _11387_ sky130_fd_sc_hd__nand2_1
XFILLER_98_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13149_ ser_C.bit_idx\[8\] _11300_ net7 VGND VGND VPWR VPWR _11301_ sky130_fd_sc_hd__a21bo_1
XFILLER_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17957_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[7\]
+ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__o21ai_2
XFILLER_22_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16908_ _04155_ _04161_ _04191_ _04189_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__o31a_1
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17888_ _05079_ _05082_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__xor2_1
X_19627_ systolic_inst.B_outs\[5\]\[7\] systolic_inst.B_outs\[1\]\[7\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__mux2_1
X_16839_ _04122_ _04089_ _04121_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__or3b_1
XFILLER_96_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19558_ _06591_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__inv_2
XFILLER_20_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18509_ _05637_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__nor2_1
XFILLER_178_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19489_ net105 systolic_inst.acc_wires\[7\]\[12\] _06531_ _06533_ VGND VGND VPWR
+ VPWR _01502_ sky130_fd_sc_hd__a22o_1
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21520_ _08311_ _08332_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_118_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21451_ _11258_ systolic_inst.acc_wires\[4\]\[29\] net63 _08286_ VGND VGND VPWR VPWR
+ _01711_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20402_ systolic_inst.B_outs\[5\]\[7\] _07338_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__nand2_1
XFILLER_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24170_ systolic_inst.A_shift\[26\]\[1\] net70 _10505_ systolic_inst.A_shift\[27\]\[1\]
+ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_228_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21382_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[19\]
+ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_21_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23121_ _09784_ _09785_ VGND VGND VPWR VPWR _09786_ sky130_fd_sc_hd__and2_1
X_20333_ _07265_ _07266_ _07269_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__a21o_1
XFILLER_135_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23052_ _09725_ _09726_ VGND VGND VPWR VPWR _09727_ sky130_fd_sc_hd__nor2_1
XFILLER_66_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20264_ _07192_ _07194_ _07205_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__and3_1
XFILLER_192_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22003_ _08782_ _08783_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__and2_1
XFILLER_131_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27860_ clknet_leaf_215_clk _01658_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_192_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20195_ _07154_ _07158_ _07155_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26811_ clknet_leaf_75_clk _00613_ net144 VGND VGND VPWR VPWR B_in\[83\] sky130_fd_sc_hd__dfrtp_1
XFILLER_88_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27791_ clknet_leaf_41_clk _01589_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_29_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29530_ clknet_leaf_262_clk _03328_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[502\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_217_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26742_ clknet_leaf_97_clk _00544_ net153 VGND VGND VPWR VPWR B_in\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_116_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23954_ systolic_inst.B_shift\[11\]\[1\] net70 net83 systolic_inst.B_shift\[15\]\[1\]
+ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__a22o_1
XFILLER_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22905_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[9\] _09584_ net122
+ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__mux2_1
X_29461_ clknet_leaf_331_clk _03259_ net136 VGND VGND VPWR VPWR C_out\[433\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23885_ _10462_ _10465_ _10468_ _10471_ VGND VGND VPWR VPWR _10472_ sky130_fd_sc_hd__o31a_1
X_26673_ clknet_leaf_9_B_in_serial_clk _00476_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28412_ clknet_leaf_60_clk _02210_ VGND VGND VPWR VPWR systolic_inst.B_shift\[23\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25624_ systolic_inst.acc_wires\[3\]\[4\] C_out\[100\] net48 VGND VGND VPWR VPWR
+ _02926_ sky130_fd_sc_hd__mux2_1
X_22836_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] _09515_ VGND
+ VGND VPWR VPWR _09517_ sky130_fd_sc_hd__a21o_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29392_ clknet_leaf_241_clk _03190_ net145 VGND VGND VPWR VPWR C_out\[364\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28343_ clknet_leaf_343_clk _02141_ VGND VGND VPWR VPWR systolic_inst.A_shift\[25\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25555_ systolic_inst.acc_wires\[0\]\[31\] C_out\[31\] net36 VGND VGND VPWR VPWR
+ _02857_ sky130_fd_sc_hd__mux2_1
X_22767_ systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[5\] systolic_inst.A_outs\[1\]\[6\]
+ systolic_inst.B_outs\[1\]\[0\] VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__a22oi_1
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24506_ net113 ser_C.shift_reg\[81\] VGND VGND VPWR VPWR _10723_ sky130_fd_sc_hd__and2_1
XFILLER_213_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21718_ _08523_ _08524_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__nor2_1
XFILLER_40_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25486_ _11279_ _11219_ _11221_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_213_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28274_ clknet_leaf_130_clk _02072_ VGND VGND VPWR VPWR systolic_inst.B_shift\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22698_ _09383_ _09384_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__or2_1
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27225_ clknet_leaf_312_clk _01023_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_24437_ C_out\[45\] _11302_ net81 ser_C.shift_reg\[45\] _10688_ VGND VGND VPWR VPWR
+ _02295_ sky130_fd_sc_hd__a221o_1
X_21649_ systolic_inst.A_outs\[3\]\[2\] systolic_inst.B_outs\[3\]\[5\] _08421_ _08420_
+ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__a31oi_1
XFILLER_240_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15170_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[14\]\[4\]
+ VGND VGND VPWR VPWR _12280_ sky130_fd_sc_hd__and2_1
X_24368_ net7 ser_C.shift_reg\[12\] VGND VGND VPWR VPWR _10654_ sky130_fd_sc_hd__and2_1
XFILLER_165_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27156_ clknet_leaf_294_clk _00954_ net138 VGND VGND VPWR VPWR systolic_inst.B_outs\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_240_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14121_ systolic_inst.A_shift\[21\]\[5\] net71 _11333_ A_in\[93\] VGND VGND VPWR
+ VPWR _00943_ sky130_fd_sc_hd__a22o_1
X_23319_ systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[3\]
+ systolic_inst.B_outs\[0\]\[1\] VGND VGND VPWR VPWR _09948_ sky130_fd_sc_hd__a22o_1
X_26107_ deser_B.serial_word\[62\] deser_B.shift_reg\[62\] net56 VGND VGND VPWR VPWR
+ _03409_ sky130_fd_sc_hd__mux2_1
XFILLER_4_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27087_ clknet_leaf_33_B_in_serial_clk _00885_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24299_ systolic_inst.A_shift\[12\]\[5\] A_in\[53\] net59 VGND VGND VPWR VPWR _10623_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14052_ deser_B.shift_reg\[86\] deser_B.shift_reg\[87\] net125 VGND VGND VPWR VPWR
+ _00878_ sky130_fd_sc_hd__mux2_1
X_26038_ systolic_inst.B_outs\[15\]\[2\] systolic_inst.B_outs\[11\]\[2\] net118 VGND
+ VGND VPWR VPWR _03340_ sky130_fd_sc_hd__mux2_1
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18860_ net63 _05970_ _05971_ systolic_inst.acc_wires\[8\]\[9\] net108 VGND VGND
+ VPWR VPWR _01435_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_160_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17811_ _05007_ _05008_ _05009_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__a21o_1
XFILLER_239_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18791_ _05694_ _05832_ _05906_ _05904_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__a31oi_1
X_27989_ clknet_leaf_100_clk _01787_ net152 VGND VGND VPWR VPWR systolic_inst.B_outs\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_82_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17742_ _04961_ _04963_ _04966_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__a21oi_2
X_14954_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[7\] VGND VGND
+ VPWR VPWR _12075_ sky130_fd_sc_hd__nand2_4
XFILLER_36_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13905_ deser_A.serial_word\[66\] deser_A.shift_reg\[66\] net57 VGND VGND VPWR VPWR
+ _00731_ sky130_fd_sc_hd__mux2_1
X_29659_ clknet_leaf_7_B_in_serial_clk _03454_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_17673_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[10\]\[13\]
+ _04902_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__a21oi_1
XFILLER_130_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_195_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_195_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14885_ systolic_inst.A_outs\[14\]\[1\] systolic_inst.B_outs\[14\]\[6\] _12007_ VGND
+ VGND VPWR VPWR _12008_ sky130_fd_sc_hd__and3_1
XFILLER_223_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19412_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[7\]\[2\]
+ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__and2_1
XFILLER_1_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16624_ systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[3\] systolic_inst.A_outs\[11\]\[4\]
+ systolic_inst.B_outs\[11\]\[0\] VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__a22o_1
XFILLER_210_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13836_ deser_B.bit_idx\[5\] _11327_ _11321_ _11285_ VGND VGND VPWR VPWR _00663_
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap70 net71 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_16
Xmax_cap81 net82 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_16
XFILLER_223_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19343_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[12\] _06403_ net119
+ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__mux2_1
Xmax_cap92 _00003_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_8
XFILLER_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16555_ _03895_ _03903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__nor2_1
X_13767_ B_in\[74\] deser_B.word_buffer\[74\] net90 VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__mux2_1
XFILLER_204_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15506_ _12564_ _12563_ VGND VGND VPWR VPWR _12565_ sky130_fd_sc_hd__nand2b_1
X_19274_ _06300_ _06301_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__nand2_1
XFILLER_91_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16486_ _03846_ _03845_ systolic_inst.acc_wires\[12\]\[16\] net108 VGND VGND VPWR
+ VPWR _01186_ sky130_fd_sc_hd__a2bb2o_1
X_13698_ B_in\[5\] deser_B.word_buffer\[5\] net84 VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18225_ _05403_ _05404_ _05396_ _05400_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__a211o_1
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15437_ _12488_ _12496_ VGND VGND VPWR VPWR _12498_ sky130_fd_sc_hd__xor2_1
XFILLER_54_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18156_ _05313_ _05317_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15368_ systolic_inst.B_outs\[12\]\[4\] systolic_inst.B_outs\[8\]\[4\] net115 VGND
+ VGND VPWR VPWR _01086_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17107_ _04396_ _04398_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__or3_1
XFILLER_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14319_ _11474_ _11504_ VGND VGND VPWR VPWR _11505_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_74_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18087_ _05222_ _05240_ _05239_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__o21a_1
X_15299_ _12387_ _12388_ _12389_ VGND VGND VPWR VPWR _12391_ sky130_fd_sc_hd__or3_1
XFILLER_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17038_ net105 systolic_inst.acc_wires\[11\]\[10\] net69 _04340_ VGND VGND VPWR VPWR
+ _01244_ sky130_fd_sc_hd__a22o_1
XFILLER_176_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18989_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[28\]
+ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__or2_1
XFILLER_140_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_219_Right_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20951_ _07801_ _07824_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_186_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_186_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_227_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23670_ _10260_ _10288_ _10264_ VGND VGND VPWR VPWR _10289_ sky130_fd_sc_hd__o21a_1
XFILLER_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_217_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20882_ systolic_inst.B_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[2\] systolic_inst.B_outs\[4\]\[2\]
+ systolic_inst.A_outs\[4\]\[3\] VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__nand4_2
XFILLER_54_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22621_ _09326_ _09330_ _09332_ net60 VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_27_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25340_ net112 ser_C.shift_reg\[498\] VGND VGND VPWR VPWR _11140_ sky130_fd_sc_hd__and2_1
XFILLER_34_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22552_ _09275_ _09276_ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21503_ _08314_ _08315_ _08304_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__a21o_1
XFILLER_179_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25271_ ser_C.parallel_data\[462\] net102 net74 ser_C.shift_reg\[462\] _11105_ VGND
+ VGND VPWR VPWR _02712_ sky130_fd_sc_hd__a221o_1
X_22483_ _09217_ VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__inv_2
XFILLER_166_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27010_ clknet_leaf_17_B_in_serial_clk _00808_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_24222_ _10596_ systolic_inst.A_shift\[19\]\[2\] net70 VGND VGND VPWR VPWR _02172_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21434_ _11258_ systolic_inst.acc_wires\[4\]\[26\] net63 _08272_ VGND VGND VPWR VPWR
+ _01708_ sky130_fd_sc_hd__a22o_1
XFILLER_148_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24153_ systolic_inst.A_shift\[28\]\[0\] A_in\[96\] net59 VGND VGND VPWR VPWR _10578_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21365_ _08212_ _08213_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_110_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_190_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23104_ _09771_ VGND VGND VPWR VPWR _09772_ sky130_fd_sc_hd__inv_2
XFILLER_174_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20316_ _07236_ _07238_ _07237_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__o21bai_1
XFILLER_107_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24084_ systolic_inst.B_shift\[2\]\[3\] _11332_ net83 systolic_inst.B_shift\[6\]\[3\]
+ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__a22o_1
X_28961_ clknet_leaf_257_clk _02759_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[509\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_162_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21296_ net63 _08152_ _08154_ systolic_inst.acc_wires\[4\]\[6\] net108 VGND VGND
+ VPWR VPWR _01688_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_57_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23035_ _09679_ _09684_ _09709_ VGND VGND VPWR VPWR _09711_ sky130_fd_sc_hd__o21ai_1
X_27912_ clknet_leaf_135_clk _01710_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_20247_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[1\]
+ systolic_inst.A_outs\[5\]\[2\] VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_57_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28892_ clknet_leaf_286_clk _02690_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[440\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_107_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_206_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27843_ clknet_leaf_206_clk _01641_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20178_ _07145_ _07146_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__or2_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_202_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27774_ clknet_leaf_179_clk _01572_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_5_5__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_198_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24986_ net111 ser_C.shift_reg\[321\] VGND VGND VPWR VPWR _10963_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_198_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29513_ clknet_leaf_260_clk _03311_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[485\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26725_ clknet_leaf_0_B_in_serial_clk _00528_ net134 VGND VGND VPWR VPWR deser_B.word_buffer\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_177_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_177_clk
+ sky130_fd_sc_hd__clkbuf_8
X_23937_ _10497_ systolic_inst.B_shift\[10\]\[0\] _11332_ VGND VGND VPWR VPWR _01986_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_24_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29444_ clknet_leaf_301_clk _03242_ net141 VGND VGND VPWR VPWR C_out\[416\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_194_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26656_ clknet_leaf_28_B_in_serial_clk _00459_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_14670_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[21\]
+ VGND VGND VPWR VPWR _11827_ sky130_fd_sc_hd__xnor2_2
X_23868_ _10451_ _10455_ _10452_ VGND VGND VPWR VPWR _10458_ sky130_fd_sc_hd__a21bo_1
XFILLER_72_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25607_ systolic_inst.acc_wires\[2\]\[19\] C_out\[83\] net52 VGND VGND VPWR VPWR
+ _02909_ sky130_fd_sc_hd__mux2_1
X_13621_ deser_B.word_buffer\[57\] deser_B.serial_word\[57\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__mux2_1
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22819_ _09487_ _09499_ VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__nand2_1
X_29375_ clknet_leaf_236_clk _03173_ net145 VGND VGND VPWR VPWR C_out\[347\] sky130_fd_sc_hd__dfrtp_1
XFILLER_207_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26587_ clknet_leaf_0_A_in_serial_clk _00390_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[117\]
+ sky130_fd_sc_hd__dfrtp_1
X_23799_ _10388_ _10394_ _10395_ VGND VGND VPWR VPWR _10400_ sky130_fd_sc_hd__o21ba_1
XFILLER_129_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16340_ _03717_ _03718_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__nand2_1
X_28326_ clknet_leaf_2_clk _02124_ VGND VGND VPWR VPWR systolic_inst.A_shift\[27\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25538_ systolic_inst.acc_wires\[0\]\[14\] C_out\[14\] net54 VGND VGND VPWR VPWR
+ _02840_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13552_ deser_A.shift_reg\[116\] deser_A.shift_reg\[117\] net130 VGND VGND VPWR VPWR
+ _00389_ sky130_fd_sc_hd__mux2_1
XFILLER_201_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28257_ clknet_leaf_97_clk _02055_ VGND VGND VPWR VPWR systolic_inst.B_shift\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16271_ _03652_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__inv_2
X_13483_ deser_A.shift_reg\[47\] deser_A.shift_reg\[48\] net130 VGND VGND VPWR VPWR
+ _00320_ sky130_fd_sc_hd__mux2_1
X_25469_ _11207_ _11208_ systolic_inst.cycle_cnt\[12\] VGND VGND VPWR VPWR _02806_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18010_ _05201_ _05200_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__nand2b_1
XFILLER_240_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15222_ _12323_ _12324_ VGND VGND VPWR VPWR _12325_ sky130_fd_sc_hd__xnor2_1
X_27208_ clknet_leaf_256_clk _01006_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_199_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28188_ clknet_leaf_124_clk _01986_ VGND VGND VPWR VPWR systolic_inst.B_shift\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27139_ clknet_leaf_87_clk _00937_ VGND VGND VPWR VPWR systolic_inst.B_shift\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_15153_ _12265_ VGND VGND VPWR VPWR _12266_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_101_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_126_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14104_ systolic_inst.A_shift\[12\]\[4\] net72 _11333_ A_in\[60\] VGND VGND VPWR
+ VPWR _00926_ sky130_fd_sc_hd__a22o_1
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19961_ _06925_ _06928_ _06926_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__o21ba_1
X_15084_ _12134_ _12138_ _12168_ _12166_ VGND VGND VPWR VPWR _12202_ sky130_fd_sc_hd__o31a_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14035_ deser_B.shift_reg\[69\] deser_B.shift_reg\[70\] net126 VGND VGND VPWR VPWR
+ _00861_ sky130_fd_sc_hd__mux2_1
X_18912_ _06015_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__nand2_1
XFILLER_84_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19892_ _06783_ _06889_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_147_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18843_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[8\]\[7\]
+ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__or2_1
XFILLER_80_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18774_ _05806_ _05895_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__nand2_1
X_15986_ _12978_ _12984_ VGND VGND VPWR VPWR _12986_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_106_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17725_ systolic_inst.acc_wires\[10\]\[20\] systolic_inst.acc_wires\[10\]\[21\] systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__o21a_1
XFILLER_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14937_ _12027_ _12057_ VGND VGND VPWR VPWR _12059_ sky130_fd_sc_hd__xor2_1
XFILLER_57_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_168_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17656_ _04876_ _04883_ _04885_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__o21a_1
X_14868_ _11961_ _11964_ _11966_ VGND VGND VPWR VPWR _11991_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_63_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16607_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.A_outs\[11\]\[1\] systolic_inst.B_outs\[11\]\[2\]
+ systolic_inst.B_outs\[11\]\[3\] VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__and4_1
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13819_ B_in\[126\] deser_B.word_buffer\[126\] net89 VGND VGND VPWR VPWR _00656_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17587_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[10\]\[0\]
+ _04828_ _04826_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__a31o_1
X_14799_ _11918_ _11924_ VGND VGND VPWR VPWR _11925_ sky130_fd_sc_hd__nor2_1
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19326_ _06355_ _06357_ _06385_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__nand3_1
XFILLER_232_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16538_ _03888_ _03889_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19257_ _06317_ _06318_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__xnor2_1
X_16469_ _03829_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__nand2b_1
XFILLER_192_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_340_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_340_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_51_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18208_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[9\]\[3\]
+ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__and2_1
XFILLER_223_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19188_ systolic_inst.A_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[5\] _06216_ _06215_
+ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_136_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18139_ _05326_ _05325_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_132_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21150_ _07976_ _07979_ _08019_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__nand3_1
XFILLER_137_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20101_ _07075_ _07079_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__nand2b_1
XFILLER_99_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21081_ _07915_ _07918_ _07920_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_242_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20032_ _07015_ _07016_ _07014_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__a21bo_1
XFILLER_113_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24840_ net113 ser_C.shift_reg\[248\] VGND VGND VPWR VPWR _10890_ sky130_fd_sc_hd__and2_1
XFILLER_230_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_219_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_159_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_159_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_230_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21983_ net106 systolic_inst.acc_wires\[3\]\[16\] net65 _08767_ VGND VGND VPWR VPWR
+ _01762_ sky130_fd_sc_hd__a22o_1
X_24771_ C_out\[212\] net98 net78 ser_C.shift_reg\[212\] _10855_ VGND VGND VPWR VPWR
+ _02462_ sky130_fd_sc_hd__a221o_1
XFILLER_27_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26510_ clknet_leaf_18_A_in_serial_clk _00313_ net143 VGND VGND VPWR VPWR deser_A.shift_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_23722_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[0\]\[5\]
+ VGND VGND VPWR VPWR _10334_ sky130_fd_sc_hd__nand2_1
X_20934_ _07775_ _07808_ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27490_ clknet_leaf_228_clk _01288_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_199_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26441_ clknet_leaf_348_clk _00248_ net132 VGND VGND VPWR VPWR A_in\[109\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23653_ _10267_ _10271_ VGND VGND VPWR VPWR _10273_ sky130_fd_sc_hd__xor2_1
XFILLER_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20865_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[3\] _07740_ _07741_
+ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__a22o_1
XFILLER_148_1168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22604_ _09318_ _09319_ _09316_ VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__o21ai_1
X_29160_ clknet_leaf_309_clk _02958_ net142 VGND VGND VPWR VPWR C_out\[132\] sky130_fd_sc_hd__dfrtp_1
XFILLER_169_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23584_ _10161_ _10164_ _10204_ VGND VGND VPWR VPWR _10206_ sky130_fd_sc_hd__nor3_1
X_26372_ clknet_leaf_23_clk _00179_ net135 VGND VGND VPWR VPWR A_in\[40\] sky130_fd_sc_hd__dfrtp_1
X_20796_ _07696_ _07698_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28111_ clknet_leaf_57_clk _01909_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22535_ _09255_ _09261_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__nand2_1
XFILLER_210_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25323_ ser_C.parallel_data\[488\] net97 net77 ser_C.shift_reg\[488\] _11131_ VGND
+ VGND VPWR VPWR _02738_ sky130_fd_sc_hd__a221o_1
XFILLER_70_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29091_ clknet_leaf_155_clk _02889_ net150 VGND VGND VPWR VPWR C_out\[63\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_331_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_331_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_194_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28042_ clknet_leaf_164_clk _01840_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22466_ _09196_ _09197_ net106 _09195_ VGND VGND VPWR VPWR _09204_ sky130_fd_sc_hd__a211o_1
XFILLER_196_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25254_ net111 ser_C.shift_reg\[455\] VGND VGND VPWR VPWR _11097_ sky130_fd_sc_hd__and2_1
XFILLER_120_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21417_ _08237_ _08257_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__nor2_1
X_24205_ systolic_inst.A_shift\[21\]\[2\] A_in\[82\] net59 VGND VGND VPWR VPWR _10588_
+ sky130_fd_sc_hd__mux2_1
X_25185_ C_out\[419\] net102 net74 ser_C.shift_reg\[419\] _11062_ VGND VGND VPWR VPWR
+ _02669_ sky130_fd_sc_hd__a221o_1
X_22397_ _09103_ _09105_ _09136_ VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_187_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_208_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24136_ _10569_ systolic_inst.A_shift\[29\]\[7\] net71 VGND VGND VPWR VPWR _02113_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21348_ _08197_ _08198_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__and2_1
XFILLER_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24067_ systolic_inst.B_shift\[19\]\[5\] B_in\[29\] net59 VGND VGND VPWR VPWR _10551_
+ sky130_fd_sc_hd__mux2_1
X_28944_ clknet_leaf_256_clk _02742_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[492\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_204_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21279_ _08138_ _08139_ _08131_ _08135_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_204_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23018_ _09627_ _09693_ VGND VGND VPWR VPWR _09694_ sky130_fd_sc_hd__nand2_1
X_28875_ clknet_leaf_290_clk _02673_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[423\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27826_ clknet_leaf_217_clk _01624_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15840_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[13\]\[12\]
+ _12873_ VGND VGND VPWR VPWR _12877_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_5_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27757_ clknet_leaf_208_clk _01555_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15771_ _12814_ _12815_ _12816_ VGND VGND VPWR VPWR _12818_ sky130_fd_sc_hd__and3_1
XFILLER_218_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24969_ C_out\[311\] net103 net76 ser_C.shift_reg\[311\] _10954_ VGND VGND VPWR VPWR
+ _02561_ sky130_fd_sc_hd__a221o_1
XFILLER_40_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17510_ _04761_ _04762_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__nor2_1
X_26708_ clknet_leaf_10_B_in_serial_clk _00511_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14722_ net69 _11870_ _11871_ systolic_inst.acc_wires\[15\]\[28\] net105 VGND VGND
+ VPWR VPWR _01006_ sky130_fd_sc_hd__a32o_1
XFILLER_218_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18490_ _05579_ _05597_ _05596_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__a21bo_1
X_27688_ clknet_leaf_199_clk _01486_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29427_ clknet_leaf_344_clk _03225_ net131 VGND VGND VPWR VPWR C_out\[399\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17441_ _04693_ _04694_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__xnor2_1
X_26639_ clknet_leaf_13_B_in_serial_clk _00442_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_14653_ systolic_inst.acc_wires\[15\]\[16\] systolic_inst.acc_wires\[15\]\[17\] systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _11813_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_16_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13604_ deser_B.word_buffer\[40\] deser_B.serial_word\[40\] net123 VGND VGND VPWR
+ VPWR _00441_ sky130_fd_sc_hd__mux2_1
XFILLER_220_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17372_ _04628_ _04598_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__nand2b_1
X_29358_ clknet_leaf_231_clk _03156_ net140 VGND VGND VPWR VPWR C_out\[330\] sky130_fd_sc_hd__dfrtp_1
X_14584_ _11753_ _11752_ systolic_inst.acc_wires\[15\]\[8\] net105 VGND VGND VPWR
+ VPWR _00986_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_242_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19111_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[4\] _06176_ _06177_
+ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__nand4_2
X_16323_ _03660_ _03702_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__xor2_1
X_28309_ clknet_leaf_348_clk _02107_ VGND VGND VPWR VPWR systolic_inst.A_shift\[29\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_201_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13535_ deser_A.shift_reg\[99\] deser_A.shift_reg\[100\] net129 VGND VGND VPWR VPWR
+ _00372_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_322_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_322_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29289_ clknet_leaf_324_clk _03087_ net142 VGND VGND VPWR VPWR C_out\[261\] sky130_fd_sc_hd__dfrtp_1
XFILLER_242_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19042_ systolic_inst.A_outs\[7\]\[1\] systolic_inst.B_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[3\]
+ systolic_inst.A_outs\[7\]\[0\] VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__a22oi_1
XFILLER_9_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16254_ _03634_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__nor2_1
X_13466_ deser_A.shift_reg\[30\] deser_A.shift_reg\[31\] deser_A.receiving VGND VGND
+ VPWR VPWR _00303_ sky130_fd_sc_hd__mux2_1
XFILLER_145_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15205_ _12306_ _12308_ VGND VGND VPWR VPWR _12310_ sky130_fd_sc_hd__nand2_1
XFILLER_51_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16185_ _03565_ _03568_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13397_ A_in\[106\] deser_A.word_buffer\[106\] net96 VGND VGND VPWR VPWR _00245_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15136_ _12199_ _12203_ _12226_ _12227_ _12249_ VGND VGND VPWR VPWR _12252_ sky130_fd_sc_hd__o311a_1
XFILLER_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19944_ _06890_ _06940_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__and2b_1
X_15067_ _12184_ _12183_ VGND VGND VPWR VPWR _12185_ sky130_fd_sc_hd__nand2b_1
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14018_ deser_B.shift_reg\[52\] deser_B.shift_reg\[53\] net125 VGND VGND VPWR VPWR
+ _00844_ sky130_fd_sc_hd__mux2_1
XFILLER_141_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19875_ _06871_ _06872_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__xor2_1
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18826_ _05941_ _05942_ _05934_ _05938_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__a211o_1
XFILLER_237_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18757_ _05880_ _05879_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__and2b_1
X_15969_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.B_outs\[7\]\[2\] net119 VGND
+ VGND VPWR VPWR _01148_ sky130_fd_sc_hd__mux2_1
XFILLER_36_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17708_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[20\]
+ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__or2_1
XFILLER_3_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18688_ _05811_ _05812_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17639_ _04876_ _04877_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__and2_1
XFILLER_91_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20650_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[5\]\[5\]
+ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__nand2_1
XFILLER_225_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19309_ _06335_ _06339_ _06367_ _06369_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__o22a_1
X_20581_ _07463_ _07512_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_313_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_313_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_143_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22320_ systolic_inst.B_outs\[2\]\[5\] systolic_inst.A_outs\[2\]\[5\] VGND VGND VPWR
+ VPWR _09063_ sky130_fd_sc_hd__nand2_1
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22251_ systolic_inst.A_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[6\]
+ systolic_inst.B_outs\[2\]\[7\] VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__and4b_1
XFILLER_164_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21202_ _08036_ _08043_ _08068_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__and3_1
XFILLER_118_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22182_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.A_outs\[2\]\[1\] systolic_inst.B_outs\[2\]\[5\]
+ systolic_inst.B_outs\[2\]\[6\] VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__and4_1
XFILLER_65_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21133_ _08001_ _08002_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26990_ clknet_leaf_30_A_in_serial_clk _00788_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_160_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21064_ _07887_ _07895_ _07894_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__a21o_1
XFILLER_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25941_ systolic_inst.acc_wires\[13\]\[1\] C_out\[417\] net27 VGND VGND VPWR VPWR
+ _03243_ sky130_fd_sc_hd__mux2_1
XFILLER_99_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20015_ net119 _07006_ _07007_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__a21oi_1
X_28660_ clknet_leaf_182_clk _02458_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[208\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25872_ systolic_inst.acc_wires\[10\]\[28\] C_out\[348\] net41 VGND VGND VPWR VPWR
+ _03174_ sky130_fd_sc_hd__mux2_1
XFILLER_101_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27611_ clknet_leaf_204_clk _01409_ net146 VGND VGND VPWR VPWR systolic_inst.B_outs\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_98_1118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24823_ C_out\[238\] net99 net79 ser_C.shift_reg\[238\] _10881_ VGND VGND VPWR VPWR
+ _02488_ sky130_fd_sc_hd__a221o_1
XFILLER_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28591_ clknet_leaf_40_clk _02389_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[139\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_228_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27542_ clknet_leaf_34_clk _01340_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_24754_ net113 ser_C.shift_reg\[205\] VGND VGND VPWR VPWR _10847_ sky130_fd_sc_hd__and2_1
X_21966_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[15\]
+ VGND VGND VPWR VPWR _08752_ sky130_fd_sc_hd__or2_1
XFILLER_15_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23705_ _10316_ _10317_ _10318_ VGND VGND VPWR VPWR _10320_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_48_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _07754_ _07791_ _07792_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__and3_1
X_27473_ clknet_leaf_221_clk _01271_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_230_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21897_ net68 _08691_ _08693_ systolic_inst.acc_wires\[3\]\[4\] net106 VGND VGND
+ VPWR VPWR _01750_ sky130_fd_sc_hd__a32o_1
X_24685_ C_out\[169\] net104 net76 ser_C.shift_reg\[169\] _10812_ VGND VGND VPWR VPWR
+ _02419_ sky130_fd_sc_hd__a221o_1
XFILLER_226_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29212_ clknet_leaf_181_clk _03010_ net148 VGND VGND VPWR VPWR C_out\[184\] sky130_fd_sc_hd__dfrtp_1
X_26424_ clknet_leaf_9_clk _00231_ net134 VGND VGND VPWR VPWR A_in\[92\] sky130_fd_sc_hd__dfrtp_1
X_23636_ _10234_ _10236_ _10233_ VGND VGND VPWR VPWR _10256_ sky130_fd_sc_hd__o21a_1
X_20848_ _07727_ _07725_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[1\]
+ net108 VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_202_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29143_ clknet_leaf_165_clk _02941_ net150 VGND VGND VPWR VPWR C_out\[115\] sky130_fd_sc_hd__dfrtp_1
XFILLER_204_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26355_ clknet_leaf_18_clk _00162_ net133 VGND VGND VPWR VPWR A_in\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20779_ systolic_inst.acc_wires\[5\]\[20\] systolic_inst.acc_wires\[5\]\[21\] systolic_inst.acc_wires\[5\]\[22\]
+ systolic_inst.acc_wires\[5\]\[23\] systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__o41a_1
X_23567_ _10185_ _10188_ VGND VGND VPWR VPWR _10189_ sky130_fd_sc_hd__and2b_1
XFILLER_70_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_304_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_304_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_189_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_189_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_189_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ A_in\[29\] deser_A.word_buffer\[29\] net91 VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__mux2_1
X_25306_ net111 ser_C.shift_reg\[481\] VGND VGND VPWR VPWR _11123_ sky130_fd_sc_hd__and2_1
X_22518_ net65 _09246_ _09247_ systolic_inst.acc_wires\[2\]\[7\] net109 VGND VGND
+ VPWR VPWR _01817_ sky130_fd_sc_hd__a32o_1
X_29074_ clknet_leaf_113_clk _02872_ net152 VGND VGND VPWR VPWR C_out\[46\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23498_ _11266_ systolic_inst.B_outs\[0\]\[7\] _10120_ VGND VGND VPWR VPWR _10122_
+ sky130_fd_sc_hd__and3_1
XFILLER_122_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26286_ clknet_leaf_26_A_in_serial_clk _00094_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28025_ clknet_leaf_161_clk _01823_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22449_ _09125_ _09187_ VGND VGND VPWR VPWR _09188_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25237_ ser_C.parallel_data\[445\] net102 net74 ser_C.shift_reg\[445\] _11088_ VGND
+ VGND VPWR VPWR _02695_ sky130_fd_sc_hd__a221o_1
X_13251_ deser_A.word_buffer\[89\] deser_A.serial_word\[89\] net127 VGND VGND VPWR
+ VPWR _00099_ sky130_fd_sc_hd__mux2_1
X_13182_ deser_A.word_buffer\[20\] deser_A.serial_word\[20\] net128 VGND VGND VPWR
+ VPWR _00030_ sky130_fd_sc_hd__mux2_1
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25168_ net110 ser_C.shift_reg\[412\] VGND VGND VPWR VPWR _11054_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_107_Left_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24119_ systolic_inst.B_shift\[27\]\[6\] net72 _11333_ B_in\[126\] VGND VGND VPWR
+ VPWR _02104_ sky130_fd_sc_hd__a22o_1
XFILLER_237_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25099_ C_out\[376\] net98 net78 ser_C.shift_reg\[376\] _11019_ VGND VGND VPWR VPWR
+ _02626_ sky130_fd_sc_hd__a221o_1
X_17990_ _05141_ _05144_ _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_144_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28927_ clknet_leaf_266_clk _02725_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[475\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_96_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16941_ _04253_ _04254_ _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19660_ systolic_inst.A_outs\[6\]\[1\] systolic_inst.B_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\]
+ systolic_inst.A_outs\[6\]\[0\] VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__a22o_1
XFILLER_49_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28858_ clknet_leaf_335_clk _02656_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[406\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16872_ _04189_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__inv_2
X_18611_ _05735_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__xnor2_1
X_27809_ clknet_leaf_139_clk _01607_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_15823_ _12860_ _12861_ VGND VGND VPWR VPWR _12862_ sky130_fd_sc_hd__nand2_1
X_19591_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[28\]
+ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__nand2_1
XFILLER_133_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28789_ clknet_leaf_212_clk _02587_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_237_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18542_ systolic_inst.A_outs\[8\]\[1\] systolic_inst.B_outs\[8\]\[6\] _05671_ VGND
+ VGND VPWR VPWR _05672_ sky130_fd_sc_hd__and3_1
X_15754_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[13\]\[1\]
+ VGND VGND VPWR VPWR _12803_ sky130_fd_sc_hd__nand2_1
XFILLER_73_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14705_ _11855_ _11856_ VGND VGND VPWR VPWR _11857_ sky130_fd_sc_hd__nand2_1
XFILLER_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18473_ _05601_ _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__xor2_1
X_15685_ _12738_ VGND VGND VPWR VPWR _12739_ sky130_fd_sc_hd__inv_2
XFILLER_221_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17424_ systolic_inst.B_outs\[10\]\[5\] systolic_inst.A_outs\[10\]\[5\] VGND VGND
+ VPWR VPWR _04679_ sky130_fd_sc_hd__nand2_1
XFILLER_178_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _11798_ _11797_ systolic_inst.acc_wires\[15\]\[15\] net105 VGND VGND VPWR
+ VPWR _00993_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_99_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ systolic_inst.A_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[5\] VGND VGND
+ VPWR VPWR _04612_ sky130_fd_sc_hd__nand2_1
X_14567_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[15\]\[6\]
+ VGND VGND VPWR VPWR _11739_ sky130_fd_sc_hd__nand2_1
XFILLER_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_894 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16306_ _03684_ _03685_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__and2_1
XFILLER_186_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13518_ deser_A.shift_reg\[82\] deser_A.shift_reg\[83\] net129 VGND VGND VPWR VPWR
+ _00355_ sky130_fd_sc_hd__mux2_1
XFILLER_174_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17286_ _04542_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__nor2_1
XFILLER_201_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14498_ _11273_ systolic_inst.A_outs\[15\]\[7\] _11626_ _11650_ VGND VGND VPWR VPWR
+ _11678_ sky130_fd_sc_hd__o211a_1
Xclkload303 clknet_leaf_187_clk VGND VGND VPWR VPWR clkload303/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_58_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19025_ systolic_inst.B_outs\[6\]\[6\] systolic_inst.B_outs\[2\]\[6\] net120 VGND
+ VGND VPWR VPWR _01472_ sky130_fd_sc_hd__mux2_1
Xclkload314 clknet_leaf_109_clk VGND VGND VPWR VPWR clkload314/Y sky130_fd_sc_hd__clkinv_4
X_16237_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__inv_2
Xclkload11 clknet_5_12__leaf_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_6
Xclkload325 clknet_leaf_149_clk VGND VGND VPWR VPWR clkload325/Y sky130_fd_sc_hd__inv_6
Xclkload22 clknet_5_27__leaf_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__clkinvlp_4
X_13449_ deser_A.shift_reg\[13\] deser_A.shift_reg\[14\] deser_A.receiving VGND VGND
+ VPWR VPWR _00286_ sky130_fd_sc_hd__mux2_1
Xclkload336 clknet_leaf_164_clk VGND VGND VPWR VPWR clkload336/Y sky130_fd_sc_hd__clkinv_4
XFILLER_220_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload33 clknet_leaf_340_clk VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__inv_8
XFILLER_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload44 clknet_leaf_289_clk VGND VGND VPWR VPWR clkload44/X sky130_fd_sc_hd__clkbuf_4
Xclkload347 clknet_leaf_22_A_in_serial_clk VGND VGND VPWR VPWR clkload347/Y sky130_fd_sc_hd__inv_8
XFILLER_161_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload55 clknet_leaf_315_clk VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__inv_6
Xclkload358 clknet_leaf_10_A_in_serial_clk VGND VGND VPWR VPWR clkload358/Y sky130_fd_sc_hd__inv_6
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload369 clknet_leaf_0_B_in_serial_clk VGND VGND VPWR VPWR clkload369/Y sky130_fd_sc_hd__bufinv_16
XFILLER_142_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16168_ _03508_ _03511_ _03550_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__or3_1
Xclkload66 clknet_leaf_9_clk VGND VGND VPWR VPWR clkload66/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_90_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload77 clknet_leaf_14_clk VGND VGND VPWR VPWR clkload77/X sky130_fd_sc_hd__clkbuf_8
Xclkload88 clknet_leaf_311_clk VGND VGND VPWR VPWR clkload88/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_90_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload99 clknet_leaf_307_clk VGND VGND VPWR VPWR clkload99/Y sky130_fd_sc_hd__inv_6
XFILLER_216_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15119_ _12146_ _12234_ VGND VGND VPWR VPWR _12235_ sky130_fd_sc_hd__nor2_1
XFILLER_114_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16099_ _13057_ _13093_ VGND VGND VPWR VPWR _13094_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19927_ _06923_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__inv_2
XFILLER_190_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19858_ systolic_inst.B_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[6\] systolic_inst.A_outs\[6\]\[7\]
+ systolic_inst.B_outs\[6\]\[3\] VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__a22o_1
XFILLER_151_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18809_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[8\]\[2\]
+ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__and2_1
XFILLER_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19789_ _06788_ _06789_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__nor2_1
XFILLER_95_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21820_ _08556_ _08622_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__or2_1
XFILLER_3_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21751_ systolic_inst.B_outs\[3\]\[5\] systolic_inst.A_outs\[3\]\[6\] VGND VGND VPWR
+ VPWR _08557_ sky130_fd_sc_hd__nand2_1
XFILLER_93_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_233_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_233_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_233_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20702_ _07615_ _07616_ _07617_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24470_ net114 ser_C.shift_reg\[63\] VGND VGND VPWR VPWR _10705_ sky130_fd_sc_hd__and2_1
XFILLER_197_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21682_ systolic_inst.A_outs\[3\]\[4\] systolic_inst.B_outs\[3\]\[5\] VGND VGND VPWR
+ VPWR _08490_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_43_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23421_ _10038_ _10046_ VGND VGND VPWR VPWR _10047_ sky130_fd_sc_hd__nand2_1
X_20633_ _07556_ _07557_ _07558_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__and3_1
X_26140_ deser_B.serial_word\[95\] deser_B.shift_reg\[95\] net56 VGND VGND VPWR VPWR
+ _03442_ sky130_fd_sc_hd__mux2_1
X_23352_ _09950_ _09952_ VGND VGND VPWR VPWR _09980_ sky130_fd_sc_hd__nand2_1
Xclkload5 clknet_5_6__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_12
X_20564_ _07494_ _07495_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22303_ _09010_ _09012_ _09046_ VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__nand3_1
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26071_ deser_B.serial_word\[26\] deser_B.shift_reg\[26\] net56 VGND VGND VPWR VPWR
+ _03373_ sky130_fd_sc_hd__mux2_1
X_23283_ systolic_inst.A_outs\[0\]\[6\] systolic_inst.A_shift\[0\]\[6\] net121 VGND
+ VGND VPWR VPWR _01912_ sky130_fd_sc_hd__mux2_1
X_20495_ systolic_inst.A_outs\[5\]\[6\] _07398_ _07399_ _07364_ VGND VGND VPWR VPWR
+ _07429_ sky130_fd_sc_hd__o2bb2a_1
X_22234_ _08978_ _08979_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__xor2_1
X_25022_ net112 ser_C.shift_reg\[339\] VGND VGND VPWR VPWR _10981_ sky130_fd_sc_hd__and2_1
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_30__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_30__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_180_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22165_ _08911_ _08912_ VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__nand2_1
XFILLER_160_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21116_ _07983_ _07985_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22096_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.A_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\]
+ systolic_inst.A_outs\[2\]\[1\] VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__and4_1
X_26973_ clknet_leaf_24_A_in_serial_clk _00771_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28712_ clknet_leaf_325_clk _02510_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[260\]
+ sky130_fd_sc_hd__dfrtp_1
X_21047_ _07914_ _07918_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__xnor2_1
X_25924_ systolic_inst.acc_wires\[12\]\[16\] C_out\[400\] net18 VGND VGND VPWR VPWR
+ _03226_ sky130_fd_sc_hd__mux2_1
X_29692_ clknet_leaf_346_clk _03487_ VGND VGND VPWR VPWR systolic_inst.A_shift\[30\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28643_ clknet_leaf_182_clk _02441_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25855_ systolic_inst.acc_wires\[10\]\[11\] C_out\[331\] net12 VGND VGND VPWR VPWR
+ _03157_ sky130_fd_sc_hd__mux2_1
XFILLER_101_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24806_ net113 ser_C.shift_reg\[231\] VGND VGND VPWR VPWR _10873_ sky130_fd_sc_hd__and2_1
XFILLER_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_A_in_serial_clk A_in_serial_clk VGND VGND VPWR VPWR clknet_0_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
X_28574_ clknet_leaf_174_clk _02372_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_25786_ systolic_inst.acc_wires\[8\]\[6\] C_out\[262\] net22 VGND VGND VPWR VPWR
+ _03088_ sky130_fd_sc_hd__mux2_1
X_22998_ _09622_ _09674_ VGND VGND VPWR VPWR _09675_ sky130_fd_sc_hd__and2b_1
XFILLER_90_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27525_ clknet_leaf_233_clk _01323_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24737_ C_out\[195\] net97 net80 ser_C.shift_reg\[195\] _10838_ VGND VGND VPWR VPWR
+ _02445_ sky130_fd_sc_hd__a221o_1
XFILLER_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21949_ _08736_ _08737_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_81_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_199_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15470_ _12527_ _12528_ _12497_ VGND VGND VPWR VPWR _12530_ sky130_fd_sc_hd__a21oi_1
XFILLER_76_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27456_ clknet_leaf_239_clk _01254_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24668_ net110 ser_C.shift_reg\[162\] VGND VGND VPWR VPWR _10804_ sky130_fd_sc_hd__and2_1
XFILLER_202_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14421_ _11602_ _11603_ VGND VGND VPWR VPWR _11604_ sky130_fd_sc_hd__nand2_1
X_26407_ clknet_leaf_30_clk _00214_ net133 VGND VGND VPWR VPWR A_in\[75\] sky130_fd_sc_hd__dfrtp_1
X_23619_ _10238_ _10239_ VGND VGND VPWR VPWR _10240_ sky130_fd_sc_hd__nand2_1
X_27387_ clknet_leaf_338_clk _01185_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_24599_ C_out\[126\] net99 net80 ser_C.shift_reg\[126\] _10769_ VGND VGND VPWR VPWR
+ _02376_ sky130_fd_sc_hd__a221o_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29126_ clknet_leaf_178_clk _02924_ net148 VGND VGND VPWR VPWR C_out\[98\] sky130_fd_sc_hd__dfrtp_1
XFILLER_156_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17140_ _04422_ _04424_ _04426_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__o21ai_1
X_26338_ clknet_leaf_58_clk _00145_ net137 VGND VGND VPWR VPWR A_in\[6\] sky130_fd_sc_hd__dfrtp_1
X_14352_ _11527_ _11536_ VGND VGND VPWR VPWR _11537_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1003 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13303_ A_in\[12\] deser_A.word_buffer\[12\] net93 VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__mux2_1
X_29057_ clknet_leaf_109_clk _02855_ net151 VGND VGND VPWR VPWR C_out\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17071_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[15\]
+ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__nor2_1
XFILLER_144_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14283_ _11435_ _11468_ VGND VGND VPWR VPWR _11470_ sky130_fd_sc_hd__nor2_1
X_26269_ clknet_leaf_21_A_in_serial_clk _00077_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_171_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28008_ clknet_leaf_149_clk _01806_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_16022_ _13019_ VGND VGND VPWR VPWR _13020_ sky130_fd_sc_hd__inv_2
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13234_ deser_A.word_buffer\[72\] deser_A.serial_word\[72\] net127 VGND VGND VPWR
+ VPWR _00082_ sky130_fd_sc_hd__mux2_1
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13165_ deser_A.word_buffer\[3\] deser_A.serial_word\[3\] net128 VGND VGND VPWR VPWR
+ _00013_ sky130_fd_sc_hd__mux2_1
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17973_ _05165_ _05164_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_163_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_163_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19712_ _06713_ _06714_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__nor2_1
X_16924_ _04238_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__nand2b_1
XFILLER_242_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19643_ net119 _06647_ _06648_ _06649_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__a31o_1
XFILLER_133_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16855_ _04171_ _04172_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__or2_1
XFILLER_225_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15806_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[13\]\[9\]
+ VGND VGND VPWR VPWR _12847_ sky130_fd_sc_hd__xor2_1
XFILLER_81_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19574_ _06600_ _06602_ _06604_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_122_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16786_ _04102_ _04105_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__xnor2_1
XFILLER_225_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13998_ deser_B.shift_reg\[32\] deser_B.shift_reg\[33\] net125 VGND VGND VPWR VPWR
+ _00824_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18525_ _05625_ _05648_ _05647_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__a21boi_1
X_15737_ _12786_ _12787_ VGND VGND VPWR VPWR _12789_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_55_1308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18456_ _05569_ _05586_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__and3_1
XFILLER_221_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15668_ _12719_ _12720_ VGND VGND VPWR VPWR _12722_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_17407_ _04660_ _04661_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14619_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[15\]\[12\]
+ _11780_ VGND VGND VPWR VPWR _11784_ sky130_fd_sc_hd__and3_1
X_18387_ _05542_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__inv_2
X_15599_ _12651_ _12654_ VGND VGND VPWR VPWR _12655_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17338_ _04558_ _04559_ _04556_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__o21ai_1
XFILLER_105_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload100 clknet_leaf_308_clk VGND VGND VPWR VPWR clkload100/Y sky130_fd_sc_hd__clkinv_8
XFILLER_105_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload111 clknet_leaf_286_clk VGND VGND VPWR VPWR clkload111/Y sky130_fd_sc_hd__clkinv_4
X_17269_ _04502_ _04528_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__xor2_1
XFILLER_162_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload122 clknet_leaf_295_clk VGND VGND VPWR VPWR clkload122/Y sky130_fd_sc_hd__bufinv_16
XFILLER_220_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload133 clknet_leaf_272_clk VGND VGND VPWR VPWR clkload133/Y sky130_fd_sc_hd__clkinvlp_4
X_19008_ _06092_ _06096_ _06097_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_77_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload144 clknet_leaf_221_clk VGND VGND VPWR VPWR clkload144/X sky130_fd_sc_hd__clkbuf_4
Xclkload155 clknet_leaf_211_clk VGND VGND VPWR VPWR clkload155/Y sky130_fd_sc_hd__inv_8
X_20280_ _07199_ _07217_ _07218_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_77_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload166 clknet_leaf_230_clk VGND VGND VPWR VPWR clkload166/X sky130_fd_sc_hd__clkbuf_8
Xclkload177 clknet_leaf_200_clk VGND VGND VPWR VPWR clkload177/Y sky130_fd_sc_hd__inv_4
Xclkload188 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload188/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_226_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload199 clknet_leaf_67_clk VGND VGND VPWR VPWR clkload199/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_226_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23970_ _10510_ systolic_inst.B_shift\[9\]\[4\] _11332_ VGND VGND VPWR VPWR _02006_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_239_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22921_ _09597_ _09598_ VGND VGND VPWR VPWR _09600_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_235_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_235_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_235_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25640_ systolic_inst.acc_wires\[3\]\[20\] C_out\[116\] net50 VGND VGND VPWR VPWR
+ _02942_ sky130_fd_sc_hd__mux2_1
X_22852_ systolic_inst.B_outs\[1\]\[7\] _09530_ _09531_ VGND VGND VPWR VPWR _09533_
+ sky130_fd_sc_hd__and3_1
XFILLER_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21803_ _08605_ _08606_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__and2_1
XFILLER_227_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25571_ systolic_inst.acc_wires\[1\]\[15\] C_out\[47\] net35 VGND VGND VPWR VPWR
+ _02873_ sky130_fd_sc_hd__mux2_1
X_22783_ _09435_ _09464_ _09465_ VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__nand3_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_63_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27310_ clknet_leaf_300_clk _01108_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24522_ net114 ser_C.shift_reg\[89\] VGND VGND VPWR VPWR _10731_ sky130_fd_sc_hd__and2_1
XFILLER_227_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21734_ _08482_ _08539_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__or2_1
X_28290_ clknet_leaf_75_clk _02088_ VGND VGND VPWR VPWR systolic_inst.B_shift\[19\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27241_ clknet_leaf_279_clk _01039_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24453_ C_out\[53\] _11302_ net81 ser_C.shift_reg\[53\] _10696_ VGND VGND VPWR VPWR
+ _02303_ sky130_fd_sc_hd__a221o_1
XFILLER_185_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21665_ _08471_ _08472_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__and2_1
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23404_ _10024_ _10029_ VGND VGND VPWR VPWR _10030_ sky130_fd_sc_hd__or2_1
XFILLER_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20616_ _07542_ _07545_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__xnor2_1
X_27172_ clknet_leaf_254_clk _00970_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24384_ net7 ser_C.shift_reg\[20\] VGND VGND VPWR VPWR _10662_ sky130_fd_sc_hd__and2_1
X_21596_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[6\]
+ systolic_inst.A_outs\[3\]\[7\] VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__nand4_1
XFILLER_197_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26123_ deser_B.serial_word\[78\] deser_B.shift_reg\[78\] net55 VGND VGND VPWR VPWR
+ _03425_ sky130_fd_sc_hd__mux2_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23335_ _09963_ VGND VGND VPWR VPWR _09964_ sky130_fd_sc_hd__inv_2
X_20547_ _07432_ _07448_ _07446_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__o21a_1
XFILLER_197_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26054_ deser_B.serial_word\[9\] deser_B.shift_reg\[9\] net55 VGND VGND VPWR VPWR
+ _03356_ sky130_fd_sc_hd__mux2_1
X_23266_ _09899_ _09902_ _09905_ _09908_ VGND VGND VPWR VPWR _09909_ sky130_fd_sc_hd__o31a_1
X_20478_ _07411_ _07412_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__nand2b_1
XFILLER_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25005_ C_out\[329\] net97 net80 ser_C.shift_reg\[329\] _10972_ VGND VGND VPWR VPWR
+ _02579_ sky130_fd_sc_hd__a221o_1
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22217_ _08928_ _08961_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23197_ _09846_ _09848_ _09845_ VGND VGND VPWR VPWR _09851_ sky130_fd_sc_hd__o21ai_1
XFILLER_193_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22148_ _08892_ _08895_ VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__xor2_1
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22079_ systolic_inst.A_outs\[2\]\[1\] systolic_inst.A_outs\[1\]\[1\] net122 VGND
+ VGND VPWR VPWR _01779_ sky130_fd_sc_hd__mux2_1
XFILLER_120_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14970_ _12089_ _12090_ VGND VGND VPWR VPWR _12091_ sky130_fd_sc_hd__nand2_1
XFILLER_48_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26956_ clknet_leaf_2_A_in_serial_clk _00754_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25907_ systolic_inst.acc_wires\[11\]\[31\] C_out\[383\] net11 VGND VGND VPWR VPWR
+ _03209_ sky130_fd_sc_hd__mux2_1
XFILLER_75_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13921_ deser_A.serial_word\[82\] deser_A.shift_reg\[82\] net57 VGND VGND VPWR VPWR
+ _00747_ sky130_fd_sc_hd__mux2_1
X_29675_ clknet_leaf_31_B_in_serial_clk _03470_ net134 VGND VGND VPWR VPWR deser_B.serial_word\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_26887_ clknet_leaf_8_A_in_serial_clk _00685_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28626_ clknet_leaf_146_clk _02424_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[174\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16640_ _03944_ _03946_ _03945_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a21bo_1
X_25838_ systolic_inst.acc_wires\[9\]\[26\] C_out\[314\] net13 VGND VGND VPWR VPWR
+ _03140_ sky130_fd_sc_hd__mux2_1
X_13852_ deser_A.serial_word\[13\] deser_A.shift_reg\[13\] net58 VGND VGND VPWR VPWR
+ _00678_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28557_ clknet_leaf_169_clk _02355_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16571_ _03912_ _03914_ _03913_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__a21bo_1
X_25769_ systolic_inst.acc_wires\[7\]\[21\] C_out\[245\] net44 VGND VGND VPWR VPWR
+ _03071_ sky130_fd_sc_hd__mux2_1
X_13783_ B_in\[90\] deser_B.word_buffer\[90\] net89 VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_54_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18310_ _05476_ _05477_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__xnor2_1
XFILLER_163_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15522_ _12575_ _12578_ VGND VGND VPWR VPWR _12580_ sky130_fd_sc_hd__xnor2_1
X_27508_ clknet_leaf_230_clk _01306_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_19290_ _06350_ _06351_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__or2_1
X_28488_ clknet_leaf_113_clk _02286_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_231_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18241_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[9\]\[8\]
+ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_239_Left_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15453_ _12508_ _12511_ VGND VGND VPWR VPWR _12513_ sky130_fd_sc_hd__xnor2_1
X_27439_ clknet_leaf_245_clk _01237_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14404_ systolic_inst.A_outs\[15\]\[6\] _11558_ _11559_ _11447_ VGND VGND VPWR VPWR
+ _11587_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18172_ _05358_ _05357_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__and2b_1
X_15384_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[2\] _12447_ VGND
+ VGND VPWR VPWR _12448_ sky130_fd_sc_hd__nand3_1
X_29109_ clknet_leaf_160_clk _02907_ net150 VGND VGND VPWR VPWR C_out\[81\] sky130_fd_sc_hd__dfrtp_1
X_17123_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[23\]
+ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__xor2_1
XFILLER_15_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14335_ _11515_ _11519_ VGND VGND VPWR VPWR _11520_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17054_ net105 systolic_inst.acc_wires\[11\]\[12\] net69 _04354_ VGND VGND VPWR VPWR
+ _01246_ sky130_fd_sc_hd__a22o_1
XFILLER_176_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14266_ systolic_inst.A_outs\[15\]\[0\] systolic_inst.B_outs\[15\]\[7\] VGND VGND
+ VPWR VPWR _11453_ sky130_fd_sc_hd__and2b_1
XFILLER_109_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16005_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[3\] _13003_ net115
+ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13217_ deser_A.word_buffer\[55\] deser_A.serial_word\[55\] net128 VGND VGND VPWR
+ VPWR _00065_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14197_ systolic_inst.A_outs\[15\]\[0\] systolic_inst.B_outs\[15\]\[5\] VGND VGND
+ VPWR VPWR _11386_ sky130_fd_sc_hd__and2_1
XFILLER_83_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ ser_C.bit_idx\[1\] ser_C.bit_idx\[2\] _11299_ VGND VGND VPWR VPWR _11300_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_72_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17956_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[7\]
+ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__o21a_1
XFILLER_239_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16907_ _04223_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__inv_2
XFILLER_238_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17887_ _05080_ _05081_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__nor2_1
XFILLER_239_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19626_ systolic_inst.B_outs\[5\]\[6\] systolic_inst.B_outs\[1\]\[6\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__mux2_1
XFILLER_54_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16838_ _04155_ _04156_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__or2_1
XFILLER_4_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19557_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[23\]
+ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__xor2_1
X_16769_ _04087_ _04088_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_45_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_20_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18508_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.A_outs\[8\]\[1\] systolic_inst.B_outs\[8\]\[5\]
+ systolic_inst.B_outs\[8\]\[6\] VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__and4_1
X_19488_ net60 _06532_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__nor2_1
XFILLER_178_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18439_ _05562_ _05571_ _05572_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__nand3_1
XFILLER_181_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21450_ _08283_ _08285_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_25_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20401_ systolic_inst.A_outs\[5\]\[0\] _07267_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_228_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21381_ net63 _08226_ _08227_ systolic_inst.acc_wires\[4\]\[18\] _11258_ VGND VGND
+ VPWR VPWR _01700_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_21_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23120_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[1\]\[8\]
+ VGND VGND VPWR VPWR _09785_ sky130_fd_sc_hd__xor2_1
X_20332_ _07265_ _07266_ _07269_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_224_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23051_ _09723_ _09724_ VGND VGND VPWR VPWR _09726_ sky130_fd_sc_hd__and2b_1
XFILLER_116_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20263_ _07198_ _07203_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22002_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[20\]
+ VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__nand2_1
XFILLER_192_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_1_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_20194_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[27\]
+ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26810_ clknet_leaf_76_clk _00612_ net144 VGND VGND VPWR VPWR B_in\[82\] sky130_fd_sc_hd__dfrtp_1
X_27790_ clknet_leaf_40_clk _01588_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_26741_ clknet_leaf_98_clk _00543_ net153 VGND VGND VPWR VPWR B_in\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23953_ systolic_inst.B_shift\[11\]\[0\] net70 net83 systolic_inst.B_shift\[15\]\[0\]
+ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__a22o_1
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22904_ _09582_ _09583_ VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__xnor2_1
X_29460_ clknet_leaf_330_clk _03258_ net136 VGND VGND VPWR VPWR C_out\[432\] sky130_fd_sc_hd__dfrtp_1
X_26672_ clknet_leaf_9_B_in_serial_clk _00475_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23884_ systolic_inst.acc_wires\[0\]\[28\] systolic_inst.acc_wires\[0\]\[29\] systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _10471_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28411_ clknet_leaf_83_clk _02209_ VGND VGND VPWR VPWR systolic_inst.B_shift\[17\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_186_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25623_ systolic_inst.acc_wires\[3\]\[3\] C_out\[99\] net48 VGND VGND VPWR VPWR _02925_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22835_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[7\]
+ VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__o21a_1
X_29391_ clknet_leaf_241_clk _03189_ net145 VGND VGND VPWR VPWR C_out\[363\] sky130_fd_sc_hd__dfrtp_1
XFILLER_112_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_36_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28342_ clknet_leaf_342_clk _02140_ VGND VGND VPWR VPWR systolic_inst.A_shift\[25\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25554_ systolic_inst.acc_wires\[0\]\[30\] C_out\[30\] net36 VGND VGND VPWR VPWR
+ _02856_ sky130_fd_sc_hd__mux2_1
XFILLER_198_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22766_ _09430_ _09432_ _09431_ VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__o21bai_1
XFILLER_13_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24505_ C_out\[79\] net100 net80 ser_C.shift_reg\[79\] _10722_ VGND VGND VPWR VPWR
+ _02329_ sky130_fd_sc_hd__a221o_1
XFILLER_213_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21717_ systolic_inst.A_outs\[3\]\[4\] systolic_inst.B_outs\[3\]\[6\] _11274_ systolic_inst.A_outs\[3\]\[3\]
+ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__o2bb2a_1
X_28273_ clknet_leaf_130_clk _02071_ VGND VGND VPWR VPWR systolic_inst.B_shift\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_25485_ _11220_ VGND VGND VPWR VPWR _11221_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_213_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22697_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[1\]
+ systolic_inst.A_outs\[1\]\[2\] VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__and4_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27224_ clknet_leaf_291_clk _01022_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_24436_ net114 ser_C.shift_reg\[46\] VGND VGND VPWR VPWR _10688_ sky130_fd_sc_hd__and2_1
X_21648_ _08453_ _08456_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27155_ clknet_leaf_294_clk _00953_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_24367_ C_out\[10\] net104 _10643_ ser_C.shift_reg\[10\] _10653_ VGND VGND VPWR VPWR
+ _02260_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_151_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21579_ _08385_ _08386_ _08388_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__or3_1
X_26106_ deser_B.serial_word\[61\] deser_B.shift_reg\[61\] net56 VGND VGND VPWR VPWR
+ _03408_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14120_ systolic_inst.A_shift\[21\]\[4\] net71 _11333_ A_in\[92\] VGND VGND VPWR
+ VPWR _00942_ sky130_fd_sc_hd__a22o_1
X_23318_ _09929_ _09946_ VGND VGND VPWR VPWR _09947_ sky130_fd_sc_hd__or2_1
X_27086_ clknet_leaf_32_B_in_serial_clk _00884_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24298_ _10622_ systolic_inst.A_shift\[11\]\[4\] net71 VGND VGND VPWR VPWR _02222_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14051_ deser_B.shift_reg\[85\] deser_B.shift_reg\[86\] net125 VGND VGND VPWR VPWR
+ _00877_ sky130_fd_sc_hd__mux2_1
X_26037_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[11\]\[1\] net118 VGND
+ VGND VPWR VPWR _03339_ sky130_fd_sc_hd__mux2_1
X_23249_ _09888_ _09892_ _09889_ VGND VGND VPWR VPWR _09895_ sky130_fd_sc_hd__a21bo_1
XFILLER_101_1383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17810_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[1\]
+ systolic_inst.A_outs\[9\]\[2\] VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__and4_1
X_18790_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[14\] _05912_ net117
+ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__mux2_1
X_27988_ clknet_leaf_121_clk _01786_ net152 VGND VGND VPWR VPWR systolic_inst.B_outs\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_94_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17741_ _04964_ _04965_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__or2_1
X_14953_ _12072_ _12073_ VGND VGND VPWR VPWR _12074_ sky130_fd_sc_hd__or2_1
X_26939_ clknet_leaf_20_A_in_serial_clk _00737_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13904_ deser_A.serial_word\[65\] deser_A.shift_reg\[65\] net57 VGND VGND VPWR VPWR
+ _00730_ sky130_fd_sc_hd__mux2_1
X_17672_ _04904_ _04905_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__nand2_1
X_29658_ clknet_leaf_7_B_in_serial_clk _03453_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14884_ systolic_inst.A_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[7\] VGND VGND
+ VPWR VPWR _12007_ sky130_fd_sc_hd__and2b_1
XFILLER_78_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19411_ net69 _06465_ _06466_ systolic_inst.acc_wires\[7\]\[1\] net105 VGND VGND
+ VPWR VPWR _01491_ sky130_fd_sc_hd__a32o_1
XFILLER_75_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16623_ _03944_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13835_ _11321_ _11326_ _11328_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__and3_1
X_28609_ clknet_leaf_134_clk _02407_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[157\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29589_ clknet_leaf_12_B_in_serial_clk _03384_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap60 _11713_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_12
XFILLER_51_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_104_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap82 _10643_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_12
X_19342_ _06401_ _06402_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__nor2_1
X_16554_ systolic_inst.acc_wires\[12\]\[26\] systolic_inst.acc_wires\[12\]\[27\] systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__o21a_1
XFILLER_91_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13766_ B_in\[73\] deser_B.word_buffer\[73\] net90 VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__mux2_1
Xmax_cap93 net95 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_8
XFILLER_31_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15505_ _12525_ _12527_ VGND VGND VPWR VPWR _12564_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_100_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19273_ _06333_ _06334_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16485_ _03841_ _03844_ net67 VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__o21ai_1
X_13697_ B_in\[4\] deser_B.word_buffer\[4\] net86 VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__mux2_1
XFILLER_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18224_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[9\]\[5\]
+ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__or2_1
XFILLER_31_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15436_ _12488_ _12496_ VGND VGND VPWR VPWR _12497_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18155_ _05341_ _05342_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__nor2_1
XFILLER_200_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15367_ systolic_inst.B_outs\[12\]\[3\] systolic_inst.B_outs\[8\]\[3\] net115 VGND
+ VGND VPWR VPWR _01085_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17106_ systolic_inst.acc_wires\[11\]\[16\] systolic_inst.acc_wires\[11\]\[17\] systolic_inst.acc_wires\[11\]\[18\]
+ systolic_inst.acc_wires\[11\]\[19\] systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__o41a_1
XFILLER_184_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14318_ _11501_ _11502_ VGND VGND VPWR VPWR _11504_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_74_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18086_ _05259_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__xor2_1
X_15298_ _12388_ _12389_ _12387_ VGND VGND VPWR VPWR _12390_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_74_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17037_ _04337_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__xor2_1
XFILLER_176_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14249_ _11381_ _11409_ _11408_ VGND VGND VPWR VPWR _11436_ sky130_fd_sc_hd__a21o_1
XFILLER_217_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18988_ _06065_ _06067_ _06079_ _06080_ _06073_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__a311oi_4
XFILLER_79_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_183_Right_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17939_ _05096_ _05131_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__and2_1
XFILLER_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20950_ _07801_ _07824_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__nor2_1
XFILLER_26_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19609_ _06629_ _06633_ _06634_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_217_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_217_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20881_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[3\] VGND VGND VPWR
+ VPWR _07758_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_18_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_187_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22620_ _09326_ _09330_ _09332_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__a21oi_1
XFILLER_228_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22551_ _09272_ _09273_ _09274_ VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21502_ _08304_ _08314_ _08315_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__nand3_1
X_25270_ net111 ser_C.shift_reg\[463\] VGND VGND VPWR VPWR _11105_ sky130_fd_sc_hd__and2_1
XFILLER_33_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22482_ _09213_ _09214_ _09215_ VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__and3_1
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24221_ systolic_inst.A_shift\[20\]\[2\] A_in\[74\] net59 VGND VGND VPWR VPWR _10596_
+ sky130_fd_sc_hd__mux2_1
X_21433_ _08269_ _08271_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21364_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[16\]
+ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__nand2_1
X_24152_ _10577_ systolic_inst.A_shift\[28\]\[7\] net71 VGND VGND VPWR VPWR _02121_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23103_ _09767_ _09768_ _09769_ VGND VGND VPWR VPWR _09771_ sky130_fd_sc_hd__and3_1
X_20315_ systolic_inst.A_outs\[5\]\[4\] _07215_ _07232_ _07231_ _07228_ VGND VGND
+ VPWR VPWR _07254_ sky130_fd_sc_hd__a32o_1
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24083_ systolic_inst.B_shift\[2\]\[2\] _11332_ net83 systolic_inst.B_shift\[6\]\[2\]
+ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__a22o_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28960_ clknet_leaf_257_clk _02758_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[508\]
+ sky130_fd_sc_hd__dfrtp_1
X_21295_ _08153_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__inv_2
XFILLER_235_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23034_ _09679_ _09684_ _09709_ VGND VGND VPWR VPWR _09710_ sky130_fd_sc_hd__or3_1
X_27911_ clknet_leaf_44_clk _01709_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_122_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20246_ systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[2\]
+ systolic_inst.B_outs\[5\]\[0\] VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_57_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28891_ clknet_leaf_287_clk _02689_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[439\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27842_ clknet_leaf_205_clk _01640_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_104_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_206_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20177_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[24\]
+ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__and2_1
XFILLER_104_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27773_ clknet_leaf_186_clk _01571_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_44_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_202_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24985_ C_out\[319\] net97 net80 ser_C.shift_reg\[319\] _10962_ VGND VGND VPWR VPWR
+ _02569_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_202_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_198_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26724_ clknet_leaf_33_B_in_serial_clk _00527_ net134 VGND VGND VPWR VPWR deser_B.word_buffer\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_29512_ clknet_leaf_261_clk _03310_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[484\]
+ sky130_fd_sc_hd__dfrtp_1
X_23936_ systolic_inst.B_shift\[14\]\[0\] B_in\[16\] _00008_ VGND VGND VPWR VPWR _10497_
+ sky130_fd_sc_hd__mux2_1
XFILLER_229_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29443_ clknet_leaf_333_clk _03241_ net131 VGND VGND VPWR VPWR C_out\[415\] sky130_fd_sc_hd__dfrtp_1
XFILLER_217_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26655_ clknet_leaf_24_B_in_serial_clk _00458_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23867_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[27\]
+ VGND VGND VPWR VPWR _10457_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_194_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25606_ systolic_inst.acc_wires\[2\]\[18\] C_out\[82\] net52 VGND VGND VPWR VPWR
+ _02908_ sky130_fd_sc_hd__mux2_1
X_13620_ deser_B.word_buffer\[56\] deser_B.serial_word\[56\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__mux2_1
XFILLER_72_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22818_ _09487_ _09499_ VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__or2_1
X_29374_ clknet_leaf_236_clk _03172_ net145 VGND VGND VPWR VPWR C_out\[346\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26586_ clknet_leaf_30_A_in_serial_clk _00389_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_23798_ _10384_ _10390_ _10398_ VGND VGND VPWR VPWR _10399_ sky130_fd_sc_hd__a21o_1
XFILLER_73_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28325_ clknet_leaf_3_clk _02123_ VGND VGND VPWR VPWR systolic_inst.A_shift\[27\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_213_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25537_ systolic_inst.acc_wires\[0\]\[13\] C_out\[13\] net33 VGND VGND VPWR VPWR
+ _02839_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13551_ deser_A.shift_reg\[115\] deser_A.shift_reg\[116\] net129 VGND VGND VPWR VPWR
+ _00388_ sky130_fd_sc_hd__mux2_1
X_22749_ _09430_ _09431_ _09432_ VGND VGND VPWR VPWR _09433_ sky130_fd_sc_hd__or3_1
XFILLER_41_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28256_ clknet_leaf_79_clk _02054_ VGND VGND VPWR VPWR systolic_inst.B_shift\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16270_ _03613_ _03615_ _03650_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__a21oi_1
X_25468_ _11208_ _11209_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13482_ deser_A.shift_reg\[46\] deser_A.shift_reg\[47\] net130 VGND VGND VPWR VPWR
+ _00319_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15221_ _12316_ _12318_ _12314_ VGND VGND VPWR VPWR _12324_ sky130_fd_sc_hd__a21bo_1
X_27207_ clknet_leaf_258_clk _01005_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_24419_ C_out\[36\] _11302_ net81 ser_C.shift_reg\[36\] _10679_ VGND VGND VPWR VPWR
+ _02286_ sky130_fd_sc_hd__a221o_1
XFILLER_240_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28187_ clknet_leaf_19_clk _01985_ VGND VGND VPWR VPWR systolic_inst.A_shift\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25399_ systolic_inst.A_shift\[3\]\[7\] A_in\[23\] net59 VGND VGND VPWR VPWR _11169_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27138_ clknet_leaf_87_clk _00936_ VGND VGND VPWR VPWR systolic_inst.B_shift\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_15152_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[14\]\[0\]
+ _12263_ _12264_ VGND VGND VPWR VPWR _12265_ sky130_fd_sc_hd__and4_1
XFILLER_153_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14103_ systolic_inst.A_shift\[12\]\[3\] net72 _11333_ A_in\[59\] VGND VGND VPWR
+ VPWR _00925_ sky130_fd_sc_hd__a22o_1
XFILLER_154_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27069_ clknet_leaf_9_B_in_serial_clk _00867_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_19960_ _06928_ _06955_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15083_ _12199_ _12200_ VGND VGND VPWR VPWR _12201_ sky130_fd_sc_hd__nor2_1
XFILLER_101_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14034_ deser_B.shift_reg\[68\] deser_B.shift_reg\[69\] net126 VGND VGND VPWR VPWR
+ _00860_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18911_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[16\]
+ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__nand2_1
X_19891_ systolic_inst.A_outs\[6\]\[6\] _06858_ _06859_ _06825_ VGND VGND VPWR VPWR
+ _06889_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_147_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18842_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[8\]\[7\]
+ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__nand2_1
XFILLER_121_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15985_ _12984_ VGND VGND VPWR VPWR _12985_ sky130_fd_sc_hd__inv_2
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18773_ _05806_ _05895_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__or2_1
XFILLER_83_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14936_ _12057_ _12027_ VGND VGND VPWR VPWR _12058_ sky130_fd_sc_hd__nand2b_1
X_17724_ _04949_ _04950_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__and2_1
XFILLER_63_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14867_ _11951_ _11981_ _11983_ VGND VGND VPWR VPWR _11990_ sky130_fd_sc_hd__o21ba_1
X_17655_ _04867_ _04891_ _04879_ _04889_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13818_ B_in\[125\] deser_B.word_buffer\[125\] net89 VGND VGND VPWR VPWR _00655_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16606_ systolic_inst.A_outs\[11\]\[1\] systolic_inst.B_outs\[11\]\[2\] systolic_inst.B_outs\[11\]\[3\]
+ systolic_inst.A_outs\[11\]\[0\] VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a22oi_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17586_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[10\]\[2\]
+ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__or2_1
XFILLER_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14798_ _11903_ _11922_ VGND VGND VPWR VPWR _11924_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19325_ _06355_ _06357_ _06385_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__a21o_1
X_16537_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[24\]
+ _03886_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a21oi_1
X_13749_ B_in\[56\] deser_B.word_buffer\[56\] net85 VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__mux2_1
XFILLER_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19256_ _06318_ _06317_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__nand2b_1
X_16468_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[15\]
+ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__nand2_1
XFILLER_108_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15419_ net107 _12479_ _12480_ VGND VGND VPWR VPWR _12481_ sky130_fd_sc_hd__or3_1
X_18207_ net66 _05387_ _05389_ systolic_inst.acc_wires\[9\]\[2\] net107 VGND VGND
+ VPWR VPWR _01364_ sky130_fd_sc_hd__a32o_1
X_19187_ _06248_ _06251_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_136_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16399_ _03768_ _03770_ _03763_ _03766_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__a211o_1
XFILLER_185_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18138_ _05293_ _05296_ _05294_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_97_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18069_ _05257_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__nand2_1
XFILLER_105_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20100_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[6\]\[12\]
+ _07077_ _07079_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_93_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21080_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[9\] _07951_ net117
+ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_99_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_242_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_242_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20031_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[6\]\[3\]
+ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__or2_1
XFILLER_8_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24770_ net113 ser_C.shift_reg\[213\] VGND VGND VPWR VPWR _10855_ sky130_fd_sc_hd__and2_1
XFILLER_227_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21982_ _08764_ _08765_ VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23721_ net63 _10331_ _10333_ systolic_inst.acc_wires\[0\]\[4\] _11258_ VGND VGND
+ VPWR VPWR _01934_ sky130_fd_sc_hd__a32o_1
XFILLER_27_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20933_ _07802_ _07806_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26440_ clknet_leaf_348_clk _00247_ net132 VGND VGND VPWR VPWR A_in\[108\] sky130_fd_sc_hd__dfrtp_1
X_23652_ _10267_ _10271_ VGND VGND VPWR VPWR _10272_ sky130_fd_sc_hd__and2b_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20864_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[3\] _07740_ _07741_
+ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__nand4_1
XFILLER_183_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22603_ _09316_ _09318_ _09319_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__or3_1
XFILLER_168_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26371_ clknet_leaf_26_clk _00178_ net143 VGND VGND VPWR VPWR A_in\[39\] sky130_fd_sc_hd__dfrtp_1
X_23583_ _10161_ _10164_ _10204_ VGND VGND VPWR VPWR _10205_ sky130_fd_sc_hd__o21a_1
XFILLER_23_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20795_ _07689_ _07691_ _07697_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__a21o_1
XFILLER_169_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28110_ clknet_leaf_57_clk _01908_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_224_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25322_ net112 ser_C.shift_reg\[489\] VGND VGND VPWR VPWR _11131_ sky130_fd_sc_hd__and2_1
X_29090_ clknet_leaf_156_clk _02888_ net150 VGND VGND VPWR VPWR C_out\[62\] sky130_fd_sc_hd__dfrtp_1
X_22534_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[2\]\[9\]
+ _09256_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28041_ clknet_leaf_162_clk _01839_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_25253_ ser_C.parallel_data\[453\] net102 net74 ser_C.shift_reg\[453\] _11096_ VGND
+ VGND VPWR VPWR _02703_ sky130_fd_sc_hd__a221o_1
X_22465_ _09199_ _09202_ VGND VGND VPWR VPWR _09203_ sky130_fd_sc_hd__xnor2_1
XFILLER_194_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24204_ _10587_ systolic_inst.A_shift\[20\]\[1\] net71 VGND VGND VPWR VPWR _02163_
+ sky130_fd_sc_hd__mux2_1
X_21416_ systolic_inst.acc_wires\[4\]\[20\] systolic_inst.acc_wires\[4\]\[21\] systolic_inst.acc_wires\[4\]\[22\]
+ systolic_inst.acc_wires\[4\]\[23\] systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__o41a_1
XFILLER_120_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25184_ net111 ser_C.shift_reg\[420\] VGND VGND VPWR VPWR _11062_ sky130_fd_sc_hd__and2_1
X_22396_ _09103_ _09105_ _09136_ VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_187_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24135_ systolic_inst.A_shift\[30\]\[7\] A_in\[119\] net59 VGND VGND VPWR VPWR _10569_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21347_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[4\]\[14\]
+ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__nand2_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_208_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24066_ _10550_ systolic_inst.B_shift\[15\]\[4\] net70 VGND VGND VPWR VPWR _02062_
+ sky130_fd_sc_hd__mux2_1
X_28943_ clknet_leaf_256_clk _02741_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[491\]
+ sky130_fd_sc_hd__dfrtp_1
X_21278_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[4\]\[4\]
+ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_204_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23017_ _09691_ _09692_ VGND VGND VPWR VPWR _09693_ sky130_fd_sc_hd__and2_1
X_20229_ systolic_inst.A_outs\[5\]\[6\] systolic_inst.A_outs\[4\]\[6\] net117 VGND
+ VGND VPWR VPWR _01592_ sky130_fd_sc_hd__mux2_1
XFILLER_238_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28874_ clknet_leaf_279_clk _02672_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[422\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27825_ clknet_leaf_217_clk _01623_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15770_ _12814_ _12815_ _12816_ VGND VGND VPWR VPWR _12817_ sky130_fd_sc_hd__a21o_1
X_27756_ clknet_leaf_208_clk _01554_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24968_ net111 ser_C.shift_reg\[312\] VGND VGND VPWR VPWR _10954_ sky130_fd_sc_hd__and2_1
XFILLER_218_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14721_ _11866_ _11869_ VGND VGND VPWR VPWR _11871_ sky130_fd_sc_hd__nand2_1
X_26707_ clknet_leaf_10_B_in_serial_clk _00510_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_23919_ _10492_ systolic_inst.B_shift\[18\]\[3\] net71 VGND VGND VPWR VPWR _01973_
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27687_ clknet_leaf_199_clk _01485_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24899_ C_out\[276\] net103 net75 ser_C.shift_reg\[276\] _10919_ VGND VGND VPWR VPWR
+ _02526_ sky130_fd_sc_hd__a221o_1
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17440_ _04694_ _04693_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__nand2b_1
X_26638_ clknet_leaf_13_B_in_serial_clk _00441_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_14652_ _11810_ _11811_ VGND VGND VPWR VPWR _11812_ sky130_fd_sc_hd__nand2_1
X_29426_ clknet_leaf_344_clk _03224_ net131 VGND VGND VPWR VPWR C_out\[398\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ deser_B.word_buffer\[39\] deser_B.serial_word\[39\] net123 VGND VGND VPWR
+ VPWR _00440_ sky130_fd_sc_hd__mux2_1
XFILLER_60_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17371_ _04625_ _04626_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__xor2_1
XFILLER_232_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26569_ clknet_leaf_23_A_in_serial_clk _00372_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_14583_ _11750_ _11751_ net69 VGND VGND VPWR VPWR _11753_ sky130_fd_sc_hd__o21ai_1
X_29357_ clknet_leaf_230_clk _03155_ net140 VGND VGND VPWR VPWR C_out\[329\] sky130_fd_sc_hd__dfrtp_1
XFILLER_158_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19110_ systolic_inst.B_outs\[7\]\[3\] systolic_inst.A_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\]
+ systolic_inst.A_outs\[7\]\[2\] VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__a22o_1
X_16322_ _03699_ _03700_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__xor2_1
XFILLER_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13534_ deser_A.shift_reg\[98\] deser_A.shift_reg\[99\] net129 VGND VGND VPWR VPWR
+ _00371_ sky130_fd_sc_hd__mux2_1
X_28308_ clknet_leaf_8_clk _02106_ VGND VGND VPWR VPWR systolic_inst.A_shift\[29\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_29288_ clknet_leaf_324_clk _03086_ net142 VGND VGND VPWR VPWR C_out\[260\] sky130_fd_sc_hd__dfrtp_1
XFILLER_199_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19041_ net119 _06110_ _06111_ _06104_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__a31o_1
X_28239_ clknet_leaf_130_clk _02037_ VGND VGND VPWR VPWR systolic_inst.B_shift\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16253_ systolic_inst.A_outs\[12\]\[5\] systolic_inst.B_outs\[12\]\[6\] _11260_ systolic_inst.A_outs\[12\]\[4\]
+ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_185_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13465_ deser_A.shift_reg\[29\] deser_A.shift_reg\[30\] deser_A.receiving VGND VGND
+ VPWR VPWR _00302_ sky130_fd_sc_hd__mux2_1
XFILLER_16_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15204_ _12303_ _12306_ _12308_ _12305_ VGND VGND VPWR VPWR _12309_ sky130_fd_sc_hd__a211o_1
X_16184_ _03566_ _03567_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__nor2_1
XFILLER_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13396_ A_in\[105\] deser_A.word_buffer\[105\] net95 VGND VGND VPWR VPWR _00244_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15135_ _12249_ _12250_ VGND VGND VPWR VPWR _12251_ sky130_fd_sc_hd__or2_1
XFILLER_103_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_189_Left_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19943_ _06937_ _06938_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__xnor2_1
X_15066_ _12147_ _12149_ _12148_ VGND VGND VPWR VPWR _12184_ sky130_fd_sc_hd__o21ba_1
XFILLER_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14017_ deser_B.shift_reg\[51\] deser_B.shift_reg\[52\] net125 VGND VGND VPWR VPWR
+ _00843_ sky130_fd_sc_hd__mux2_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19874_ _06871_ _06872_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__nand2b_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18825_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[8\]\[4\]
+ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__or2_1
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18756_ _05835_ _05847_ _05845_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__o21a_1
X_15968_ systolic_inst.B_outs\[11\]\[1\] systolic_inst.B_outs\[7\]\[1\] net119 VGND
+ VGND VPWR VPWR _01147_ sky130_fd_sc_hd__mux2_1
XFILLER_114_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17707_ net106 systolic_inst.acc_wires\[10\]\[19\] _11712_ _04936_ VGND VGND VPWR
+ VPWR _01317_ sky130_fd_sc_hd__a22o_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14919_ systolic_inst.A_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[5\] VGND VGND
+ VPWR VPWR _12041_ sky130_fd_sc_hd__nand2_1
X_15899_ systolic_inst.acc_wires\[13\]\[20\] systolic_inst.acc_wires\[13\]\[21\] systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12927_ sky130_fd_sc_hd__o21a_1
X_18687_ _05812_ _05811_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_198_Left_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17638_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[10\]\[10\]
+ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__or2_1
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17569_ _04742_ _04804_ _04802_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19308_ _06335_ _06339_ _06367_ _06369_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__nor4_1
X_20580_ _07510_ _07511_ VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__nor2_1
XFILLER_108_1153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19239_ _06299_ _06300_ _06301_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22250_ systolic_inst.A_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[5\] VGND VGND VPWR
+ VPWR _08995_ sky130_fd_sc_hd__nand2_1
XFILLER_180_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21201_ _08036_ _08043_ _08068_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__a21oi_1
X_22181_ systolic_inst.A_outs\[2\]\[1\] systolic_inst.B_outs\[2\]\[6\] VGND VGND VPWR
+ VPWR _08928_ sky130_fd_sc_hd__nand2_1
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21132_ systolic_inst.A_outs\[4\]\[4\] _07852_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21063_ _07926_ _07934_ VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__xnor2_1
X_25940_ systolic_inst.acc_wires\[13\]\[0\] C_out\[416\] net27 VGND VGND VPWR VPWR
+ _03242_ sky130_fd_sc_hd__mux2_1
XFILLER_232_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20014_ net119 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[6\]\[0\]
+ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25871_ systolic_inst.acc_wires\[10\]\[27\] C_out\[347\] net11 VGND VGND VPWR VPWR
+ _03173_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27610_ clknet_leaf_204_clk _01408_ net146 VGND VGND VPWR VPWR systolic_inst.B_outs\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_24822_ net113 ser_C.shift_reg\[239\] VGND VGND VPWR VPWR _10881_ sky130_fd_sc_hd__and2_1
X_28590_ clknet_leaf_40_clk _02388_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[138\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27541_ clknet_leaf_34_clk _01339_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_24753_ C_out\[203\] net99 net79 ser_C.shift_reg\[203\] _10846_ VGND VGND VPWR VPWR
+ _02453_ sky130_fd_sc_hd__a221o_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21965_ net68 _08750_ _08751_ systolic_inst.acc_wires\[3\]\[14\] net106 VGND VGND
+ VPWR VPWR _01760_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_191_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _10316_ _10317_ _10318_ VGND VGND VPWR VPWR _10319_ sky130_fd_sc_hd__a21o_1
XFILLER_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27472_ clknet_leaf_222_clk _01270_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_20916_ _07788_ _07789_ _07790_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__a21o_1
X_24684_ net112 ser_C.shift_reg\[170\] VGND VGND VPWR VPWR _10812_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21896_ _08692_ VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__inv_2
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29211_ clknet_leaf_181_clk _03009_ net148 VGND VGND VPWR VPWR C_out\[183\] sky130_fd_sc_hd__dfrtp_1
X_26423_ clknet_leaf_13_clk _00230_ net134 VGND VGND VPWR VPWR A_in\[91\] sky130_fd_sc_hd__dfrtp_1
X_23635_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[12\] _10255_ systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__mux2_1
XFILLER_39_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20847_ net117 _07726_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__nand2_1
XFILLER_168_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29142_ clknet_leaf_166_clk _02940_ net150 VGND VGND VPWR VPWR C_out\[114\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_202_Left_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26354_ clknet_leaf_19_clk _00161_ net133 VGND VGND VPWR VPWR A_in\[22\] sky130_fd_sc_hd__dfrtp_1
X_23566_ _10186_ _10187_ VGND VGND VPWR VPWR _10188_ sky130_fd_sc_hd__nor2_1
XFILLER_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20778_ _07639_ _07640_ _07662_ _07682_ VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_189_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25305_ ser_C.parallel_data\[479\] net102 net74 ser_C.shift_reg\[479\] _11122_ VGND
+ VGND VPWR VPWR _02729_ sky130_fd_sc_hd__a221o_1
X_22517_ _09243_ _09244_ _09245_ VGND VGND VPWR VPWR _09247_ sky130_fd_sc_hd__nand3_1
X_29073_ clknet_leaf_116_clk _02871_ net152 VGND VGND VPWR VPWR C_out\[45\] sky130_fd_sc_hd__dfrtp_1
XFILLER_126_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26285_ clknet_leaf_26_A_in_serial_clk _00093_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_23497_ _11266_ systolic_inst.B_outs\[0\]\[7\] _10120_ VGND VGND VPWR VPWR _10121_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_11_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28024_ clknet_leaf_167_clk _01822_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_202_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25236_ net111 ser_C.shift_reg\[446\] VGND VGND VPWR VPWR _11088_ sky130_fd_sc_hd__and2_1
XFILLER_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13250_ deser_A.word_buffer\[88\] deser_A.serial_word\[88\] net127 VGND VGND VPWR
+ VPWR _00098_ sky130_fd_sc_hd__mux2_1
XFILLER_202_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22448_ _09185_ _09186_ VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__nor2_1
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13181_ deser_A.word_buffer\[19\] deser_A.serial_word\[19\] net128 VGND VGND VPWR
+ VPWR _00029_ sky130_fd_sc_hd__mux2_1
X_25167_ C_out\[410\] net101 net73 ser_C.shift_reg\[410\] _11053_ VGND VGND VPWR VPWR
+ _02660_ sky130_fd_sc_hd__a221o_1
X_22379_ net122 _09120_ VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__nand2_1
XFILLER_191_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24118_ systolic_inst.B_shift\[27\]\[5\] net72 _11333_ B_in\[125\] VGND VGND VPWR
+ VPWR _02103_ sky130_fd_sc_hd__a22o_1
X_25098_ net113 ser_C.shift_reg\[377\] VGND VGND VPWR VPWR _11019_ sky130_fd_sc_hd__and2_1
XFILLER_123_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_211_Left_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24049_ systolic_inst.B_shift\[4\]\[4\] B_in\[4\] _00008_ VGND VGND VPWR VPWR _10542_
+ sky130_fd_sc_hd__mux2_1
X_28926_ clknet_leaf_267_clk _02724_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[474\]
+ sky130_fd_sc_hd__dfrtp_1
X_16940_ _11262_ systolic_inst.A_outs\[11\]\[7\] _04204_ _04227_ VGND VGND VPWR VPWR
+ _04255_ sky130_fd_sc_hd__o211a_1
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28857_ clknet_leaf_335_clk _02655_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[405\]
+ sky130_fd_sc_hd__dfrtp_1
X_16871_ _04150_ _04152_ _04188_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nand3_1
XFILLER_49_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18610_ _05736_ _05737_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_240_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_240_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_219_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27808_ clknet_leaf_217_clk _01606_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_15822_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[13\]\[11\]
+ VGND VGND VPWR VPWR _12861_ sky130_fd_sc_hd__nand2_1
X_19590_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[28\]
+ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__or2_1
XFILLER_213_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28788_ clknet_leaf_225_clk _02586_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[336\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15753_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[13\]\[1\]
+ VGND VGND VPWR VPWR _12802_ sky130_fd_sc_hd__and2_1
X_18541_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[7\] VGND VGND VPWR
+ VPWR _05671_ sky130_fd_sc_hd__and2b_1
XFILLER_92_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27739_ clknet_leaf_132_clk _01537_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_166_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14704_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[26\]
+ VGND VGND VPWR VPWR _11856_ sky130_fd_sc_hd__nand2_1
XFILLER_79_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15684_ _12736_ _12737_ VGND VGND VPWR VPWR _12738_ sky130_fd_sc_hd__or2_1
X_18472_ _05602_ _05603_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__nor2_1
XFILLER_61_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_220_Left_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29409_ clknet_leaf_237_clk _03207_ net147 VGND VGND VPWR VPWR C_out\[381\] sky130_fd_sc_hd__dfrtp_1
X_14635_ _11787_ _11792_ _11796_ net61 VGND VGND VPWR VPWR _11798_ sky130_fd_sc_hd__a31o_1
X_17423_ _04643_ _04677_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_174_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14566_ net69 _11736_ _11738_ systolic_inst.acc_wires\[15\]\[5\] net107 VGND VGND
+ VPWR VPWR _00983_ sky130_fd_sc_hd__a32o_1
X_17354_ _04609_ _04610_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16305_ _03620_ _03624_ _03653_ _03684_ _03651_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__a311oi_4
X_13517_ deser_A.shift_reg\[81\] deser_A.shift_reg\[82\] net129 VGND VGND VPWR VPWR
+ _00354_ sky130_fd_sc_hd__mux2_1
X_17285_ systolic_inst.A_outs\[10\]\[0\] systolic_inst.A_outs\[10\]\[1\] systolic_inst.B_outs\[10\]\[5\]
+ systolic_inst.B_outs\[10\]\[6\] VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__and4_1
XFILLER_144_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14497_ systolic_inst.B_outs\[15\]\[5\] systolic_inst.B_outs\[15\]\[6\] systolic_inst.A_outs\[15\]\[7\]
+ VGND VGND VPWR VPWR _11677_ sky130_fd_sc_hd__nand3_1
XFILLER_186_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload304 clknet_leaf_205_clk VGND VGND VPWR VPWR clkload304/Y sky130_fd_sc_hd__inv_8
X_19024_ systolic_inst.B_outs\[6\]\[5\] systolic_inst.B_outs\[2\]\[5\] net120 VGND
+ VGND VPWR VPWR _01471_ sky130_fd_sc_hd__mux2_1
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16236_ _03617_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_58_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload315 clknet_leaf_110_clk VGND VGND VPWR VPWR clkload315/Y sky130_fd_sc_hd__clkinvlp_4
X_13448_ deser_A.shift_reg\[12\] deser_A.shift_reg\[13\] deser_A.receiving VGND VGND
+ VPWR VPWR _00285_ sky130_fd_sc_hd__mux2_1
XFILLER_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload12 clknet_5_14__leaf_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_8
Xclkload326 clknet_leaf_167_clk VGND VGND VPWR VPWR clkload326/Y sky130_fd_sc_hd__bufinv_16
Xclkload23 clknet_5_28__leaf_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__inv_8
Xclkload337 clknet_leaf_166_clk VGND VGND VPWR VPWR clkload337/Y sky130_fd_sc_hd__bufinv_16
Xclkload34 clknet_leaf_344_clk VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__clkinv_4
XFILLER_220_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload348 clknet_leaf_23_A_in_serial_clk VGND VGND VPWR VPWR clkload348/X sky130_fd_sc_hd__clkbuf_4
Xclkload45 clknet_leaf_326_clk VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__bufinv_16
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16167_ _03508_ _03511_ _03550_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__o21ai_1
Xclkload56 clknet_leaf_318_clk VGND VGND VPWR VPWR clkload56/Y sky130_fd_sc_hd__inv_12
Xclkload359 clknet_leaf_11_A_in_serial_clk VGND VGND VPWR VPWR clkload359/X sky130_fd_sc_hd__clkbuf_8
Xclkload67 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload67/Y sky130_fd_sc_hd__clkinv_8
X_13379_ A_in\[88\] deser_A.word_buffer\[88\] net95 VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__mux2_1
XFILLER_126_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload78 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload78/Y sky130_fd_sc_hd__inv_6
XFILLER_142_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15118_ _12231_ _12232_ _12233_ VGND VGND VPWR VPWR _12234_ sky130_fd_sc_hd__a21oi_1
Xclkload89 clknet_leaf_312_clk VGND VGND VPWR VPWR clkload89/X sky130_fd_sc_hd__clkbuf_8
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16098_ _13091_ _13092_ VGND VGND VPWR VPWR _13093_ sky130_fd_sc_hd__nor2_1
XFILLER_173_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19926_ _06921_ _06922_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__nand2_1
X_15049_ _12128_ _12130_ _12165_ VGND VGND VPWR VPWR _12168_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19857_ _06854_ _06855_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_231_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_231_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18808_ net63 _05926_ _05927_ systolic_inst.acc_wires\[8\]\[1\] net108 VGND VGND
+ VPWR VPWR _01427_ sky130_fd_sc_hd__a32o_1
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19788_ systolic_inst.B_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[5\]
+ systolic_inst.B_outs\[6\]\[3\] VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_88_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18739_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[12\] _05863_ net117
+ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__mux2_1
XFILLER_97_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_237_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1095 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21750_ _08485_ _08555_ VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__xnor2_4
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_233_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_233_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20701_ _07615_ _07616_ _07617_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__and3_1
XFILLER_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21681_ _08485_ _08488_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23420_ _10045_ VGND VGND VPWR VPWR _10046_ sky130_fd_sc_hd__inv_2
X_20632_ _07556_ _07557_ _07558_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_43_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_298_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_298_clk
+ sky130_fd_sc_hd__clkbuf_8
X_23351_ _09973_ _09978_ VGND VGND VPWR VPWR _09979_ sky130_fd_sc_hd__xnor2_1
X_20563_ systolic_inst.A_outs\[5\]\[6\] _11276_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__nor2_1
Xclkload6 clknet_5_7__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_6
XFILLER_165_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22302_ _09020_ _09045_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26070_ deser_B.serial_word\[25\] deser_B.shift_reg\[25\] net56 VGND VGND VPWR VPWR
+ _03372_ sky130_fd_sc_hd__mux2_1
XFILLER_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23282_ systolic_inst.A_outs\[0\]\[5\] systolic_inst.A_shift\[0\]\[5\] net121 VGND
+ VGND VPWR VPWR _01911_ sky130_fd_sc_hd__mux2_1
X_20494_ _07428_ _07426_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[10\]
+ net109 VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25021_ C_out\[337\] net97 net80 ser_C.shift_reg\[337\] _10980_ VGND VGND VPWR VPWR
+ _02587_ sky130_fd_sc_hd__a221o_1
X_22233_ _08911_ _08912_ _08943_ _08941_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__a31o_1
XFILLER_117_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_180_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22164_ _08870_ _08887_ _08886_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__a21bo_1
XFILLER_133_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21115_ _07907_ _07910_ _07946_ _07948_ _07984_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__o311a_1
XFILLER_182_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22095_ net109 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[0\] _08847_
+ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__a21o_1
X_26972_ clknet_leaf_25_A_in_serial_clk _00770_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28711_ clknet_leaf_325_clk _02509_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[259\]
+ sky130_fd_sc_hd__dfrtp_1
X_21046_ _07876_ _07916_ _07917_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__a21o_1
X_25923_ systolic_inst.acc_wires\[12\]\[15\] C_out\[399\] net18 VGND VGND VPWR VPWR
+ _03225_ sky130_fd_sc_hd__mux2_1
X_29691_ clknet_leaf_347_clk _03486_ VGND VGND VPWR VPWR systolic_inst.A_shift\[30\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_219_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_222_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_222_clk
+ sky130_fd_sc_hd__clkbuf_8
X_28642_ clknet_leaf_181_clk _02440_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[190\]
+ sky130_fd_sc_hd__dfrtp_1
X_25854_ systolic_inst.acc_wires\[10\]\[10\] C_out\[330\] net12 VGND VGND VPWR VPWR
+ _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_178_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24805_ C_out\[229\] net99 net79 ser_C.shift_reg\[229\] _10872_ VGND VGND VPWR VPWR
+ _02479_ sky130_fd_sc_hd__a221o_1
X_28573_ clknet_leaf_174_clk _02371_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25785_ systolic_inst.acc_wires\[8\]\[5\] C_out\[261\] net22 VGND VGND VPWR VPWR
+ _03087_ sky130_fd_sc_hd__mux2_1
X_22997_ _09672_ _09673_ VGND VGND VPWR VPWR _09674_ sky130_fd_sc_hd__nor2_1
XFILLER_55_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_886 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24736_ net112 ser_C.shift_reg\[196\] VGND VGND VPWR VPWR _10838_ sky130_fd_sc_hd__and2_1
X_27524_ clknet_leaf_233_clk _01322_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21948_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[3\]\[12\]
+ VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__nand2_1
XFILLER_15_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27455_ clknet_leaf_239_clk _01253_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_24667_ C_out\[160\] net103 net76 ser_C.shift_reg\[160\] _10803_ VGND VGND VPWR VPWR
+ _02410_ sky130_fd_sc_hd__a221o_1
X_21879_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[3\]\[2\]
+ VGND VGND VPWR VPWR _08678_ sky130_fd_sc_hd__or2_1
XFILLER_128_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14420_ _11593_ _11601_ VGND VGND VPWR VPWR _11603_ sky130_fd_sc_hd__or2_1
X_26406_ clknet_leaf_29_clk _00213_ net133 VGND VGND VPWR VPWR A_in\[74\] sky130_fd_sc_hd__dfrtp_1
X_23618_ _10201_ _10203_ _10237_ VGND VGND VPWR VPWR _10239_ sky130_fd_sc_hd__or3_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27386_ clknet_leaf_344_clk _01184_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24598_ net113 ser_C.shift_reg\[127\] VGND VGND VPWR VPWR _10769_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_289_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_289_clk
+ sky130_fd_sc_hd__clkbuf_8
X_29125_ clknet_leaf_178_clk _02923_ net148 VGND VGND VPWR VPWR C_out\[97\] sky130_fd_sc_hd__dfrtp_1
X_26337_ clknet_leaf_25_clk _00144_ net137 VGND VGND VPWR VPWR A_in\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14351_ _11533_ _11534_ VGND VGND VPWR VPWR _11536_ sky130_fd_sc_hd__xor2_1
X_23549_ _10130_ _10132_ _10171_ VGND VGND VPWR VPWR _10172_ sky130_fd_sc_hd__o21a_1
XFILLER_126_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13302_ A_in\[11\] deser_A.word_buffer\[11\] net93 VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__mux2_1
X_29056_ clknet_leaf_110_clk _02854_ net151 VGND VGND VPWR VPWR C_out\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_195_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17070_ net69 _04367_ _04368_ systolic_inst.acc_wires\[11\]\[14\] net105 VGND VGND
+ VPWR VPWR _01248_ sky130_fd_sc_hd__a32o_1
XFILLER_196_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14282_ _11435_ _11468_ VGND VGND VPWR VPWR _11469_ sky130_fd_sc_hd__and2_1
X_26268_ clknet_leaf_16_A_in_serial_clk _00076_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_1253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16021_ _12996_ _12999_ _13018_ VGND VGND VPWR VPWR _13019_ sky130_fd_sc_hd__a21o_1
X_28007_ clknet_5_30__leaf_clk _01805_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_25219_ C_out\[436\] net101 net73 ser_C.shift_reg\[436\] _11079_ VGND VGND VPWR VPWR
+ _02686_ sky130_fd_sc_hd__a221o_1
X_13233_ deser_A.word_buffer\[71\] deser_A.serial_word\[71\] net127 VGND VGND VPWR
+ VPWR _00081_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26199_ systolic_inst.A_shift\[30\]\[5\] net71 _11333_ A_in\[125\] VGND VGND VPWR
+ VPWR _03489_ sky130_fd_sc_hd__a22o_1
XFILLER_87_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13164_ deser_A.word_buffer\[2\] deser_A.serial_word\[2\] net128 VGND VGND VPWR VPWR
+ _00012_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17972_ systolic_inst.A_outs\[9\]\[2\] systolic_inst.B_outs\[9\]\[5\] _05127_ _05126_
+ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__a31oi_2
XFILLER_105_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19711_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[5\]
+ systolic_inst.A_outs\[6\]\[6\] VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__and4_1
X_28909_ clknet_leaf_281_clk _02707_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16923_ _04169_ _04208_ _04207_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a21bo_1
XFILLER_172_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_213_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_213_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19642_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _06649_ sky130_fd_sc_hd__and2_1
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16854_ systolic_inst.A_outs\[11\]\[5\] systolic_inst.B_outs\[11\]\[6\] _11262_ systolic_inst.A_outs\[11\]\[4\]
+ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15805_ _12846_ _12845_ systolic_inst.acc_wires\[13\]\[8\] net107 VGND VGND VPWR
+ VPWR _01114_ sky130_fd_sc_hd__a2bb2o_1
X_19573_ _06600_ _06602_ _06604_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__or3_1
XFILLER_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13997_ deser_B.shift_reg\[31\] deser_B.shift_reg\[32\] net125 VGND VGND VPWR VPWR
+ _00823_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16785_ _04103_ _04104_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__nor2_1
XFILLER_207_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18524_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[6\] _05654_ net115
+ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__mux2_1
XFILLER_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15736_ _12787_ _12786_ VGND VGND VPWR VPWR _12788_ sky130_fd_sc_hd__nand2b_1
XFILLER_34_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18455_ systolic_inst.A_outs\[8\]\[4\] _05587_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__nand2_1
X_15667_ systolic_inst.B_outs\[13\]\[5\] systolic_inst.A_outs\[13\]\[7\] _12719_ VGND
+ VGND VPWR VPWR _12721_ sky130_fd_sc_hd__and3_1
XFILLER_178_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17406_ _04661_ _04660_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__nand2b_1
X_14618_ _11774_ _11775_ _11782_ VGND VGND VPWR VPWR _11783_ sky130_fd_sc_hd__a21o_1
XFILLER_60_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18386_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[29\]
+ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__xor2_1
XFILLER_33_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15598_ _12652_ _12653_ VGND VGND VPWR VPWR _12654_ sky130_fd_sc_hd__nor2_1
XFILLER_92_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14549_ _11721_ _11722_ _11723_ VGND VGND VPWR VPWR _11724_ sky130_fd_sc_hd__a21o_1
X_17337_ _04562_ _04593_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17268_ _04498_ _04526_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__xnor2_1
Xclkload101 clknet_leaf_309_clk VGND VGND VPWR VPWR clkload101/X sky130_fd_sc_hd__clkbuf_4
Xclkload112 clknet_leaf_290_clk VGND VGND VPWR VPWR clkload112/X sky130_fd_sc_hd__clkbuf_8
XFILLER_105_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload123 clknet_leaf_296_clk VGND VGND VPWR VPWR clkload123/X sky130_fd_sc_hd__clkbuf_8
Xclkload134 clknet_leaf_273_clk VGND VGND VPWR VPWR clkload134/X sky130_fd_sc_hd__clkbuf_4
X_19007_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[31\]
+ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__xnor2_1
X_16219_ _03565_ _03567_ _03566_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_77_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload145 clknet_leaf_222_clk VGND VGND VPWR VPWR clkload145/Y sky130_fd_sc_hd__clkinv_4
XFILLER_220_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17199_ net120 _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload156 clknet_leaf_212_clk VGND VGND VPWR VPWR clkload156/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload167 clknet_leaf_240_clk VGND VGND VPWR VPWR clkload167/Y sky130_fd_sc_hd__bufinv_16
XFILLER_143_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload178 clknet_leaf_234_clk VGND VGND VPWR VPWR clkload178/Y sky130_fd_sc_hd__clkinv_4
XFILLER_143_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload189 clknet_leaf_24_clk VGND VGND VPWR VPWR clkload189/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_226_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19909_ _06867_ _06869_ _06905_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__nand3_1
XFILLER_216_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1004 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_239_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_204_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_204_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22920_ _09598_ _09597_ VGND VGND VPWR VPWR _09599_ sky130_fd_sc_hd__nand2b_1
XFILLER_151_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_235_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_235_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22851_ systolic_inst.B_outs\[1\]\[7\] _09531_ VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__nand2_1
XFILLER_84_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21802_ _08605_ _08606_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__nor2_1
XFILLER_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25570_ systolic_inst.acc_wires\[1\]\[14\] C_out\[46\] net35 VGND VGND VPWR VPWR
+ _02872_ sky130_fd_sc_hd__mux2_1
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22782_ _09459_ _09460_ _09463_ VGND VGND VPWR VPWR _09465_ sky130_fd_sc_hd__a21o_1
XFILLER_227_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24521_ C_out\[87\] net100 net82 ser_C.shift_reg\[87\] _10730_ VGND VGND VPWR VPWR
+ _02337_ sky130_fd_sc_hd__a221o_1
XFILLER_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21733_ _08482_ _08539_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__nand2_1
XFILLER_101_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27240_ clknet_leaf_279_clk _01038_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24452_ net114 ser_C.shift_reg\[54\] VGND VGND VPWR VPWR _10696_ sky130_fd_sc_hd__and2_1
XFILLER_197_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21664_ _08471_ _08472_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__nor2_1
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_135_Left_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23403_ systolic_inst.B_outs\[0\]\[7\] _10028_ VGND VGND VPWR VPWR _10029_ sky130_fd_sc_hd__xor2_1
X_20615_ _07543_ _07544_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__xnor2_1
X_27171_ clknet_leaf_253_clk _00969_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24383_ C_out\[18\] net104 _10643_ ser_C.shift_reg\[18\] _10661_ VGND VGND VPWR VPWR
+ _02268_ sky130_fd_sc_hd__a221o_1
XFILLER_193_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21595_ systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[6\] systolic_inst.A_outs\[3\]\[7\]
+ systolic_inst.B_outs\[3\]\[0\] VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__a22o_1
XFILLER_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26122_ deser_B.serial_word\[77\] deser_B.shift_reg\[77\] net55 VGND VGND VPWR VPWR
+ _03424_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23334_ _09961_ _09962_ _09941_ VGND VGND VPWR VPWR _09963_ sky130_fd_sc_hd__mux2_1
XFILLER_20_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20546_ _07465_ _07478_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_211_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26053_ deser_B.serial_word\[8\] deser_B.shift_reg\[8\] net55 VGND VGND VPWR VPWR
+ _03355_ sky130_fd_sc_hd__mux2_1
XFILLER_193_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23265_ systolic_inst.acc_wires\[1\]\[28\] systolic_inst.acc_wires\[1\]\[29\] systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09908_ sky130_fd_sc_hd__o21ai_1
XFILLER_192_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20477_ _07368_ _07376_ _07375_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__a21bo_1
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25004_ net111 ser_C.shift_reg\[330\] VGND VGND VPWR VPWR _10972_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_197_Right_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22216_ systolic_inst.A_outs\[2\]\[1\] systolic_inst.B_outs\[2\]\[6\] _08961_ VGND
+ VGND VPWR VPWR _08962_ sky130_fd_sc_hd__and3_1
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23196_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[19\]
+ VGND VGND VPWR VPWR _09850_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22147_ _08893_ _08894_ VGND VGND VPWR VPWR _08895_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_144_Left_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22078_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.A_outs\[1\]\[0\] net122 VGND
+ VGND VPWR VPWR _01778_ sky130_fd_sc_hd__mux2_1
XFILLER_134_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26955_ clknet_leaf_2_A_in_serial_clk _00753_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25906_ systolic_inst.acc_wires\[11\]\[30\] C_out\[382\] net40 VGND VGND VPWR VPWR
+ _03208_ sky130_fd_sc_hd__mux2_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13920_ deser_A.serial_word\[81\] deser_A.shift_reg\[81\] net57 VGND VGND VPWR VPWR
+ _00746_ sky130_fd_sc_hd__mux2_1
X_21029_ _07843_ _07861_ _07859_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__o21a_1
X_29674_ clknet_leaf_31_B_in_serial_clk _03469_ net134 VGND VGND VPWR VPWR deser_B.serial_word\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26886_ clknet_leaf_8_A_in_serial_clk _00684_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28625_ clknet_leaf_147_clk _02423_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[173\]
+ sky130_fd_sc_hd__dfrtp_1
X_13851_ deser_A.serial_word\[12\] deser_A.shift_reg\[12\] net58 VGND VGND VPWR VPWR
+ _00677_ sky130_fd_sc_hd__mux2_1
XFILLER_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25837_ systolic_inst.acc_wires\[9\]\[25\] C_out\[313\] net13 VGND VGND VPWR VPWR
+ _03139_ sky130_fd_sc_hd__mux2_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28556_ clknet_leaf_172_clk _02354_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_13782_ B_in\[89\] deser_B.word_buffer\[89\] net89 VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__mux2_1
X_16570_ net108 systolic_inst.acc_wires\[12\]\[30\] net67 _03916_ VGND VGND VPWR VPWR
+ _01200_ sky130_fd_sc_hd__a22o_1
XFILLER_222_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25768_ systolic_inst.acc_wires\[7\]\[20\] C_out\[244\] net44 VGND VGND VPWR VPWR
+ _03070_ sky130_fd_sc_hd__mux2_1
XFILLER_55_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15521_ _12578_ _12575_ VGND VGND VPWR VPWR _12579_ sky130_fd_sc_hd__and2b_1
X_27507_ clknet_leaf_229_clk _01305_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24719_ C_out\[186\] net99 net79 ser_C.shift_reg\[186\] _10829_ VGND VGND VPWR VPWR
+ _02436_ sky130_fd_sc_hd__a221o_1
X_28487_ clknet_leaf_113_clk _02285_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_25699_ systolic_inst.acc_wires\[5\]\[15\] C_out\[175\] net31 VGND VGND VPWR VPWR
+ _03001_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_153_Left_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15452_ _12511_ _12508_ VGND VGND VPWR VPWR _12512_ sky130_fd_sc_hd__and2b_1
XFILLER_54_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18240_ net66 _05416_ _05417_ systolic_inst.acc_wires\[9\]\[7\] net107 VGND VGND
+ VPWR VPWR _01369_ sky130_fd_sc_hd__a32o_1
XFILLER_31_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27438_ clknet_leaf_247_clk _01236_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_230_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _11580_ _11584_ VGND VGND VPWR VPWR _11586_ sky130_fd_sc_hd__or2_1
X_15383_ _12439_ _12445_ VGND VGND VPWR VPWR _12447_ sky130_fd_sc_hd__xnor2_1
X_18171_ _05291_ _05334_ _05333_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__o21a_1
XFILLER_169_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27369_ clknet_leaf_339_clk _01167_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29108_ clknet_leaf_162_clk _02906_ net150 VGND VGND VPWR VPWR C_out\[80\] sky130_fd_sc_hd__dfrtp_1
XFILLER_168_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17122_ net62 _04411_ _04412_ systolic_inst.acc_wires\[11\]\[22\] net105 VGND VGND
+ VPWR VPWR _01256_ sky130_fd_sc_hd__a32o_1
X_14334_ _11516_ _11517_ VGND VGND VPWR VPWR _11519_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_169_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17053_ _04352_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__nor2_1
X_29039_ clknet_leaf_122_clk _02837_ net153 VGND VGND VPWR VPWR C_out\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14265_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[5\] VGND VGND
+ VPWR VPWR _11452_ sky130_fd_sc_hd__nand2_1
XFILLER_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16004_ _13000_ _13001_ VGND VGND VPWR VPWR _13003_ sky130_fd_sc_hd__xnor2_1
X_13216_ deser_A.word_buffer\[54\] deser_A.serial_word\[54\] net128 VGND VGND VPWR
+ VPWR _00064_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14196_ _11360_ _11384_ VGND VGND VPWR VPWR _11385_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13147_ ser_C.bit_idx\[0\] ser_C.bit_idx\[3\] _11298_ VGND VGND VPWR VPWR _11299_
+ sky130_fd_sc_hd__and3_1
XFILLER_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17955_ _05119_ _05121_ _05120_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__o21bai_1
XFILLER_61_1324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16906_ _04221_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__nand2_1
X_17886_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[5\]
+ systolic_inst.A_outs\[9\]\[6\] VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__and4_1
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19625_ systolic_inst.B_outs\[5\]\[5\] systolic_inst.B_outs\[1\]\[5\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__mux2_1
X_16837_ _04153_ _04154_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__and2_1
XFILLER_66_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19556_ net62 _06589_ _06590_ systolic_inst.acc_wires\[7\]\[22\] net105 VGND VGND
+ VPWR VPWR _01512_ sky130_fd_sc_hd__a32o_1
X_16768_ _04087_ _04088_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__nand2_1
XFILLER_34_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18507_ systolic_inst.A_outs\[8\]\[1\] systolic_inst.B_outs\[8\]\[6\] VGND VGND VPWR
+ VPWR _05638_ sky130_fd_sc_hd__nand2_1
XFILLER_206_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15719_ net108 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[13\] _12771_
+ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19487_ _06528_ _06529_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__nor2_1
X_16699_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[6\]
+ systolic_inst.A_outs\[11\]\[7\] VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__nand4_1
XFILLER_224_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18438_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[2\]
+ systolic_inst.A_outs\[8\]\[3\] VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__nand4_2
XFILLER_107_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18369_ systolic_inst.acc_wires\[9\]\[24\] systolic_inst.acc_wires\[9\]\[25\] systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_79_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20400_ _07296_ _07336_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__xnor2_1
X_21380_ _08223_ _08224_ _08225_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_228_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20331_ _07265_ _07266_ _07269_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__and3_1
XFILLER_179_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23050_ _09724_ _09723_ VGND VGND VPWR VPWR _09725_ sky130_fd_sc_hd__and2b_1
X_20262_ _07198_ _07203_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22001_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[20\]
+ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__or2_1
XFILLER_89_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20193_ net106 systolic_inst.acc_wires\[6\]\[26\] net62 _07159_ VGND VGND VPWR VPWR
+ _01580_ sky130_fd_sc_hd__a22o_1
XFILLER_66_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26740_ clknet_leaf_98_clk _00542_ net5 VGND VGND VPWR VPWR B_in\[12\] sky130_fd_sc_hd__dfrtp_1
X_23952_ net115 net131 VGND VGND VPWR VPWR _10505_ sky130_fd_sc_hd__and2_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22903_ _09546_ _09549_ VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__nand2_1
X_26671_ clknet_leaf_8_B_in_serial_clk _00474_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23883_ _11258_ systolic_inst.acc_wires\[0\]\[29\] net64 _10470_ VGND VGND VPWR VPWR
+ _01959_ sky130_fd_sc_hd__a22o_1
XFILLER_45_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28410_ clknet_leaf_82_clk _02208_ VGND VGND VPWR VPWR systolic_inst.B_shift\[17\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25622_ systolic_inst.acc_wires\[3\]\[2\] C_out\[98\] net48 VGND VGND VPWR VPWR _02924_
+ sky130_fd_sc_hd__mux2_1
X_22834_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[7\]
+ VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__o21ai_2
XFILLER_38_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29390_ clknet_leaf_241_clk _03188_ net145 VGND VGND VPWR VPWR C_out\[362\] sky130_fd_sc_hd__dfrtp_1
XFILLER_112_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25553_ systolic_inst.acc_wires\[0\]\[29\] C_out\[29\] net53 VGND VGND VPWR VPWR
+ _02855_ sky130_fd_sc_hd__mux2_1
XFILLER_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28341_ clknet_leaf_342_clk _02139_ VGND VGND VPWR VPWR systolic_inst.A_shift\[25\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_22765_ systolic_inst.A_outs\[1\]\[4\] _09409_ _09426_ _09425_ _09422_ VGND VGND
+ VPWR VPWR _09448_ sky130_fd_sc_hd__a32o_1
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24504_ net113 ser_C.shift_reg\[80\] VGND VGND VPWR VPWR _10722_ sky130_fd_sc_hd__and2_1
XFILLER_197_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21716_ systolic_inst.A_outs\[3\]\[3\] systolic_inst.A_outs\[3\]\[4\] systolic_inst.B_outs\[3\]\[6\]
+ systolic_inst.B_outs\[3\]\[7\] VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__and4b_1
X_28272_ clknet_leaf_134_clk _02070_ VGND VGND VPWR VPWR systolic_inst.B_shift\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25484_ systolic_inst.cycle_cnt\[17\] systolic_inst.cycle_cnt\[16\] _11216_ VGND
+ VGND VPWR VPWR _11220_ sky130_fd_sc_hd__and3_1
XFILLER_164_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22696_ systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[2\]
+ systolic_inst.B_outs\[1\]\[0\] VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__a22oi_1
XFILLER_197_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_213_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24435_ C_out\[44\] _11302_ net81 ser_C.shift_reg\[44\] _10687_ VGND VGND VPWR VPWR
+ _02294_ sky130_fd_sc_hd__a221o_1
XFILLER_40_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27223_ clknet_leaf_291_clk _01021_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_21647_ _08454_ _08455_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__nor2_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27154_ clknet_leaf_251_clk _00952_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_24366_ net7 ser_C.shift_reg\[11\] VGND VGND VPWR VPWR _10653_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_151_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21578_ _08386_ _08388_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_151_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26105_ deser_B.serial_word\[60\] deser_B.shift_reg\[60\] net56 VGND VGND VPWR VPWR
+ _03407_ sky130_fd_sc_hd__mux2_1
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23317_ systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[4\] VGND VGND VPWR
+ VPWR _09946_ sky130_fd_sc_hd__nand2_1
X_20529_ _07323_ _07461_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__or2_1
XFILLER_158_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27085_ clknet_leaf_32_B_in_serial_clk _00883_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_24297_ systolic_inst.A_shift\[12\]\[4\] A_in\[52\] net59 VGND VGND VPWR VPWR _10622_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14050_ deser_B.shift_reg\[84\] deser_B.shift_reg\[85\] net125 VGND VGND VPWR VPWR
+ _00876_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26036_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.B_outs\[11\]\[0\] net118 VGND
+ VGND VPWR VPWR _03338_ sky130_fd_sc_hd__mux2_1
X_23248_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[27\]
+ VGND VGND VPWR VPWR _09894_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23179_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[16\]
+ VGND VGND VPWR VPWR _09836_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_27987_ clknet_leaf_144_clk _01785_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_82_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17740_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[24\]
+ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__and2_1
X_14952_ _12031_ _12071_ VGND VGND VPWR VPWR _12073_ sky130_fd_sc_hd__and2_1
X_26938_ clknet_leaf_20_A_in_serial_clk _00736_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13903_ deser_A.serial_word\[64\] deser_A.shift_reg\[64\] net57 VGND VGND VPWR VPWR
+ _00729_ sky130_fd_sc_hd__mux2_1
X_29657_ clknet_leaf_7_B_in_serial_clk _03452_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_17671_ _04904_ _04905_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__and2_1
X_26869_ clknet_leaf_14_A_in_serial_clk _00667_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14883_ systolic_inst.A_outs\[14\]\[2\] systolic_inst.B_outs\[14\]\[5\] VGND VGND
+ VPWR VPWR _12006_ sky130_fd_sc_hd__nand2_1
XFILLER_75_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19410_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[7\]\[0\]
+ _06462_ _06463_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__a22o_1
XFILLER_1_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28608_ clknet_leaf_135_clk _02406_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16622_ _03945_ _03946_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__nand2_1
XFILLER_210_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13834_ _11327_ VGND VGND VPWR VPWR _11328_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap50 net51 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_8
X_29588_ clknet_leaf_12_B_in_serial_clk _03383_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_161_Left_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap61 _11713_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_104_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap72 _11332_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_12
XFILLER_216_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19341_ _06399_ _06400_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__nor2_1
X_28539_ clknet_leaf_159_clk _02337_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_13765_ B_in\[72\] deser_B.word_buffer\[72\] net88 VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__mux2_1
X_16553_ _03884_ _03885_ _03898_ _03901_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__or4_1
Xmax_cap83 _10505_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_12
Xmax_cap94 net95 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_8
XFILLER_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15504_ _12546_ _12562_ VGND VGND VPWR VPWR _12563_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_100_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19272_ _06333_ _06334_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__nor2_1
XFILLER_43_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13696_ B_in\[3\] deser_B.word_buffer\[3\] net86 VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__mux2_1
X_16484_ _03841_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__and2_1
XFILLER_94_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_233_Right_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18223_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[9\]\[5\]
+ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__nand2_1
XFILLER_188_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15435_ _12494_ _12495_ VGND VGND VPWR VPWR _12496_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_61_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15366_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.B_outs\[8\]\[2\] net115 VGND
+ VGND VPWR VPWR _01084_ sky130_fd_sc_hd__mux2_1
X_18154_ _05307_ _05310_ _05340_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_113_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17105_ _04376_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__nor2_1
XFILLER_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14317_ _11502_ _11501_ VGND VGND VPWR VPWR _11503_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_74_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15297_ _12379_ _12381_ VGND VGND VPWR VPWR _12389_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_74_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18085_ _05273_ _05274_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_170_Left_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14248_ _11426_ _11428_ VGND VGND VPWR VPWR _11435_ sky130_fd_sc_hd__nor2_1
X_17036_ _04332_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__nand2_1
XFILLER_109_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14179_ _11365_ _11368_ VGND VGND VPWR VPWR _11369_ sky130_fd_sc_hd__xnor2_1
XFILLER_217_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18987_ systolic_inst.acc_wires\[8\]\[26\] systolic_inst.acc_wires\[8\]\[27\] systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__o21a_1
XFILLER_140_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17938_ _05096_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__or2_1
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17869_ _05059_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__nand2b_1
XFILLER_226_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19608_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[31\]
+ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_217_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20880_ systolic_inst.A_outs\[4\]\[2\] systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[3\]
+ systolic_inst.B_outs\[4\]\[1\] VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_217_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_217_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19539_ _06554_ _06575_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__nor2_1
XFILLER_53_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22550_ _09272_ _09273_ _09274_ VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__and3_1
XFILLER_22_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_200_Right_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21501_ systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[3\]
+ systolic_inst.B_outs\[3\]\[0\] VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__a22o_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22481_ _09213_ _09214_ _09215_ VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__a21o_1
XFILLER_72_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24220_ _10595_ systolic_inst.A_shift\[19\]\[1\] net70 VGND VGND VPWR VPWR _02171_
+ sky130_fd_sc_hd__mux2_1
X_21432_ _08262_ _08264_ _08270_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__a21o_1
XFILLER_72_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24151_ systolic_inst.A_shift\[29\]\[7\] A_in\[111\] net59 VGND VGND VPWR VPWR _10577_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21363_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[16\]
+ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__or2_1
X_23102_ _09767_ _09768_ _09769_ VGND VGND VPWR VPWR _09770_ sky130_fd_sc_hd__a21o_1
XFILLER_200_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20314_ net109 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[5\] _07252_
+ _07253_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__a22o_1
X_24082_ systolic_inst.B_shift\[2\]\[1\] _11332_ net83 systolic_inst.B_shift\[6\]\[1\]
+ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__a22o_1
XFILLER_116_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21294_ _08143_ _08147_ _08150_ _08151_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__o211a_1
XFILLER_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23033_ _09706_ _09707_ VGND VGND VPWR VPWR _09709_ sky130_fd_sc_hd__nor2_1
X_27910_ clknet_leaf_44_clk _01708_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20245_ net107 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _07188_ sky130_fd_sc_hd__and2_1
XFILLER_162_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28890_ clknet_leaf_287_clk _02688_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[438\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_206_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27841_ clknet_leaf_205_clk _01639_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_20176_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[24\]
+ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_206_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27772_ clknet_leaf_186_clk _01570_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_170_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_202_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24984_ net111 ser_C.shift_reg\[320\] VGND VGND VPWR VPWR _10962_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_198_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_835 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29511_ clknet_leaf_264_clk _03309_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[483\]
+ sky130_fd_sc_hd__dfrtp_1
X_26723_ clknet_leaf_32_B_in_serial_clk _00526_ net134 VGND VGND VPWR VPWR deser_B.word_buffer\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_198_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23935_ systolic_inst.A_shift\[3\]\[7\] net71 _11333_ A_in\[31\] VGND VGND VPWR VPWR
+ _01985_ sky130_fd_sc_hd__a22o_1
XFILLER_218_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29442_ clknet_leaf_333_clk _03240_ net131 VGND VGND VPWR VPWR C_out\[414\] sky130_fd_sc_hd__dfrtp_1
X_23866_ _11258_ systolic_inst.acc_wires\[0\]\[26\] net64 _10456_ VGND VGND VPWR VPWR
+ _01956_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26654_ clknet_leaf_24_B_in_serial_clk _00457_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25605_ systolic_inst.acc_wires\[2\]\[17\] C_out\[81\] net52 VGND VGND VPWR VPWR
+ _02907_ sky130_fd_sc_hd__mux2_1
X_22817_ _09464_ _09498_ VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__xnor2_1
X_29373_ clknet_leaf_234_clk _03171_ net145 VGND VGND VPWR VPWR C_out\[345\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23797_ _10394_ _10395_ _10389_ VGND VGND VPWR VPWR _10398_ sky130_fd_sc_hd__or3b_1
X_26585_ clknet_leaf_29_A_in_serial_clk _00388_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_13550_ deser_A.shift_reg\[114\] deser_A.shift_reg\[115\] net129 VGND VGND VPWR VPWR
+ _00387_ sky130_fd_sc_hd__mux2_1
X_28324_ clknet_leaf_3_clk _02122_ VGND VGND VPWR VPWR systolic_inst.A_shift\[27\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25536_ systolic_inst.acc_wires\[0\]\[12\] C_out\[12\] net33 VGND VGND VPWR VPWR
+ _02838_ sky130_fd_sc_hd__mux2_1
X_22748_ systolic_inst.A_outs\[1\]\[2\] systolic_inst.B_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\]
+ systolic_inst.A_outs\[1\]\[1\] VGND VGND VPWR VPWR _09432_ sky130_fd_sc_hd__a22oi_2
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25467_ systolic_inst.cycle_cnt\[10\] _11306_ _11199_ _11202_ systolic_inst.cycle_cnt\[11\]
+ VGND VGND VPWR VPWR _11209_ sky130_fd_sc_hd__a41o_1
X_28255_ clknet_leaf_79_clk _02053_ VGND VGND VPWR VPWR systolic_inst.B_shift\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13481_ deser_A.shift_reg\[45\] deser_A.shift_reg\[46\] net130 VGND VGND VPWR VPWR
+ _00318_ sky130_fd_sc_hd__mux2_1
X_22679_ systolic_inst.A_outs\[1\]\[6\] systolic_inst.A_outs\[0\]\[6\] net121 VGND
+ VGND VPWR VPWR _01848_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15220_ _12321_ _12322_ VGND VGND VPWR VPWR _12323_ sky130_fd_sc_hd__nand2_1
X_24418_ net114 ser_C.shift_reg\[37\] VGND VGND VPWR VPWR _10679_ sky130_fd_sc_hd__and2_1
X_27206_ clknet_leaf_258_clk _01004_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28186_ clknet_leaf_17_clk _01984_ VGND VGND VPWR VPWR systolic_inst.A_shift\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25398_ _11168_ systolic_inst.A_shift\[2\]\[6\] net71 VGND VGND VPWR VPWR _02776_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15151_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[14\]\[1\]
+ VGND VGND VPWR VPWR _12264_ sky130_fd_sc_hd__or2_1
XFILLER_51_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27137_ clknet_leaf_86_clk _00935_ VGND VGND VPWR VPWR systolic_inst.B_shift\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_24349_ C_out\[1\] net104 _10643_ ser_C.shift_reg\[1\] _10644_ VGND VGND VPWR VPWR
+ _02251_ sky130_fd_sc_hd__a221o_1
XFILLER_154_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14102_ systolic_inst.A_shift\[12\]\[2\] net72 _11333_ A_in\[58\] VGND VGND VPWR
+ VPWR _00924_ sky130_fd_sc_hd__a22o_1
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27068_ clknet_leaf_9_B_in_serial_clk _00866_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_15082_ _12197_ _12198_ VGND VGND VPWR VPWR _12200_ sky130_fd_sc_hd__and2_1
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14033_ deser_B.shift_reg\[67\] deser_B.shift_reg\[68\] net126 VGND VGND VPWR VPWR
+ _00859_ sky130_fd_sc_hd__mux2_1
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26019_ systolic_inst.acc_wires\[15\]\[15\] ser_C.parallel_data\[495\] net37 VGND
+ VGND VPWR VPWR _03321_ sky130_fd_sc_hd__mux2_1
X_18910_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[16\]
+ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__or2_1
XFILLER_101_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19890_ net119 _06887_ _06888_ _06852_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18841_ net63 _05954_ _05955_ systolic_inst.acc_wires\[8\]\[6\] net108 VGND VGND
+ VPWR VPWR _01432_ sky130_fd_sc_hd__a32o_1
XFILLER_110_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18772_ _05892_ _05893_ _05894_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__a21oi_1
X_15984_ _12981_ _12982_ _12983_ VGND VGND VPWR VPWR _12984_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_106_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[22\]
+ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__nand2_1
X_14935_ _12054_ _12055_ VGND VGND VPWR VPWR _12057_ sky130_fd_sc_hd__xor2_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17654_ _04868_ _04871_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__and3b_1
XFILLER_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14866_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[6\] _11987_
+ _11989_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16605_ net118 _03930_ _03931_ _03924_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__a31o_1
X_13817_ B_in\[124\] deser_B.word_buffer\[124\] net89 VGND VGND VPWR VPWR _00654_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17585_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[10\]\[2\]
+ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__nand2_1
X_14797_ _11903_ _11922_ VGND VGND VPWR VPWR _11923_ sky130_fd_sc_hd__nor2_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19324_ _06348_ _06384_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16536_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[25\]
+ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__xor2_1
XFILLER_204_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13748_ B_in\[55\] deser_B.word_buffer\[55\] net85 VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__mux2_1
XFILLER_73_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19255_ _06282_ _06284_ _06283_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__o21ba_1
XFILLER_143_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16467_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[15\]
+ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__nor2_1
X_13679_ deser_B.word_buffer\[115\] deser_B.serial_word\[115\] net124 VGND VGND VPWR
+ VPWR _00516_ sky130_fd_sc_hd__mux2_1
X_18206_ _05388_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__inv_2
X_15418_ _12461_ _12477_ _12478_ VGND VGND VPWR VPWR _12480_ sky130_fd_sc_hd__and3_1
XFILLER_192_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19186_ _06249_ _06250_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__nor2_1
XFILLER_145_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16398_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[12\]\[5\]
+ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_136_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18137_ _05296_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__xnor2_1
X_15349_ _12429_ _12432_ VGND VGND VPWR VPWR _12433_ sky130_fd_sc_hd__nand2_1
XFILLER_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18068_ _05150_ _05256_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17019_ net69 _04323_ _04324_ systolic_inst.acc_wires\[11\]\[7\] net105 VGND VGND
+ VPWR VPWR _01241_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_93_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_242_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20030_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[6\]\[3\]
+ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__nand2_1
XFILLER_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21981_ _08765_ _08764_ VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__and2b_1
XFILLER_67_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23720_ _10332_ VGND VGND VPWR VPWR _10333_ sky130_fd_sc_hd__inv_2
XFILLER_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20932_ _07780_ _07782_ _07806_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__a21oi_1
XFILLER_226_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23651_ _10269_ _10270_ VGND VGND VPWR VPWR _10271_ sky130_fd_sc_hd__nor2_1
XFILLER_82_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20863_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[2\]
+ systolic_inst.B_outs\[4\]\[2\] VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__nand4_2
XFILLER_242_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22602_ systolic_inst.acc_wires\[2\]\[16\] systolic_inst.acc_wires\[2\]\[17\] systolic_inst.acc_wires\[2\]\[18\]
+ systolic_inst.acc_wires\[2\]\[19\] systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__o41a_1
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26370_ clknet_leaf_27_clk _00177_ net133 VGND VGND VPWR VPWR A_in\[38\] sky130_fd_sc_hd__dfrtp_1
XFILLER_241_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23582_ _10196_ _10202_ VGND VGND VPWR VPWR _10204_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_18_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20794_ systolic_inst.acc_wires\[5\]\[24\] systolic_inst.acc_wires\[5\]\[25\] systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__o21a_1
XFILLER_223_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25321_ ser_C.parallel_data\[487\] net97 net77 ser_C.shift_reg\[487\] _11130_ VGND
+ VGND VPWR VPWR _02737_ sky130_fd_sc_hd__a221o_1
X_22533_ _09258_ _09259_ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_46_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28040_ clknet_leaf_163_clk _01838_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_25252_ net111 ser_C.shift_reg\[454\] VGND VGND VPWR VPWR _11096_ sky130_fd_sc_hd__and2_1
X_22464_ _09200_ _09201_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__xnor2_1
XFILLER_210_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24203_ systolic_inst.A_shift\[21\]\[1\] A_in\[81\] net59 VGND VGND VPWR VPWR _10587_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21415_ _08209_ _08210_ _08235_ _08255_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__a211o_1
XFILLER_124_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25183_ C_out\[418\] net103 net75 ser_C.shift_reg\[418\] _11061_ VGND VGND VPWR VPWR
+ _02668_ sky130_fd_sc_hd__a221o_1
X_22395_ _09096_ _09135_ VGND VGND VPWR VPWR _09136_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24134_ _10568_ systolic_inst.A_shift\[29\]\[6\] net71 VGND VGND VPWR VPWR _02112_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21346_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[4\]\[14\]
+ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_208_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_208_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24065_ systolic_inst.B_shift\[19\]\[4\] B_in\[28\] net59 VGND VGND VPWR VPWR _10550_
+ sky130_fd_sc_hd__mux2_1
XFILLER_118_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28942_ clknet_leaf_246_clk _02740_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21277_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[4\]\[4\]
+ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__nand2_1
XFILLER_104_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_13__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_13__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_204_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23016_ _09658_ _09661_ _09690_ VGND VGND VPWR VPWR _09692_ sky130_fd_sc_hd__or3_1
XFILLER_150_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20228_ systolic_inst.A_outs\[5\]\[5\] systolic_inst.A_outs\[4\]\[5\] net116 VGND
+ VGND VPWR VPWR _01591_ sky130_fd_sc_hd__mux2_1
X_28873_ clknet_leaf_293_clk _02671_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[421\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27824_ clknet_leaf_217_clk _01622_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_196_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[22\]
+ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_142_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27755_ clknet_leaf_207_clk _01553_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24967_ C_out\[310\] net103 net76 ser_C.shift_reg\[310\] _10953_ VGND VGND VPWR VPWR
+ _02560_ sky130_fd_sc_hd__a221o_1
XFILLER_91_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26706_ clknet_leaf_9_B_in_serial_clk _00509_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_14720_ _11866_ _11869_ VGND VGND VPWR VPWR _11870_ sky130_fd_sc_hd__or2_1
X_23918_ systolic_inst.B_shift\[22\]\[3\] B_in\[83\] net59 VGND VGND VPWR VPWR _10492_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27686_ clknet_leaf_198_clk _01484_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24898_ net110 ser_C.shift_reg\[277\] VGND VGND VPWR VPWR _10919_ sky130_fd_sc_hd__and2_1
XFILLER_73_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29425_ clknet_leaf_338_clk _03223_ net131 VGND VGND VPWR VPWR C_out\[397\] sky130_fd_sc_hd__dfrtp_1
XFILLER_205_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26637_ clknet_leaf_12_B_in_serial_clk _00440_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14651_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[18\]
+ VGND VGND VPWR VPWR _11811_ sky130_fd_sc_hd__nand2_1
XFILLER_33_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23849_ _10422_ _10441_ VGND VGND VPWR VPWR _10442_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13602_ deser_B.word_buffer\[38\] deser_B.serial_word\[38\] net123 VGND VGND VPWR
+ VPWR _00439_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29356_ clknet_leaf_230_clk _03154_ net140 VGND VGND VPWR VPWR C_out\[328\] sky130_fd_sc_hd__dfrtp_1
X_17370_ _04626_ _04625_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__nand2b_1
X_26568_ clknet_leaf_23_A_in_serial_clk _00371_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_14582_ _11750_ _11751_ VGND VGND VPWR VPWR _11752_ sky130_fd_sc_hd__and2_1
XFILLER_232_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28307_ clknet_leaf_71_clk _02105_ VGND VGND VPWR VPWR systolic_inst.B_shift\[27\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16321_ _03699_ _03700_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nand2b_1
X_25519_ systolic_inst.cycle_cnt\[30\] _11279_ _11239_ VGND VGND VPWR VPWR _11242_
+ sky130_fd_sc_hd__a21o_1
XFILLER_185_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13533_ deser_A.shift_reg\[97\] deser_A.shift_reg\[98\] net129 VGND VGND VPWR VPWR
+ _00370_ sky130_fd_sc_hd__mux2_1
X_29287_ clknet_leaf_323_clk _03085_ net142 VGND VGND VPWR VPWR C_out\[259\] sky130_fd_sc_hd__dfrtp_1
X_26499_ clknet_leaf_6_A_in_serial_clk _00302_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_207_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19040_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[2\] _06109_ VGND
+ VGND VPWR VPWR _06111_ sky130_fd_sc_hd__a21o_1
XFILLER_186_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28238_ clknet_leaf_130_clk _02036_ VGND VGND VPWR VPWR systolic_inst.B_shift\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13464_ deser_A.shift_reg\[28\] deser_A.shift_reg\[29\] deser_A.receiving VGND VGND
+ VPWR VPWR _00301_ sky130_fd_sc_hd__mux2_1
X_16252_ systolic_inst.A_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[5\] systolic_inst.B_outs\[12\]\[6\]
+ systolic_inst.B_outs\[12\]\[7\] VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__and4b_1
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15203_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[14\]\[9\]
+ VGND VGND VPWR VPWR _12308_ sky130_fd_sc_hd__xor2_1
X_28169_ clknet_leaf_81_clk _01967_ VGND VGND VPWR VPWR systolic_inst.B_shift\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16183_ systolic_inst.A_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[6\] _11260_ systolic_inst.A_outs\[12\]\[2\]
+ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__o2bb2a_1
X_13395_ A_in\[104\] deser_A.word_buffer\[104\] net96 VGND VGND VPWR VPWR _00243_
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15134_ _12199_ _12203_ _12226_ _12227_ VGND VGND VPWR VPWR _12250_ sky130_fd_sc_hd__o31a_1
XFILLER_127_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19942_ _06938_ _06937_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__and2b_1
XFILLER_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15065_ _12180_ _12181_ VGND VGND VPWR VPWR _12183_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14016_ deser_B.shift_reg\[50\] deser_B.shift_reg\[51\] net125 VGND VGND VPWR VPWR
+ _00842_ sky130_fd_sc_hd__mux2_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19873_ _06829_ _06837_ _06836_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__a21bo_1
XFILLER_141_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18824_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[8\]\[4\]
+ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__nand2_1
XFILLER_68_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18755_ _05835_ _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__xor2_1
X_15967_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[7\]\[0\] net119 VGND
+ VGND VPWR VPWR _01146_ sky130_fd_sc_hd__mux2_1
XFILLER_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17706_ _04934_ _04935_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14918_ _12038_ _12039_ VGND VGND VPWR VPWR _12040_ sky130_fd_sc_hd__xnor2_1
XFILLER_237_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18686_ _05771_ _05773_ _05772_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__o21ba_1
XFILLER_97_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15898_ _12924_ _12925_ VGND VGND VPWR VPWR _12926_ sky130_fd_sc_hd__and2_1
XFILLER_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17637_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[10\]\[10\]
+ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__nand2_1
XFILLER_224_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14849_ _11969_ _11972_ VGND VGND VPWR VPWR _11973_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17568_ _04601_ _04738_ _04809_ _04807_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__a31o_1
XFILLER_189_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19307_ _06329_ _06331_ _06366_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__a21oi_1
X_16519_ _03866_ _03867_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__and2b_1
XFILLER_20_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17499_ _04714_ _04751_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19238_ _06299_ _06300_ _06301_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__and3_1
XFILLER_34_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19169_ _06171_ _06206_ _06205_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__a21bo_1
XFILLER_121_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21200_ _08066_ _08067_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__or2_1
XFILLER_195_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22180_ systolic_inst.A_outs\[2\]\[1\] systolic_inst.B_outs\[2\]\[5\] systolic_inst.B_outs\[2\]\[6\]
+ systolic_inst.A_outs\[2\]\[0\] VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__a22oi_1
XFILLER_133_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21131_ systolic_inst.A_outs\[4\]\[4\] _11271_ _07850_ VGND VGND VPWR VPWR _08001_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_54_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21062_ _07931_ _07932_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__xor2_1
XFILLER_8_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20013_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[6\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__a21o_1
XFILLER_24_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25870_ systolic_inst.acc_wires\[10\]\[26\] C_out\[346\] net11 VGND VGND VPWR VPWR
+ _03172_ sky130_fd_sc_hd__mux2_1
XFILLER_28_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24821_ C_out\[237\] net99 net79 ser_C.shift_reg\[237\] _10880_ VGND VGND VPWR VPWR
+ _02487_ sky130_fd_sc_hd__a221o_1
XFILLER_101_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27540_ clknet_leaf_34_clk _01338_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_21964_ _08742_ _08746_ _08749_ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__a21o_1
X_24752_ net113 ser_C.shift_reg\[204\] VGND VGND VPWR VPWR _10846_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_191_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23703_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[0\]\[0\]
+ _10312_ _10310_ VGND VGND VPWR VPWR _10318_ sky130_fd_sc_hd__a31o_1
XFILLER_76_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20915_ _07788_ _07789_ _07790_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__nand3_1
X_24683_ C_out\[168\] net104 net76 ser_C.shift_reg\[168\] _10811_ VGND VGND VPWR VPWR
+ _02418_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_48_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27471_ clknet_leaf_222_clk _01269_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_21895_ _08682_ _08686_ _08689_ _08690_ VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__o211a_1
XFILLER_82_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29210_ clknet_leaf_181_clk _03008_ net146 VGND VGND VPWR VPWR C_out\[182\] sky130_fd_sc_hd__dfrtp_1
XFILLER_202_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23634_ _10253_ _10254_ VGND VGND VPWR VPWR _10255_ sky130_fd_sc_hd__nor2_1
X_26422_ clknet_leaf_12_clk _00229_ net134 VGND VGND VPWR VPWR A_in\[90\] sky130_fd_sc_hd__dfrtp_1
X_20846_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[1\]
+ systolic_inst.A_outs\[4\]\[0\] VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__a22o_1
X_29141_ clknet_leaf_166_clk _02939_ net152 VGND VGND VPWR VPWR C_out\[113\] sky130_fd_sc_hd__dfrtp_1
XFILLER_168_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23565_ systolic_inst.B_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[6\] _10025_ VGND
+ VGND VPWR VPWR _10187_ sky130_fd_sc_hd__a21oi_1
X_26353_ clknet_leaf_19_clk _00160_ net133 VGND VGND VPWR VPWR A_in\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_211_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20777_ _07661_ _07668_ _07673_ _07678_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__nand4_1
XFILLER_204_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22516_ _09243_ _09244_ _09245_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__a21o_1
XFILLER_195_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25304_ net111 ser_C.shift_reg\[480\] VGND VGND VPWR VPWR _11122_ sky130_fd_sc_hd__and2_1
XFILLER_211_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29072_ clknet_leaf_116_clk _02870_ net152 VGND VGND VPWR VPWR C_out\[44\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26284_ clknet_leaf_3_A_in_serial_clk _00092_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23496_ _10080_ _10119_ VGND VGND VPWR VPWR _10120_ sky130_fd_sc_hd__nor2_2
XFILLER_161_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28023_ clknet_leaf_167_clk _01821_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22447_ _09159_ _09162_ _09184_ VGND VGND VPWR VPWR _09186_ sky130_fd_sc_hd__and3_1
X_25235_ ser_C.parallel_data\[444\] net102 net74 ser_C.shift_reg\[444\] _11087_ VGND
+ VGND VPWR VPWR _02694_ sky130_fd_sc_hd__a221o_1
XFILLER_148_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13180_ deser_A.word_buffer\[18\] deser_A.serial_word\[18\] net128 VGND VGND VPWR
+ VPWR _00028_ sky130_fd_sc_hd__mux2_1
X_25166_ net110 ser_C.shift_reg\[411\] VGND VGND VPWR VPWR _11053_ sky130_fd_sc_hd__and2_1
X_22378_ _09085_ _09088_ _09117_ _09118_ VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__or4_1
XFILLER_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24117_ systolic_inst.B_shift\[27\]\[4\] net72 _11333_ B_in\[124\] VGND VGND VPWR
+ VPWR _02102_ sky130_fd_sc_hd__a22o_1
XFILLER_108_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21329_ _08155_ _08157_ _08161_ _08181_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__a211o_1
X_25097_ C_out\[375\] net98 net78 ser_C.shift_reg\[375\] _11018_ VGND VGND VPWR VPWR
+ _02625_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_144_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24048_ _10541_ systolic_inst.B_shift\[0\]\[3\] _11332_ VGND VGND VPWR VPWR _02053_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28925_ clknet_leaf_267_clk _02723_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[473\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28856_ clknet_leaf_336_clk _02654_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[404\]
+ sky130_fd_sc_hd__dfrtp_1
X_16870_ _04128_ _04187_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27807_ clknet_leaf_217_clk _01605_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15821_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[13\]\[11\]
+ VGND VGND VPWR VPWR _12860_ sky130_fd_sc_hd__or2_1
XFILLER_49_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28787_ clknet_leaf_225_clk _02585_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[335\]
+ sky130_fd_sc_hd__dfrtp_1
X_25999_ systolic_inst.acc_wires\[14\]\[27\] ser_C.parallel_data\[475\] net24 VGND
+ VGND VPWR VPWR _03301_ sky130_fd_sc_hd__mux2_1
XFILLER_93_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18540_ systolic_inst.A_outs\[8\]\[2\] systolic_inst.B_outs\[8\]\[5\] VGND VGND VPWR
+ VPWR _05670_ sky130_fd_sc_hd__nand2_1
X_27738_ clknet_leaf_133_clk _01536_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_15752_ net116 _12800_ _12801_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__a21oi_1
X_14703_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[26\]
+ VGND VGND VPWR VPWR _11855_ sky130_fd_sc_hd__or2_1
X_18471_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[4\]
+ systolic_inst.A_outs\[8\]\[5\] VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__and4_1
X_27669_ clknet_leaf_146_clk _01467_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15683_ _12644_ _12705_ _12703_ VGND VGND VPWR VPWR _12737_ sky130_fd_sc_hd__a21oi_1
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29408_ clknet_leaf_196_clk _03206_ net146 VGND VGND VPWR VPWR C_out\[380\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ systolic_inst.A_outs\[10\]\[6\] _04676_ _04675_ VGND VGND VPWR VPWR _04677_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_127_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _11787_ _11792_ _11796_ VGND VGND VPWR VPWR _11797_ sky130_fd_sc_hd__a21oi_1
XFILLER_57_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29339_ clknet_leaf_214_clk _03137_ net149 VGND VGND VPWR VPWR C_out\[311\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17353_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[6\] VGND VGND
+ VPWR VPWR _04610_ sky130_fd_sc_hd__nand2_1
X_14565_ _11737_ VGND VGND VPWR VPWR _11738_ sky130_fd_sc_hd__inv_2
XFILLER_57_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16304_ _03620_ _03624_ _03653_ _03651_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__a31o_1
XFILLER_53_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13516_ deser_A.shift_reg\[80\] deser_A.shift_reg\[81\] net129 VGND VGND VPWR VPWR
+ _00353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17284_ systolic_inst.A_outs\[10\]\[1\] systolic_inst.B_outs\[10\]\[6\] VGND VGND
+ VPWR VPWR _04543_ sky130_fd_sc_hd__nand2_1
X_14496_ systolic_inst.B_outs\[15\]\[5\] systolic_inst.A_outs\[15\]\[7\] _11654_ _11653_
+ VGND VGND VPWR VPWR _11676_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_133_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19023_ systolic_inst.B_outs\[6\]\[4\] systolic_inst.B_outs\[2\]\[4\] net120 VGND
+ VGND VPWR VPWR _01470_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16235_ _03555_ _03580_ _03579_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_58_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload305 clknet_leaf_115_clk VGND VGND VPWR VPWR clkload305/Y sky130_fd_sc_hd__inv_6
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13447_ deser_A.shift_reg\[11\] deser_A.shift_reg\[12\] deser_A.receiving VGND VGND
+ VPWR VPWR _00284_ sky130_fd_sc_hd__mux2_1
Xclkload316 clknet_leaf_111_clk VGND VGND VPWR VPWR clkload316/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload13 clknet_5_15__leaf_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_6
Xclkload24 clknet_5_29__leaf_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__inv_6
Xclkload327 clknet_leaf_168_clk VGND VGND VPWR VPWR clkload327/X sky130_fd_sc_hd__clkbuf_4
XFILLER_127_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload338 clknet_leaf_175_clk VGND VGND VPWR VPWR clkload338/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload35 clknet_leaf_345_clk VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__clkinv_8
XFILLER_103_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload46 clknet_leaf_327_clk VGND VGND VPWR VPWR clkload46/X sky130_fd_sc_hd__clkbuf_4
Xclkload349 clknet_leaf_24_A_in_serial_clk VGND VGND VPWR VPWR clkload349/X sky130_fd_sc_hd__clkbuf_8
XFILLER_220_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16166_ _03508_ _03511_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__o21a_1
X_13378_ A_in\[87\] deser_A.word_buffer\[87\] net95 VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__mux2_1
Xclkload57 clknet_leaf_321_clk VGND VGND VPWR VPWR clkload57/Y sky130_fd_sc_hd__clkinv_8
XFILLER_127_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload68 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload68/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_90_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload79 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload79/Y sky130_fd_sc_hd__clkinvlp_4
X_15117_ _11264_ systolic_inst.A_outs\[14\]\[7\] _12181_ _12205_ VGND VGND VPWR VPWR
+ _12233_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_90_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16097_ _13086_ _13090_ VGND VGND VPWR VPWR _13092_ sky130_fd_sc_hd__and2_1
XFILLER_138_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19925_ _06782_ _06920_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__nand2_1
X_15048_ _12166_ VGND VGND VPWR VPWR _12167_ sky130_fd_sc_hd__inv_2
XFILLER_214_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19856_ _06783_ _06853_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__and2_1
XFILLER_190_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18807_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[8\]\[0\]
+ _05923_ _05924_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__a22o_1
X_19787_ systolic_inst.B_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[4\]
+ systolic_inst.A_outs\[6\]\[5\] VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__and4_1
X_16999_ net69 _04305_ _04307_ systolic_inst.acc_wires\[11\]\[4\] net105 VGND VGND
+ VPWR VPWR _01238_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_88_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18738_ _05861_ _05862_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_237_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_237_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18669_ _05724_ _05757_ _05758_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_48_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_233_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20700_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[5\]\[12\]
+ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__xnor2_1
XFILLER_240_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_233_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21680_ _08486_ _08487_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__nor2_1
XFILLER_196_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20631_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[5\]\[0\]
+ _07552_ _07550_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_43_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_178_Right_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23350_ _09976_ _09977_ VGND VGND VPWR VPWR _09978_ sky130_fd_sc_hd__nor2_1
X_20562_ systolic_inst.B_outs\[5\]\[6\] systolic_inst.A_outs\[5\]\[7\] VGND VGND VPWR
+ VPWR _07494_ sky130_fd_sc_hd__nand2_1
XFILLER_220_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload7 clknet_5_8__leaf_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__bufinv_16
X_22301_ _09042_ _09043_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23281_ systolic_inst.A_outs\[0\]\[4\] systolic_inst.A_shift\[0\]\[4\] net121 VGND
+ VGND VPWR VPWR _01910_ sky130_fd_sc_hd__mux2_1
XFILLER_192_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20493_ net120 _07427_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__nand2_1
XFILLER_20_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_184_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25020_ net112 ser_C.shift_reg\[338\] VGND VGND VPWR VPWR _10980_ sky130_fd_sc_hd__and2_1
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22232_ _08945_ _08976_ VGND VGND VPWR VPWR _08978_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_184_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22163_ _08891_ _08909_ VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__xnor2_1
XFILLER_191_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_180_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21114_ _07907_ _07910_ _07946_ _07948_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__o31a_1
X_22094_ net122 systolic_inst.B_outs\[2\]\[0\] systolic_inst.A_outs\[2\]\[0\] VGND
+ VGND VPWR VPWR _08847_ sky130_fd_sc_hd__and3_1
X_26971_ clknet_leaf_25_A_in_serial_clk _00769_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28710_ clknet_leaf_325_clk _02508_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[258\]
+ sky130_fd_sc_hd__dfrtp_1
X_21045_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\] systolic_inst.A_outs\[4\]\[5\]
+ systolic_inst.A_outs\[4\]\[6\] VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__and4_1
X_25922_ systolic_inst.acc_wires\[12\]\[14\] C_out\[398\] net18 VGND VGND VPWR VPWR
+ _03224_ sky130_fd_sc_hd__mux2_1
XFILLER_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29690_ clknet_leaf_347_clk _03485_ VGND VGND VPWR VPWR systolic_inst.A_shift\[30\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28641_ clknet_leaf_179_clk _02439_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[189\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25853_ systolic_inst.acc_wires\[10\]\[9\] C_out\[329\] net12 VGND VGND VPWR VPWR
+ _03155_ sky130_fd_sc_hd__mux2_1
XFILLER_28_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24804_ net113 ser_C.shift_reg\[230\] VGND VGND VPWR VPWR _10872_ sky130_fd_sc_hd__and2_1
X_28572_ clknet_leaf_174_clk _02370_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_178_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25784_ systolic_inst.acc_wires\[8\]\[4\] C_out\[260\] net22 VGND VGND VPWR VPWR
+ _03086_ sky130_fd_sc_hd__mux2_1
X_22996_ _09670_ _09671_ VGND VGND VPWR VPWR _09673_ sky130_fd_sc_hd__and2b_1
XFILLER_216_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27523_ clknet_leaf_232_clk _01321_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_24735_ C_out\[194\] net97 net80 ser_C.shift_reg\[194\] _10837_ VGND VGND VPWR VPWR
+ _02444_ sky130_fd_sc_hd__a221o_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21947_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[3\]\[12\]
+ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__or2_1
XFILLER_167_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27454_ clknet_leaf_239_clk _01252_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_21878_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[3\]\[2\]
+ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__nand2_1
X_24666_ net110 ser_C.shift_reg\[161\] VGND VGND VPWR VPWR _10803_ sky130_fd_sc_hd__and2_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26405_ clknet_leaf_30_clk _00212_ net133 VGND VGND VPWR VPWR A_in\[73\] sky130_fd_sc_hd__dfrtp_1
X_23617_ _10201_ _10203_ _10237_ VGND VGND VPWR VPWR _10238_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20829_ systolic_inst.A_outs\[4\]\[2\] systolic_inst.A_shift\[8\]\[2\] net121 VGND
+ VGND VPWR VPWR _01652_ sky130_fd_sc_hd__mux2_1
X_27385_ clknet_leaf_338_clk _01183_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_208_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24597_ C_out\[125\] net99 net80 ser_C.shift_reg\[125\] _10768_ VGND VGND VPWR VPWR
+ _02375_ sky130_fd_sc_hd__a221o_1
X_29124_ clknet_leaf_173_clk _02922_ net148 VGND VGND VPWR VPWR C_out\[96\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26336_ clknet_leaf_58_clk _00143_ net137 VGND VGND VPWR VPWR A_in\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14350_ _11533_ _11534_ VGND VGND VPWR VPWR _11535_ sky130_fd_sc_hd__and2_1
X_23548_ _10152_ _10169_ VGND VGND VPWR VPWR _10171_ sky130_fd_sc_hd__xor2_1
XFILLER_128_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13301_ A_in\[10\] deser_A.word_buffer\[10\] net93 VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__mux2_1
XFILLER_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29055_ clknet_leaf_110_clk _02853_ net151 VGND VGND VPWR VPWR C_out\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14281_ _11436_ _11467_ VGND VGND VPWR VPWR _11468_ sky130_fd_sc_hd__xnor2_1
X_23479_ _10102_ _10103_ net121 VGND VGND VPWR VPWR _10104_ sky130_fd_sc_hd__and3b_1
X_26267_ clknet_leaf_16_A_in_serial_clk _00075_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28006_ clknet_leaf_153_clk _01804_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_16020_ _13016_ _13017_ VGND VGND VPWR VPWR _13018_ sky130_fd_sc_hd__or2_1
X_13232_ deser_A.word_buffer\[70\] deser_A.serial_word\[70\] net127 VGND VGND VPWR
+ VPWR _00080_ sky130_fd_sc_hd__mux2_1
XFILLER_104_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25218_ net110 ser_C.shift_reg\[437\] VGND VGND VPWR VPWR _11079_ sky130_fd_sc_hd__and2_1
XFILLER_104_1382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26198_ systolic_inst.A_shift\[30\]\[4\] net71 _11333_ A_in\[124\] VGND VGND VPWR
+ VPWR _03488_ sky130_fd_sc_hd__a22o_1
XFILLER_108_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13163_ deser_A.word_buffer\[1\] deser_A.serial_word\[1\] net128 VGND VGND VPWR VPWR
+ _00011_ sky130_fd_sc_hd__mux2_1
XFILLER_48_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25149_ C_out\[401\] net101 net73 ser_C.shift_reg\[401\] _11044_ VGND VGND VPWR VPWR
+ _02651_ sky130_fd_sc_hd__a221o_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17971_ _05160_ _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19710_ systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[5\] systolic_inst.A_outs\[6\]\[6\]
+ systolic_inst.B_outs\[6\]\[0\] VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__a22oi_1
X_28908_ clknet_leaf_271_clk _02706_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[456\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_105_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16922_ _04236_ _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__nand2_1
XFILLER_172_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19641_ systolic_inst.A_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[2\] _06646_ VGND
+ VGND VPWR VPWR _06648_ sky130_fd_sc_hd__a21o_1
X_28839_ clknet_leaf_328_clk _02637_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[387\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16853_ systolic_inst.A_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[5\] systolic_inst.B_outs\[11\]\[6\]
+ systolic_inst.B_outs\[11\]\[7\] VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__and4b_1
XFILLER_215_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15804_ _12843_ _12844_ net67 VGND VGND VPWR VPWR _12846_ sky130_fd_sc_hd__o21ai_1
XFILLER_92_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19572_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[25\]
+ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_122_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16784_ systolic_inst.A_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[6\] _11262_ systolic_inst.A_outs\[11\]\[2\]
+ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__o2bb2a_1
X_13996_ deser_B.shift_reg\[30\] deser_B.shift_reg\[31\] net125 VGND VGND VPWR VPWR
+ _00822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18523_ _05623_ _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__xnor2_1
X_15735_ _12714_ _12763_ _12762_ VGND VGND VPWR VPWR _12787_ sky130_fd_sc_hd__o21ba_1
XFILLER_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18454_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[3\]
+ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__and3_1
XFILLER_233_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15666_ systolic_inst.B_outs\[13\]\[5\] systolic_inst.A_outs\[13\]\[7\] VGND VGND
+ VPWR VPWR _12720_ sky130_fd_sc_hd__nand2_1
XFILLER_222_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17405_ _04621_ _04622_ _04624_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__o21a_1
XFILLER_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14617_ _11776_ _11780_ VGND VGND VPWR VPWR _11782_ sky130_fd_sc_hd__nand2b_1
X_18385_ net66 _05540_ _05541_ systolic_inst.acc_wires\[9\]\[28\] net105 VGND VGND
+ VPWR VPWR _01390_ sky130_fd_sc_hd__a32o_1
XFILLER_92_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15597_ systolic_inst.A_outs\[13\]\[4\] systolic_inst.B_outs\[13\]\[6\] _11272_ systolic_inst.A_outs\[13\]\[3\]
+ VGND VGND VPWR VPWR _12653_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_222_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_A_in_serial_clk clknet_2_0__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_28_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17336_ _04562_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__and2b_1
XFILLER_144_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14548_ _11716_ _11717_ _11715_ VGND VGND VPWR VPWR _11723_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17267_ _04498_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__and2b_1
Xclkload102 clknet_leaf_268_clk VGND VGND VPWR VPWR clkload102/X sky130_fd_sc_hd__clkbuf_8
X_14479_ _11593_ _11658_ VGND VGND VPWR VPWR _11660_ sky130_fd_sc_hd__or2_1
Xclkload113 clknet_leaf_251_clk VGND VGND VPWR VPWR clkload113/Y sky130_fd_sc_hd__clkinvlp_4
X_19006_ net66 _06095_ _06096_ systolic_inst.acc_wires\[8\]\[30\] net108 VGND VGND
+ VPWR VPWR _01456_ sky130_fd_sc_hd__a32o_1
XFILLER_162_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload124 clknet_leaf_253_clk VGND VGND VPWR VPWR clkload124/Y sky130_fd_sc_hd__clkinv_2
X_16218_ _03597_ _03600_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__xnor2_1
Xclkload135 clknet_leaf_246_clk VGND VGND VPWR VPWR clkload135/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_155_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17198_ systolic_inst.A_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[1\]
+ systolic_inst.B_outs\[10\]\[0\] VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload146 clknet_leaf_226_clk VGND VGND VPWR VPWR clkload146/Y sky130_fd_sc_hd__clkinv_2
Xclkload157 clknet_leaf_213_clk VGND VGND VPWR VPWR clkload157/Y sky130_fd_sc_hd__clkinv_8
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload168 clknet_leaf_241_clk VGND VGND VPWR VPWR clkload168/X sky130_fd_sc_hd__clkbuf_8
XFILLER_127_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16149_ _03531_ _03532_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__xnor2_1
Xclkload179 clknet_leaf_235_clk VGND VGND VPWR VPWR clkload179/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_226_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_226_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19908_ _06867_ _06869_ _06905_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_239_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19839_ _06799_ _06801_ _06838_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__a21o_1
XFILLER_9_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_235_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_235_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22850_ systolic_inst.A_outs\[1\]\[0\] _09461_ VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__nand2_1
XFILLER_209_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21801_ _08515_ _08573_ _08572_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__a21oi_1
XFILLER_232_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22781_ _09459_ _09460_ _09463_ VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__nand3_2
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24520_ net114 ser_C.shift_reg\[88\] VGND VGND VPWR VPWR _10730_ sky130_fd_sc_hd__and2_1
X_21732_ _08536_ _08537_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24451_ C_out\[52\] _11302_ net81 ser_C.shift_reg\[52\] _10695_ VGND VGND VPWR VPWR
+ _02302_ sky130_fd_sc_hd__a221o_1
X_21663_ _08431_ _08433_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__and2_1
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20614_ _07462_ _07525_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__xnor2_1
X_23402_ _10026_ _10027_ VGND VGND VPWR VPWR _10028_ sky130_fd_sc_hd__nand2_1
X_24382_ net7 ser_C.shift_reg\[19\] VGND VGND VPWR VPWR _10661_ sky130_fd_sc_hd__and2_1
XFILLER_184_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27170_ clknet_leaf_253_clk _00968_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_21594_ _08381_ _08383_ _08382_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__o21ba_1
XFILLER_138_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26121_ deser_B.serial_word\[76\] deser_B.shift_reg\[76\] net55 VGND VGND VPWR VPWR
+ _03423_ sky130_fd_sc_hd__mux2_1
XFILLER_193_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23333_ _09939_ _09961_ VGND VGND VPWR VPWR _09962_ sky130_fd_sc_hd__xor2_1
X_20545_ _07476_ _07477_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__nand2_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_140_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_137_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23264_ net109 systolic_inst.acc_wires\[1\]\[29\] net65 _09907_ VGND VGND VPWR VPWR
+ _01903_ sky130_fd_sc_hd__a22o_1
X_26052_ deser_B.serial_word\[7\] deser_B.shift_reg\[7\] net55 VGND VGND VPWR VPWR
+ _03354_ sky130_fd_sc_hd__mux2_1
XFILLER_165_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20476_ _07409_ _07410_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__nand2_1
XFILLER_152_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22215_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[7\] VGND VGND VPWR
+ VPWR _08961_ sky130_fd_sc_hd__and2b_1
X_25003_ C_out\[328\] net97 net80 ser_C.shift_reg\[328\] _10971_ VGND VGND VPWR VPWR
+ _02578_ sky130_fd_sc_hd__a221o_1
X_23195_ net109 systolic_inst.acc_wires\[1\]\[18\] net65 _09849_ VGND VGND VPWR VPWR
+ _01892_ sky130_fd_sc_hd__a22o_1
XFILLER_133_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22146_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[4\]
+ systolic_inst.A_outs\[2\]\[5\] VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__and4_1
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22077_ _08846_ _08845_ systolic_inst.acc_wires\[3\]\[31\] net106 VGND VGND VPWR
+ VPWR _01777_ sky130_fd_sc_hd__a2bb2o_1
X_26954_ clknet_leaf_27_A_in_serial_clk _00752_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25905_ systolic_inst.acc_wires\[11\]\[29\] C_out\[381\] net40 VGND VGND VPWR VPWR
+ _03207_ sky130_fd_sc_hd__mux2_1
X_21028_ _07899_ _07900_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__nor2_1
X_29673_ clknet_leaf_31_B_in_serial_clk _03468_ net134 VGND VGND VPWR VPWR deser_B.serial_word\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26885_ clknet_leaf_8_A_in_serial_clk _00683_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28624_ clknet_leaf_147_clk _02422_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[172\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13850_ deser_A.serial_word\[11\] deser_A.shift_reg\[11\] net58 VGND VGND VPWR VPWR
+ _00676_ sky130_fd_sc_hd__mux2_1
X_25836_ systolic_inst.acc_wires\[9\]\[24\] C_out\[312\] net13 VGND VGND VPWR VPWR
+ _03138_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_214_Right_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28555_ clknet_leaf_172_clk _02353_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25767_ systolic_inst.acc_wires\[7\]\[19\] C_out\[243\] net44 VGND VGND VPWR VPWR
+ _03069_ sky130_fd_sc_hd__mux2_1
X_13781_ B_in\[88\] deser_B.word_buffer\[88\] net89 VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__mux2_1
XFILLER_204_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22979_ _09655_ VGND VGND VPWR VPWR _09656_ sky130_fd_sc_hd__inv_2
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15520_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] _12577_ VGND
+ VGND VPWR VPWR _12578_ sky130_fd_sc_hd__a21o_1
XFILLER_76_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27506_ clknet_leaf_229_clk _01304_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24718_ net113 ser_C.shift_reg\[187\] VGND VGND VPWR VPWR _10829_ sky130_fd_sc_hd__and2_1
X_28486_ clknet_leaf_114_clk _02284_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25698_ systolic_inst.acc_wires\[5\]\[14\] C_out\[174\] net31 VGND VGND VPWR VPWR
+ _03000_ sky130_fd_sc_hd__mux2_1
XFILLER_31_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15451_ _12509_ _12510_ VGND VGND VPWR VPWR _12511_ sky130_fd_sc_hd__or2_1
X_27437_ clknet_leaf_247_clk _01235_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24649_ C_out\[151\] net104 _10643_ ser_C.shift_reg\[151\] _10794_ VGND VGND VPWR
+ VPWR _02401_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_156_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14402_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[10\] _11585_ net118
+ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__mux2_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18170_ _05291_ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__xnor2_1
X_27368_ clknet_leaf_339_clk _01166_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15382_ _12443_ _12444_ _12439_ VGND VGND VPWR VPWR _12446_ sky130_fd_sc_hd__or3b_1
XFILLER_180_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29107_ clknet_leaf_162_clk _02905_ net150 VGND VGND VPWR VPWR C_out\[79\] sky130_fd_sc_hd__dfrtp_1
X_17121_ _04408_ _04409_ _04410_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14333_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[7\]
+ VGND VGND VPWR VPWR _11518_ sky130_fd_sc_hd__o21ai_1
X_26319_ clknet_leaf_0_A_in_serial_clk _00127_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_141_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_131_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27299_ clknet_leaf_290_clk _01097_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29038_ clknet_leaf_122_clk _02836_ net153 VGND VGND VPWR VPWR C_out\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17052_ _04349_ _04350_ _04351_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14264_ _11447_ _11450_ VGND VGND VPWR VPWR _11451_ sky130_fd_sc_hd__xor2_1
XFILLER_171_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16003_ _13000_ _13001_ VGND VGND VPWR VPWR _13002_ sky130_fd_sc_hd__and2b_1
X_13215_ deser_A.word_buffer\[53\] deser_A.serial_word\[53\] net128 VGND VGND VPWR
+ VPWR _00063_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14195_ _11379_ _11382_ VGND VGND VPWR VPWR _11384_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_111_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13146_ ser_C.bit_idx\[4\] ser_C.bit_idx\[5\] ser_C.bit_idx\[6\] ser_C.bit_idx\[7\]
+ VGND VGND VPWR VPWR _11298_ sky130_fd_sc_hd__and4_1
XFILLER_151_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1038 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17954_ systolic_inst.B_outs\[9\]\[7\] _05111_ _05112_ VGND VGND VPWR VPWR _05147_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_239_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16905_ _04219_ _04220_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_198_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_198_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17885_ systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[5\] systolic_inst.A_outs\[9\]\[6\]
+ systolic_inst.B_outs\[9\]\[0\] VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__a22oi_1
XFILLER_239_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19624_ systolic_inst.B_outs\[5\]\[4\] systolic_inst.B_outs\[1\]\[4\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__mux2_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16836_ _04153_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__nor2_1
XFILLER_65_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19555_ _06586_ _06587_ _06588_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__or3_1
XFILLER_0_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16767_ _04050_ _04051_ _04049_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__a21o_1
X_13979_ deser_B.shift_reg\[13\] deser_B.shift_reg\[14\] net125 VGND VGND VPWR VPWR
+ _00805_ sky130_fd_sc_hd__mux2_1
XFILLER_207_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18506_ systolic_inst.A_outs\[8\]\[1\] systolic_inst.B_outs\[8\]\[5\] systolic_inst.B_outs\[8\]\[6\]
+ systolic_inst.A_outs\[8\]\[0\] VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__a22oi_1
XFILLER_207_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15718_ net115 _12769_ _12770_ VGND VGND VPWR VPWR _12771_ sky130_fd_sc_hd__and3_1
XFILLER_0_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19486_ _06528_ _06529_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__nand2_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16698_ systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[6\] systolic_inst.A_outs\[11\]\[7\]
+ systolic_inst.B_outs\[11\]\[0\] VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__a22o_1
XFILLER_181_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18437_ systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[3\]
+ systolic_inst.B_outs\[8\]\[0\] VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__a22o_1
X_15649_ _12701_ _12702_ VGND VGND VPWR VPWR _12704_ sky130_fd_sc_hd__and2b_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18368_ _05525_ _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__nand2_1
XFILLER_222_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17319_ systolic_inst.A_outs\[10\]\[2\] systolic_inst.B_outs\[10\]\[5\] VGND VGND
+ VPWR VPWR _04577_ sky130_fd_sc_hd__nand2_1
XFILLER_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18299_ _05457_ _05462_ _05463_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_228_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20330_ _07235_ _07267_ _07268_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__o21a_1
XFILLER_135_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20261_ _07201_ _07202_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22000_ _08781_ _08780_ systolic_inst.acc_wires\[3\]\[19\] net109 VGND VGND VPWR
+ VPWR _01765_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20192_ _07156_ _07158_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23951_ _10504_ systolic_inst.B_shift\[10\]\[7\] net70 VGND VGND VPWR VPWR _01993_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_189_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_189_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_84_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22902_ _09580_ _09581_ VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__nand2_1
X_26670_ clknet_leaf_8_B_in_serial_clk _00473_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_23882_ _10467_ _10469_ VGND VGND VPWR VPWR _10470_ sky130_fd_sc_hd__xnor2_1
X_25621_ systolic_inst.acc_wires\[3\]\[1\] C_out\[97\] net48 VGND VGND VPWR VPWR _02923_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22833_ systolic_inst.B_outs\[1\]\[3\] systolic_inst.A_outs\[1\]\[4\] _09491_ _09490_
+ VGND VGND VPWR VPWR _09514_ sky130_fd_sc_hd__a31o_1
XFILLER_232_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28340_ clknet_leaf_319_clk _02138_ VGND VGND VPWR VPWR systolic_inst.A_shift\[25\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25552_ systolic_inst.acc_wires\[0\]\[28\] C_out\[28\] net53 VGND VGND VPWR VPWR
+ _02854_ sky130_fd_sc_hd__mux2_1
XFILLER_129_1422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22764_ _11258_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[5\] _09446_
+ _09447_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__a22o_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24503_ C_out\[78\] net100 net80 ser_C.shift_reg\[78\] _10721_ VGND VGND VPWR VPWR
+ _02328_ sky130_fd_sc_hd__a221o_1
XFILLER_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21715_ systolic_inst.B_outs\[3\]\[5\] systolic_inst.A_outs\[3\]\[5\] VGND VGND VPWR
+ VPWR _08522_ sky130_fd_sc_hd__nand2_1
X_28271_ clknet_leaf_129_clk _02069_ VGND VGND VPWR VPWR systolic_inst.B_shift\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25483_ systolic_inst.cycle_cnt\[16\] _11306_ _11215_ systolic_inst.cycle_cnt\[17\]
+ VGND VGND VPWR VPWR _11219_ sky130_fd_sc_hd__a31o_1
X_22695_ _11258_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _09382_ sky130_fd_sc_hd__and2_1
XFILLER_197_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27222_ clknet_leaf_291_clk _01020_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_213_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24434_ net114 ser_C.shift_reg\[45\] VGND VGND VPWR VPWR _10687_ sky130_fd_sc_hd__and2_1
X_21646_ systolic_inst.A_outs\[3\]\[2\] systolic_inst.B_outs\[3\]\[6\] _11274_ systolic_inst.A_outs\[3\]\[1\]
+ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_169_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27153_ clknet_leaf_277_clk _00951_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_113_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_24365_ C_out\[9\] net104 _10643_ ser_C.shift_reg\[9\] _10652_ VGND VGND VPWR VPWR
+ _02259_ sky130_fd_sc_hd__a221o_1
X_21577_ _08354_ _08387_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__nor2_1
XFILLER_166_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26104_ deser_B.serial_word\[59\] deser_B.shift_reg\[59\] net56 VGND VGND VPWR VPWR
+ _03406_ sky130_fd_sc_hd__mux2_1
X_23316_ systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[4\]
+ systolic_inst.A_outs\[0\]\[0\] VGND VGND VPWR VPWR _09945_ sky130_fd_sc_hd__a22o_1
XFILLER_165_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20528_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[7\] _07433_ _07398_
+ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__a31o_1
XFILLER_138_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27084_ clknet_leaf_31_B_in_serial_clk _00882_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24296_ _10621_ systolic_inst.A_shift\[11\]\[3\] net71 VGND VGND VPWR VPWR _02221_
+ sky130_fd_sc_hd__mux2_1
XFILLER_115_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26035_ systolic_inst.acc_wires\[15\]\[31\] ser_C.parallel_data\[511\] net38 VGND
+ VGND VPWR VPWR _03337_ sky130_fd_sc_hd__mux2_1
X_23247_ net109 systolic_inst.acc_wires\[1\]\[26\] net65 _09893_ VGND VGND VPWR VPWR
+ _01900_ sky130_fd_sc_hd__a22o_1
X_20459_ _07322_ _07393_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__nor2_1
XFILLER_238_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23178_ _09833_ _09834_ VGND VGND VPWR VPWR _09835_ sky130_fd_sc_hd__and2_1
XFILLER_238_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22129_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[3\]
+ VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_160_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27986_ clknet_leaf_145_clk _01784_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14951_ _12031_ _12071_ VGND VGND VPWR VPWR _12072_ sky130_fd_sc_hd__nor2_1
X_26937_ clknet_leaf_21_A_in_serial_clk _00735_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13902_ deser_A.serial_word\[63\] deser_A.shift_reg\[63\] net57 VGND VGND VPWR VPWR
+ _00728_ sky130_fd_sc_hd__mux2_1
X_29656_ clknet_leaf_7_B_in_serial_clk _03451_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_17670_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[10\]\[14\]
+ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__nand2_1
X_26868_ clknet_leaf_14_A_in_serial_clk _00666_ net143 VGND VGND VPWR VPWR deser_A.serial_word\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14882_ _12001_ _12004_ VGND VGND VPWR VPWR _12005_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28607_ clknet_leaf_44_clk _02405_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[155\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16621_ systolic_inst.A_outs\[11\]\[1\] systolic_inst.B_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\]
+ systolic_inst.A_outs\[11\]\[0\] VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__a22o_1
X_13833_ deser_B.bit_idx\[3\] deser_B.bit_idx\[4\] _11323_ VGND VGND VPWR VPWR _11327_
+ sky130_fd_sc_hd__and3_1
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25819_ systolic_inst.acc_wires\[9\]\[7\] C_out\[295\] net15 VGND VGND VPWR VPWR
+ _03121_ sky130_fd_sc_hd__mux2_1
X_29587_ clknet_leaf_11_B_in_serial_clk _03382_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26799_ clknet_leaf_87_clk _00601_ net144 VGND VGND VPWR VPWR B_in\[71\] sky130_fd_sc_hd__dfrtp_1
Xmax_cap40 net42 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_3_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19340_ _06335_ _06339_ _06369_ _06399_ _06368_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__o311a_1
Xmax_cap62 net69 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_104_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28538_ clknet_leaf_158_clk _02336_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16552_ _03888_ _03893_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__nand2_1
Xmax_cap73 net75 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_12
XFILLER_90_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13764_ B_in\[71\] deser_B.word_buffer\[71\] net87 VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__mux2_1
Xmax_cap84 net90 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_8
Xmax_cap95 net96 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_12
X_15503_ _12523_ _12559_ VGND VGND VPWR VPWR _12562_ sky130_fd_sc_hd__xor2_1
X_19271_ _06272_ _06297_ _06296_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__a21boi_1
XFILLER_91_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28469_ clknet_leaf_101_clk _02267_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_204_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16483_ _03842_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13695_ B_in\[2\] deser_B.word_buffer\[2\] net86 VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__mux2_1
XFILLER_43_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18222_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[9\]\[5\]
+ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_117_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15434_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[5\] _12492_ _12493_
+ VGND VGND VPWR VPWR _12495_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ _05307_ _05310_ _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_104_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_168_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15365_ systolic_inst.B_outs\[12\]\[1\] systolic_inst.B_outs\[8\]\[1\] net115 VGND
+ VGND VPWR VPWR _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17104_ _04377_ _04382_ _04387_ _04391_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__or4_1
XFILLER_190_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14316_ _11446_ _11462_ _11461_ VGND VGND VPWR VPWR _11502_ sky130_fd_sc_hd__o21a_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18084_ _05233_ _05235_ _05272_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__nand3_1
XFILLER_116_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15296_ systolic_inst.acc_wires\[14\]\[20\] systolic_inst.acc_wires\[14\]\[21\] systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12388_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_74_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17035_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[11\]\[9\]
+ _04333_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__a21oi_1
XFILLER_144_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14247_ _11401_ _11431_ _11430_ VGND VGND VPWR VPWR _11434_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_223_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14178_ _11366_ _11367_ VGND VGND VPWR VPWR _11368_ sky130_fd_sc_hd__nand2_1
XFILLER_112_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13129_ net126 deser_B.bit_idx\[1\] deser_B.bit_idx\[0\] deser_B.bit_idx\[2\] VGND
+ VGND VPWR VPWR _11283_ sky130_fd_sc_hd__and4_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18986_ _06072_ _06076_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__nor2_1
XFILLER_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17937_ _05123_ _05129_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17868_ _05060_ _05063_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19607_ net62 _06632_ _06633_ systolic_inst.acc_wires\[7\]\[30\] net105 VGND VGND
+ VPWR VPWR _01520_ sky130_fd_sc_hd__a32o_1
XFILLER_113_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_896 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16819_ _04136_ _04137_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_217_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17799_ systolic_inst.B_outs\[8\]\[6\] systolic_inst.B_outs\[4\]\[6\] net121 VGND
+ VGND VPWR VPWR _01344_ sky130_fd_sc_hd__mux2_1
XFILLER_241_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_217_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19538_ _06555_ _06560_ _06565_ _06569_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__or4_1
XFILLER_241_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19469_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[7\]\[9\]
+ _06511_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_343_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_343_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_224_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21500_ _08303_ _08313_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__or2_1
X_22480_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[2\]\[0\]
+ _09209_ _09207_ VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__a31o_1
XFILLER_195_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21431_ systolic_inst.acc_wires\[4\]\[24\] systolic_inst.acc_wires\[4\]\[25\] systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__o21a_1
XFILLER_124_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24150_ _10576_ systolic_inst.A_shift\[28\]\[6\] net71 VGND VGND VPWR VPWR _02120_
+ sky130_fd_sc_hd__mux2_1
X_21362_ _08209_ _08210_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__and2_1
XFILLER_163_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23101_ _09762_ _09763_ _09761_ VGND VGND VPWR VPWR _09769_ sky130_fd_sc_hd__a21bo_1
X_20313_ _07250_ _07251_ net120 VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__o21a_1
XFILLER_107_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24081_ systolic_inst.B_shift\[2\]\[0\] _11332_ net83 systolic_inst.B_shift\[6\]\[0\]
+ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__a22o_1
XFILLER_174_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21293_ _08150_ _08151_ _08143_ _08147_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__a211o_1
XFILLER_190_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23032_ _09707_ VGND VGND VPWR VPWR _09708_ sky130_fd_sc_hd__inv_2
X_20244_ _07187_ _07185_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[1\]
+ net109 VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_235_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27840_ clknet_leaf_205_clk _01638_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20175_ _07123_ _07143_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_206_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27771_ clknet_leaf_183_clk _01569_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_24983_ C_out\[318\] net97 net80 ser_C.shift_reg\[318\] _10961_ VGND VGND VPWR VPWR
+ _02568_ sky130_fd_sc_hd__a221o_1
XFILLER_97_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_202_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29510_ clknet_leaf_264_clk _03308_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_198_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26722_ clknet_leaf_32_B_in_serial_clk _00525_ net134 VGND VGND VPWR VPWR deser_B.word_buffer\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23934_ systolic_inst.A_shift\[3\]\[6\] net72 _11333_ A_in\[30\] VGND VGND VPWR VPWR
+ _01984_ sky130_fd_sc_hd__a22o_1
XFILLER_218_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_198_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29441_ clknet_leaf_332_clk _03239_ net131 VGND VGND VPWR VPWR C_out\[413\] sky130_fd_sc_hd__dfrtp_1
X_26653_ clknet_leaf_23_B_in_serial_clk _00456_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_140_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23865_ _10453_ _10455_ VGND VGND VPWR VPWR _10456_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_194_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25604_ systolic_inst.acc_wires\[2\]\[16\] C_out\[80\] net51 VGND VGND VPWR VPWR
+ _02906_ sky130_fd_sc_hd__mux2_1
X_22816_ _09493_ _09496_ VGND VGND VPWR VPWR _09498_ sky130_fd_sc_hd__xnor2_1
X_29372_ clknet_leaf_233_clk _03170_ net145 VGND VGND VPWR VPWR C_out\[344\] sky130_fd_sc_hd__dfrtp_1
X_26584_ clknet_leaf_29_A_in_serial_clk _00387_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_23796_ net63 _10396_ _10397_ systolic_inst.acc_wires\[0\]\[15\] _11258_ VGND VGND
+ VPWR VPWR _01945_ sky130_fd_sc_hd__a32o_1
XFILLER_60_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28323_ clknet_leaf_347_clk _02121_ VGND VGND VPWR VPWR systolic_inst.A_shift\[28\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25535_ systolic_inst.acc_wires\[0\]\[11\] C_out\[11\] net33 VGND VGND VPWR VPWR
+ _02837_ sky130_fd_sc_hd__mux2_1
XFILLER_198_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22747_ systolic_inst.A_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[2\] systolic_inst.B_outs\[1\]\[3\]
+ systolic_inst.B_outs\[1\]\[4\] VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_334_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_334_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_242_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28254_ clknet_leaf_51_clk _02052_ VGND VGND VPWR VPWR systolic_inst.B_shift\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25466_ _00008_ _11207_ VGND VGND VPWR VPWR _11208_ sky130_fd_sc_hd__nor2_1
XFILLER_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13480_ deser_A.shift_reg\[44\] deser_A.shift_reg\[45\] net130 VGND VGND VPWR VPWR
+ _00317_ sky130_fd_sc_hd__mux2_1
XFILLER_232_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22678_ systolic_inst.A_outs\[1\]\[5\] systolic_inst.A_outs\[0\]\[5\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__mux2_1
XFILLER_139_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27205_ clknet_leaf_260_clk _01003_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24417_ C_out\[35\] _11302_ net81 ser_C.shift_reg\[35\] _10678_ VGND VGND VPWR VPWR
+ _02285_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_11_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21629_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[7\] _08437_
+ _08438_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__a22o_1
XFILLER_185_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28185_ clknet_leaf_17_clk _01983_ VGND VGND VPWR VPWR systolic_inst.A_shift\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25397_ systolic_inst.A_shift\[3\]\[6\] A_in\[22\] net59 VGND VGND VPWR VPWR _11168_
+ sky130_fd_sc_hd__mux2_1
XFILLER_148_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27136_ clknet_leaf_86_clk _00934_ VGND VGND VPWR VPWR systolic_inst.B_shift\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15150_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[14\]\[1\]
+ VGND VGND VPWR VPWR _12263_ sky130_fd_sc_hd__nand2_1
X_24348_ net7 ser_C.shift_reg\[2\] VGND VGND VPWR VPWR _10644_ sky130_fd_sc_hd__and2_1
XFILLER_154_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14101_ systolic_inst.A_shift\[12\]\[1\] net72 _11333_ A_in\[57\] VGND VGND VPWR
+ VPWR _00923_ sky130_fd_sc_hd__a22o_1
XFILLER_181_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27067_ clknet_leaf_9_B_in_serial_clk _00865_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_15081_ _12197_ _12198_ VGND VGND VPWR VPWR _12199_ sky130_fd_sc_hd__nor2_1
X_24279_ systolic_inst.B_shift\[27\]\[3\] B_in\[91\] _00008_ VGND VGND VPWR VPWR _10613_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14032_ deser_B.shift_reg\[66\] deser_B.shift_reg\[67\] net126 VGND VGND VPWR VPWR
+ _00858_ sky130_fd_sc_hd__mux2_1
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26018_ systolic_inst.acc_wires\[15\]\[14\] ser_C.parallel_data\[494\] net37 VGND
+ VGND VPWR VPWR _03320_ sky130_fd_sc_hd__mux2_1
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18840_ _05952_ _05953_ _05946_ _05950_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__a211o_1
XFILLER_79_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18771_ _11259_ systolic_inst.A_outs\[8\]\[7\] _05839_ _05864_ VGND VGND VPWR VPWR
+ _05894_ sky130_fd_sc_hd__o211a_1
X_27969_ clknet_leaf_165_clk _01767_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_15983_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[1\]
+ systolic_inst.A_outs\[12\]\[2\] VGND VGND VPWR VPWR _12983_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_106_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[22\]
+ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__or2_1
X_14934_ _12055_ _12054_ VGND VGND VPWR VPWR _12056_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_106_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__inv_2
XFILLER_110_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1__f_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_2_1__leaf_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
X_29639_ clknet_leaf_28_B_in_serial_clk _03434_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_14865_ net107 _11988_ VGND VGND VPWR VPWR _11989_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_102_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16604_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[2\] _03929_ VGND
+ VGND VPWR VPWR _03931_ sky130_fd_sc_hd__a21o_1
X_13816_ B_in\[123\] deser_B.word_buffer\[123\] net89 VGND VGND VPWR VPWR _00653_
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17584_ _11712_ _04830_ _04831_ systolic_inst.acc_wires\[10\]\[1\] net107 VGND VGND
+ VPWR VPWR _01299_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_11_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14796_ _11900_ _11921_ VGND VGND VPWR VPWR _11922_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_63_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19323_ _06381_ _06382_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16535_ _03887_ _03886_ systolic_inst.acc_wires\[12\]\[24\] net108 VGND VGND VPWR
+ VPWR _01194_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13747_ B_in\[54\] deser_B.word_buffer\[54\] net85 VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__mux2_1
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_325_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_325_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_56_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19254_ _06313_ _06316_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__xnor2_1
X_16466_ net67 _03827_ _03828_ systolic_inst.acc_wires\[12\]\[14\] net108 VGND VGND
+ VPWR VPWR _01184_ sky130_fd_sc_hd__a32o_1
XFILLER_32_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13678_ deser_B.word_buffer\[114\] deser_B.serial_word\[114\] net124 VGND VGND VPWR
+ VPWR _00515_ sky130_fd_sc_hd__mux2_1
XFILLER_31_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18205_ _05378_ _05381_ _05385_ _05386_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__o211a_1
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15417_ _12477_ _12478_ _12461_ VGND VGND VPWR VPWR _12479_ sky130_fd_sc_hd__a21oi_1
X_19185_ systolic_inst.A_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[6\] _11261_ systolic_inst.A_outs\[7\]\[1\]
+ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16397_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18136_ _05322_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__nor2_1
X_15348_ _12430_ _12431_ VGND VGND VPWR VPWR _12432_ sky130_fd_sc_hd__nand2_1
XFILLER_106_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18067_ _05150_ _05256_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_20_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15279_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[20\]
+ VGND VGND VPWR VPWR _12373_ sky130_fd_sc_hd__or2_1
XFILLER_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17018_ _04320_ _04321_ _04322_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_93_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_242_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _06059_ _06061_ _06064_ net61 VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__a31o_1
XFILLER_227_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_219_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_219_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21980_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[16\]
+ VGND VGND VPWR VPWR _08765_ sky130_fd_sc_hd__xnor2_1
XFILLER_226_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20931_ _07803_ _07805_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__or2_1
XFILLER_187_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23650_ _10222_ _10268_ VGND VGND VPWR VPWR _10270_ sky130_fd_sc_hd__and2_1
XFILLER_42_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20862_ systolic_inst.B_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[2\] systolic_inst.B_outs\[4\]\[2\]
+ systolic_inst.A_outs\[4\]\[1\] VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__a22o_1
XFILLER_242_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22601_ _09298_ _09317_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__nor2_1
XFILLER_240_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20793_ _07694_ _07695_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__nand2_1
X_23581_ _10196_ _10202_ VGND VGND VPWR VPWR _10203_ sky130_fd_sc_hd__nor2_1
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_316_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_316_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_223_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25320_ net112 ser_C.shift_reg\[488\] VGND VGND VPWR VPWR _11130_ sky130_fd_sc_hd__and2_1
XFILLER_224_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22532_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[2\]\[10\]
+ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__or2_1
XFILLER_23_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25251_ ser_C.parallel_data\[452\] net102 net74 ser_C.shift_reg\[452\] _11095_ VGND
+ VGND VPWR VPWR _02702_ sky130_fd_sc_hd__a221o_1
X_22463_ _09123_ _09182_ VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24202_ _10586_ systolic_inst.A_shift\[20\]\[0\] net71 VGND VGND VPWR VPWR _02162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21414_ _08233_ _08241_ _08246_ _08251_ VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__nand4_1
X_22394_ _09132_ _09133_ VGND VGND VPWR VPWR _09135_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25182_ net111 ser_C.shift_reg\[419\] VGND VGND VPWR VPWR _11061_ sky130_fd_sc_hd__and2_1
XFILLER_198_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21345_ _08196_ _08194_ systolic_inst.acc_wires\[4\]\[13\] _11258_ VGND VGND VPWR
+ VPWR _01695_ sky130_fd_sc_hd__a2bb2o_1
X_24133_ systolic_inst.A_shift\[30\]\[6\] A_in\[118\] net59 VGND VGND VPWR VPWR _10568_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_208_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24064_ _10549_ systolic_inst.B_shift\[15\]\[3\] net71 VGND VGND VPWR VPWR _02061_
+ sky130_fd_sc_hd__mux2_1
X_28941_ clknet_leaf_256_clk _02739_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[489\]
+ sky130_fd_sc_hd__dfrtp_1
X_21276_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[4\]\[4\]
+ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__and2_1
XFILLER_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23015_ _09658_ _09661_ _09690_ VGND VGND VPWR VPWR _09691_ sky130_fd_sc_hd__o21ai_1
X_20227_ systolic_inst.A_outs\[5\]\[4\] systolic_inst.A_outs\[4\]\[4\] net116 VGND
+ VGND VPWR VPWR _01590_ sky130_fd_sc_hd__mux2_1
X_28872_ clknet_leaf_293_clk _02670_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[420\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27823_ clknet_leaf_218_clk _01621_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20158_ _07129_ _07128_ systolic_inst.acc_wires\[6\]\[21\] net106 VGND VGND VPWR
+ VPWR _01575_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27754_ clknet_leaf_207_clk _01552_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_20089_ net106 systolic_inst.acc_wires\[6\]\[11\] net68 _07070_ VGND VGND VPWR VPWR
+ _01565_ sky130_fd_sc_hd__a22o_1
X_24966_ net111 ser_C.shift_reg\[311\] VGND VGND VPWR VPWR _10953_ sky130_fd_sc_hd__and2_1
XFILLER_40_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26705_ clknet_leaf_8_B_in_serial_clk _00508_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_23917_ _10491_ systolic_inst.B_shift\[18\]\[2\] net71 VGND VGND VPWR VPWR _01972_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27685_ clknet_leaf_198_clk _01483_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24897_ C_out\[275\] net101 net73 ser_C.shift_reg\[275\] _10918_ VGND VGND VPWR VPWR
+ _02525_ sky130_fd_sc_hd__a221o_1
XFILLER_166_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29424_ clknet_leaf_338_clk _03222_ net131 VGND VGND VPWR VPWR C_out\[396\] sky130_fd_sc_hd__dfrtp_1
X_26636_ clknet_leaf_12_B_in_serial_clk _00439_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_14650_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[18\]
+ VGND VGND VPWR VPWR _11810_ sky130_fd_sc_hd__or2_1
X_23848_ systolic_inst.acc_wires\[0\]\[20\] systolic_inst.acc_wires\[0\]\[21\] systolic_inst.acc_wires\[0\]\[22\]
+ systolic_inst.acc_wires\[0\]\[23\] systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _10441_ sky130_fd_sc_hd__o41a_1
XFILLER_60_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13601_ deser_B.word_buffer\[37\] deser_B.serial_word\[37\] net123 VGND VGND VPWR
+ VPWR _00438_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29355_ clknet_leaf_229_clk _03153_ net140 VGND VGND VPWR VPWR C_out\[327\] sky130_fd_sc_hd__dfrtp_1
XFILLER_207_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_307_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_307_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14581_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[15\]\[8\]
+ VGND VGND VPWR VPWR _11751_ sky130_fd_sc_hd__xor2_1
X_26567_ clknet_leaf_23_A_in_serial_clk _00370_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23779_ _10377_ _10381_ VGND VGND VPWR VPWR _10383_ sky130_fd_sc_hd__nand2b_1
XFILLER_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28306_ clknet_leaf_70_clk _02104_ VGND VGND VPWR VPWR systolic_inst.B_shift\[27\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16320_ _03632_ _03669_ _03668_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__a21bo_1
XFILLER_41_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25518_ systolic_inst.cycle_cnt\[30\] _11239_ VGND VGND VPWR VPWR _11241_ sky130_fd_sc_hd__nand2_1
XFILLER_186_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13532_ deser_A.shift_reg\[96\] deser_A.shift_reg\[97\] net129 VGND VGND VPWR VPWR
+ _00369_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29286_ clknet_leaf_323_clk _03084_ net136 VGND VGND VPWR VPWR C_out\[258\] sky130_fd_sc_hd__dfrtp_1
XFILLER_213_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26498_ clknet_leaf_7_A_in_serial_clk _00301_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28237_ clknet_leaf_126_clk _02035_ VGND VGND VPWR VPWR systolic_inst.B_shift\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16251_ systolic_inst.B_outs\[12\]\[5\] systolic_inst.A_outs\[12\]\[6\] VGND VGND
+ VPWR VPWR _03633_ sky130_fd_sc_hd__nand2_1
X_25449_ _00008_ _11196_ VGND VGND VPWR VPWR _11197_ sky130_fd_sc_hd__nor2_1
X_13463_ deser_A.shift_reg\[27\] deser_A.shift_reg\[28\] deser_A.receiving VGND VGND
+ VPWR VPWR _00300_ sky130_fd_sc_hd__mux2_1
X_15202_ net107 systolic_inst.acc_wires\[14\]\[8\] _11712_ _12307_ VGND VGND VPWR
+ VPWR _01050_ sky130_fd_sc_hd__a22o_1
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28168_ clknet_leaf_96_clk _01966_ VGND VGND VPWR VPWR systolic_inst.B_shift\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16182_ systolic_inst.A_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[6\]
+ systolic_inst.B_outs\[12\]\[7\] VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__and4b_1
XFILLER_103_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13394_ A_in\[103\] deser_A.word_buffer\[103\] net96 VGND VGND VPWR VPWR _00242_
+ sky130_fd_sc_hd__mux2_1
X_27119_ clknet_leaf_32_B_in_serial_clk _00917_ net134 VGND VGND VPWR VPWR deser_B.shift_reg\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15133_ _12246_ _12247_ VGND VGND VPWR VPWR _12249_ sky130_fd_sc_hd__xnor2_1
X_28099_ clknet_leaf_110_clk _01897_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_177_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19941_ _06892_ _06908_ _06906_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__o21a_1
X_15064_ systolic_inst.B_outs\[14\]\[5\] systolic_inst.A_outs\[14\]\[7\] _12180_ VGND
+ VGND VPWR VPWR _12182_ sky130_fd_sc_hd__and3_1
XFILLER_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14015_ deser_B.shift_reg\[49\] deser_B.shift_reg\[50\] net125 VGND VGND VPWR VPWR
+ _00841_ sky130_fd_sc_hd__mux2_1
XFILLER_136_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19872_ _06869_ _06870_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__nand2_1
XFILLER_122_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18823_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[8\]\[4\]
+ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__and2_1
XFILLER_228_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15966_ systolic_inst.A_outs\[12\]\[7\] systolic_inst.A_shift\[24\]\[7\] net115 VGND
+ VGND VPWR VPWR _01145_ sky130_fd_sc_hd__mux2_1
X_18754_ _05875_ _05876_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__xor2_1
XFILLER_114_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17705_ _04930_ _04932_ _04929_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14917_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[6\] VGND VGND
+ VPWR VPWR _12039_ sky130_fd_sc_hd__nand2_1
XFILLER_97_1324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15897_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[22\]
+ VGND VGND VPWR VPWR _12925_ sky130_fd_sc_hd__nand2_1
XFILLER_64_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18685_ _05807_ _05810_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14848_ _11970_ _11971_ VGND VGND VPWR VPWR _11972_ sky130_fd_sc_hd__or2_1
X_17636_ _04872_ _04873_ _04875_ systolic_inst.acc_wires\[10\]\[9\] net105 VGND VGND
+ VPWR VPWR _01307_ sky130_fd_sc_hd__a32o_1
XFILLER_90_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17567_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[14\] _04817_ net118
+ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__mux2_1
XFILLER_225_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14779_ _11903_ _11904_ _11893_ VGND VGND VPWR VPWR _11906_ sky130_fd_sc_hd__a21o_1
XFILLER_56_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19306_ _06367_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__inv_2
X_16518_ systolic_inst.acc_wires\[12\]\[20\] systolic_inst.acc_wires\[12\]\[21\] systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__o21a_1
XFILLER_225_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17498_ _04748_ _04749_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19237_ _06269_ _06270_ _06268_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__a21o_1
X_16449_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__inv_2
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19168_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[7\] _06233_ net119
+ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__mux2_1
XFILLER_118_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18119_ _05305_ _05306_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__and2b_1
X_19099_ _06164_ _06165_ net119 VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__o21a_1
XFILLER_160_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21130_ _07923_ _07999_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__xor2_1
XFILLER_117_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21061_ _07931_ _07932_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__and2_1
XFILLER_67_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20012_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] _06998_
+ _07005_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__a22o_1
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24820_ net113 ser_C.shift_reg\[238\] VGND VGND VPWR VPWR _10880_ sky130_fd_sc_hd__and2_1
XFILLER_86_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24751_ C_out\[202\] net97 net80 ser_C.shift_reg\[202\] _10845_ VGND VGND VPWR VPWR
+ _02452_ sky130_fd_sc_hd__a221o_1
XFILLER_95_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21963_ _08742_ _08746_ _08749_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_93_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_215_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23702_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[0\]\[2\]
+ VGND VGND VPWR VPWR _10317_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27470_ clknet_leaf_304_clk _01268_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_20914_ _07756_ _07763_ _07762_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__a21bo_1
XFILLER_242_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24682_ net111 ser_C.shift_reg\[169\] VGND VGND VPWR VPWR _10811_ sky130_fd_sc_hd__and2_1
X_21894_ _08689_ _08690_ _08682_ _08686_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__a211o_1
XFILLER_215_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26421_ clknet_leaf_14_clk _00228_ net133 VGND VGND VPWR VPWR A_in\[89\] sky130_fd_sc_hd__dfrtp_1
XFILLER_199_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23633_ _10251_ _10252_ VGND VGND VPWR VPWR _10254_ sky130_fd_sc_hd__nor2_1
XFILLER_70_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20845_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[1\]
+ systolic_inst.B_outs\[4\]\[1\] VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__and4_1
XFILLER_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29140_ clknet_leaf_168_clk _02938_ net152 VGND VGND VPWR VPWR C_out\[112\] sky130_fd_sc_hd__dfrtp_1
X_26352_ clknet_leaf_19_clk _00159_ net134 VGND VGND VPWR VPWR A_in\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23564_ systolic_inst.B_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[6\] _10025_ VGND
+ VGND VPWR VPWR _10186_ sky130_fd_sc_hd__and3_1
XFILLER_126_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20776_ net68 _07680_ _07681_ systolic_inst.acc_wires\[5\]\[23\] net106 VGND VGND
+ VPWR VPWR _01641_ sky130_fd_sc_hd__a32o_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25303_ ser_C.parallel_data\[478\] net102 net74 ser_C.shift_reg\[478\] _11121_ VGND
+ VGND VPWR VPWR _02728_ sky130_fd_sc_hd__a221o_1
XFILLER_80_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22515_ _09238_ _09239_ _09237_ VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__a21bo_1
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29071_ clknet_leaf_118_clk _02869_ net152 VGND VGND VPWR VPWR C_out\[43\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26283_ clknet_leaf_19_A_in_serial_clk _00091_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23495_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[7\]
+ VGND VGND VPWR VPWR _10119_ sky130_fd_sc_hd__o21ai_1
XFILLER_210_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28022_ clknet_leaf_161_clk _01820_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_202_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25234_ net111 ser_C.shift_reg\[445\] VGND VGND VPWR VPWR _11087_ sky130_fd_sc_hd__and2_1
XFILLER_13_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22446_ _09159_ _09162_ _09184_ VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__a21oi_1
XFILLER_136_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25165_ C_out\[409\] net101 net73 ser_C.shift_reg\[409\] _11052_ VGND VGND VPWR VPWR
+ _02659_ sky130_fd_sc_hd__a221o_1
X_22377_ _09085_ _09088_ _09117_ _09118_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__o22a_1
XFILLER_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24116_ systolic_inst.B_shift\[27\]\[3\] net72 _11333_ B_in\[123\] VGND VGND VPWR
+ VPWR _02101_ sky130_fd_sc_hd__a22o_1
XFILLER_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21328_ _08166_ _08180_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__nand2_1
X_25096_ net113 ser_C.shift_reg\[376\] VGND VGND VPWR VPWR _11018_ sky130_fd_sc_hd__and2_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24047_ systolic_inst.B_shift\[4\]\[3\] B_in\[3\] _00008_ VGND VGND VPWR VPWR _10541_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28924_ clknet_leaf_267_clk _02722_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[472\]
+ sky130_fd_sc_hd__dfrtp_1
X_21259_ _08122_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__inv_2
XFILLER_81_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28855_ clknet_leaf_337_clk _02653_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[403\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_237_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15820_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[13\]\[11\]
+ VGND VGND VPWR VPWR _12859_ sky130_fd_sc_hd__nor2_1
X_27806_ clknet_leaf_218_clk _01604_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_28786_ clknet_leaf_226_clk _02584_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[334\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_237_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25998_ systolic_inst.acc_wires\[14\]\[26\] ser_C.parallel_data\[474\] net24 VGND
+ VGND VPWR VPWR _03300_ sky130_fd_sc_hd__mux2_1
XFILLER_93_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27737_ clknet_leaf_132_clk _01535_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_15751_ net116 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[13\]\[0\]
+ VGND VGND VPWR VPWR _12801_ sky130_fd_sc_hd__a21oi_1
X_24949_ C_out\[301\] net103 net76 ser_C.shift_reg\[301\] _10944_ VGND VGND VPWR VPWR
+ _02551_ sky130_fd_sc_hd__a221o_1
XFILLER_20_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_84_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
X_14702_ net69 _11853_ _11854_ systolic_inst.acc_wires\[15\]\[25\] net105 VGND VGND
+ VPWR VPWR _01003_ sky130_fd_sc_hd__a32o_1
XFILLER_46_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18470_ systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[5\]
+ systolic_inst.B_outs\[8\]\[0\] VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__a22oi_1
X_27668_ clknet_leaf_147_clk _01466_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_15682_ _12682_ _12734_ VGND VGND VPWR VPWR _12736_ sky130_fd_sc_hd__xor2_1
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17421_ systolic_inst.B_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[7\]
+ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__and3_1
X_26619_ clknet_leaf_22_B_in_serial_clk _00422_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_29407_ clknet_leaf_196_clk _03205_ net146 VGND VGND VPWR VPWR C_out\[379\] sky130_fd_sc_hd__dfrtp_1
X_14633_ _11794_ _11795_ VGND VGND VPWR VPWR _11796_ sky130_fd_sc_hd__or2_1
XFILLER_60_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27599_ clknet_leaf_32_clk _01397_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_120_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17352_ _04607_ _04608_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__nor2_1
XFILLER_158_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29338_ clknet_leaf_215_clk _03136_ net149 VGND VGND VPWR VPWR C_out\[310\] sky130_fd_sc_hd__dfrtp_1
X_14564_ _11733_ _11734_ _11735_ VGND VGND VPWR VPWR _11737_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16303_ _03683_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__inv_2
XFILLER_14_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13515_ deser_A.shift_reg\[79\] deser_A.shift_reg\[80\] net129 VGND VGND VPWR VPWR
+ _00352_ sky130_fd_sc_hd__mux2_1
X_29269_ clknet_leaf_194_clk _03067_ net146 VGND VGND VPWR VPWR C_out\[241\] sky130_fd_sc_hd__dfrtp_1
X_17283_ systolic_inst.A_outs\[10\]\[1\] systolic_inst.B_outs\[10\]\[5\] systolic_inst.B_outs\[10\]\[6\]
+ systolic_inst.A_outs\[10\]\[0\] VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__a22oi_1
X_14495_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[13\] _11675_ net118
+ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19022_ systolic_inst.B_outs\[6\]\[3\] systolic_inst.B_outs\[2\]\[3\] net120 VGND
+ VGND VPWR VPWR _01469_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16234_ _03615_ _03616_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__nand2_1
XFILLER_158_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13446_ deser_A.shift_reg\[10\] deser_A.shift_reg\[11\] deser_A.receiving VGND VGND
+ VPWR VPWR _00283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload306 clknet_leaf_116_clk VGND VGND VPWR VPWR clkload306/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_58_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload317 clknet_leaf_112_clk VGND VGND VPWR VPWR clkload317/Y sky130_fd_sc_hd__bufinv_16
Xclkload14 clknet_5_16__leaf_clk VGND VGND VPWR VPWR clkload14/X sky130_fd_sc_hd__clkbuf_8
XFILLER_16_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload25 clknet_5_30__leaf_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__clkinv_8
Xclkload328 clknet_leaf_169_clk VGND VGND VPWR VPWR clkload328/Y sky130_fd_sc_hd__clkinv_2
XFILLER_127_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16165_ _03547_ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__nor2_1
Xclkload36 clknet_leaf_0_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__clkinv_2
Xclkload339 clknet_2_0__leaf_A_in_serial_clk VGND VGND VPWR VPWR clkload339/X sky130_fd_sc_hd__clkbuf_8
XFILLER_115_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload47 clknet_leaf_329_clk VGND VGND VPWR VPWR clkload47/X sky130_fd_sc_hd__clkbuf_4
X_13377_ A_in\[86\] deser_A.word_buffer\[86\] net95 VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__mux2_1
XFILLER_86_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload58 clknet_leaf_323_clk VGND VGND VPWR VPWR clkload58/Y sky130_fd_sc_hd__clkinv_4
XFILLER_103_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload69 clknet_leaf_319_clk VGND VGND VPWR VPWR clkload69/Y sky130_fd_sc_hd__clkinv_2
X_15116_ systolic_inst.B_outs\[14\]\[5\] systolic_inst.B_outs\[14\]\[6\] systolic_inst.A_outs\[14\]\[7\]
+ VGND VGND VPWR VPWR _12232_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_90_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16096_ _13086_ _13090_ VGND VGND VPWR VPWR _13091_ sky130_fd_sc_hd__nor2_1
XFILLER_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19924_ _06782_ _06920_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__or2_1
XFILLER_142_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15047_ _12128_ _12130_ _12165_ VGND VGND VPWR VPWR _12166_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_228_Right_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19855_ _06783_ _06853_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__nor2_1
XFILLER_123_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1058 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18806_ _05925_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__inv_2
X_19786_ _06780_ _06786_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16998_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18737_ _05859_ _05860_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__nor2_1
X_15949_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[30\]
+ VGND VGND VPWR VPWR _12969_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_75_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_237_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_237_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18668_ _05758_ _05727_ _05757_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__or3b_1
XFILLER_224_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_233_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17619_ _11712_ _04859_ _04861_ systolic_inst.acc_wires\[10\]\[6\] net105 VGND VGND
+ VPWR VPWR _01304_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_233_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18599_ _05725_ _05726_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__or2_1
XFILLER_225_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20630_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[5\]\[2\]
+ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20561_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[12\] _07493_ net120
+ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__mux2_1
XFILLER_165_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload8 clknet_5_9__leaf_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinvlp_4
X_22300_ _09043_ _09042_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__nand2b_1
X_20492_ _07387_ _07425_ _07424_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__a21o_1
X_23280_ systolic_inst.A_outs\[0\]\[3\] systolic_inst.A_shift\[0\]\[3\] net121 VGND
+ VGND VPWR VPWR _01909_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_184_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22231_ _08945_ _08976_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__and2b_1
XFILLER_195_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22162_ _08891_ _08909_ VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__nand2b_1
XFILLER_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_180_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21113_ _07983_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22093_ systolic_inst.B_outs\[1\]\[7\] systolic_inst.B_shift\[1\]\[7\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__mux2_1
XFILLER_156_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26970_ clknet_leaf_25_A_in_serial_clk _00768_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_236_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21044_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.A_outs\[4\]\[6\] VGND VGND VPWR
+ VPWR _07916_ sky130_fd_sc_hd__nand2_1
X_25921_ systolic_inst.acc_wires\[12\]\[13\] C_out\[397\] net18 VGND VGND VPWR VPWR
+ _03223_ sky130_fd_sc_hd__mux2_1
XFILLER_160_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28640_ clknet_leaf_179_clk _02438_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[188\]
+ sky130_fd_sc_hd__dfrtp_1
X_25852_ systolic_inst.acc_wires\[10\]\[8\] C_out\[328\] net12 VGND VGND VPWR VPWR
+ _03154_ sky130_fd_sc_hd__mux2_1
XFILLER_219_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24803_ C_out\[228\] net99 net79 ser_C.shift_reg\[228\] _10871_ VGND VGND VPWR VPWR
+ _02478_ sky130_fd_sc_hd__a221o_1
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28571_ clknet_leaf_175_clk _02369_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_178_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25783_ systolic_inst.acc_wires\[8\]\[3\] C_out\[259\] net22 VGND VGND VPWR VPWR
+ _03085_ sky130_fd_sc_hd__mux2_1
XFILLER_216_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22995_ _09671_ _09670_ VGND VGND VPWR VPWR _09672_ sky130_fd_sc_hd__and2b_1
XFILLER_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_83_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27522_ clknet_leaf_232_clk _01320_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_24734_ net112 ser_C.shift_reg\[195\] VGND VGND VPWR VPWR _10837_ sky130_fd_sc_hd__and2_1
XFILLER_76_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21946_ _08706_ _08709_ _08734_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__a21oi_1
XFILLER_227_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27453_ clknet_leaf_241_clk _01251_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_203_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24665_ C_out\[159\] net104 net76 ser_C.shift_reg\[159\] _10802_ VGND VGND VPWR VPWR
+ _02409_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_137_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21877_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[3\]\[2\]
+ VGND VGND VPWR VPWR _08676_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26404_ clknet_leaf_30_clk _00211_ net133 VGND VGND VPWR VPWR A_in\[72\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23616_ _10234_ _10236_ VGND VGND VPWR VPWR _10237_ sky130_fd_sc_hd__xor2_1
X_20828_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.A_shift\[8\]\[1\] net121 VGND
+ VGND VPWR VPWR _01651_ sky130_fd_sc_hd__mux2_1
X_27384_ clknet_leaf_338_clk _01182_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24596_ net113 ser_C.shift_reg\[126\] VGND VGND VPWR VPWR _10768_ sky130_fd_sc_hd__and2_1
XFILLER_204_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29123_ clknet_leaf_164_clk _02921_ net150 VGND VGND VPWR VPWR C_out\[95\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26335_ clknet_leaf_58_clk _00142_ net137 VGND VGND VPWR VPWR A_in\[3\] sky130_fd_sc_hd__dfrtp_1
X_23547_ _10152_ _10169_ VGND VGND VPWR VPWR _10170_ sky130_fd_sc_hd__nor2_1
X_20759_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[21\]
+ VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__xnor2_2
XFILLER_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13300_ A_in\[9\] deser_A.word_buffer\[9\] net93 VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__mux2_1
X_29054_ clknet_leaf_106_clk _02852_ net151 VGND VGND VPWR VPWR C_out\[26\] sky130_fd_sc_hd__dfrtp_1
X_14280_ _11464_ _11465_ VGND VGND VPWR VPWR _11467_ sky130_fd_sc_hd__xnor2_1
X_26266_ clknet_leaf_16_A_in_serial_clk _00074_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_23478_ _10100_ _10101_ _10058_ _10061_ VGND VGND VPWR VPWR _10103_ sky130_fd_sc_hd__a211o_1
XFILLER_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28005_ clknet_leaf_153_clk _01803_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25217_ C_out\[435\] net101 net73 ser_C.shift_reg\[435\] _11078_ VGND VGND VPWR VPWR
+ _02685_ sky130_fd_sc_hd__a221o_1
X_13231_ deser_A.word_buffer\[69\] deser_A.serial_word\[69\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__mux2_1
X_22429_ _09125_ _09139_ _09137_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__o21a_1
XFILLER_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26197_ systolic_inst.A_shift\[30\]\[3\] net71 _11333_ A_in\[123\] VGND VGND VPWR
+ VPWR _03487_ sky130_fd_sc_hd__a22o_1
XFILLER_100_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_15_A_in_serial_clk clknet_2_3__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_15_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_13_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13162_ deser_A.word_buffer\[0\] deser_A.serial_word\[0\] net127 VGND VGND VPWR VPWR
+ _00010_ sky130_fd_sc_hd__mux2_1
XFILLER_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25148_ net110 ser_C.shift_reg\[402\] VGND VGND VPWR VPWR _11044_ sky130_fd_sc_hd__and2_1
XFILLER_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17970_ _05161_ _05162_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__nor2_1
X_25079_ C_out\[366\] net97 net77 ser_C.shift_reg\[366\] _11009_ VGND VGND VPWR VPWR
+ _02616_ sky130_fd_sc_hd__a221o_1
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28907_ clknet_leaf_270_clk _02705_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[455\]
+ sky130_fd_sc_hd__dfrtp_1
X_16921_ _04169_ _04235_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__or2_1
XFILLER_215_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19640_ systolic_inst.A_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[2\] _06646_ VGND
+ VGND VPWR VPWR _06647_ sky130_fd_sc_hd__nand3_1
X_28838_ clknet_leaf_328_clk _02636_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[386\]
+ sky130_fd_sc_hd__dfrtp_1
X_16852_ systolic_inst.B_outs\[11\]\[5\] systolic_inst.A_outs\[11\]\[6\] VGND VGND
+ VPWR VPWR _04170_ sky130_fd_sc_hd__nand2_1
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15803_ _12843_ _12844_ VGND VGND VPWR VPWR _12845_ sky130_fd_sc_hd__and2_1
X_19571_ _06603_ _06602_ systolic_inst.acc_wires\[7\]\[24\] net105 VGND VGND VPWR
+ VPWR _01514_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_122_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16783_ systolic_inst.A_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[6\]
+ systolic_inst.B_outs\[11\]\[7\] VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__and4b_1
X_13995_ deser_B.shift_reg\[29\] deser_B.shift_reg\[30\] net125 VGND VGND VPWR VPWR
+ _00821_ sky130_fd_sc_hd__mux2_1
X_28769_ clknet_leaf_225_clk _02567_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_57_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_122_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15734_ _12714_ _12785_ VGND VGND VPWR VPWR _12786_ sky130_fd_sc_hd__xnor2_1
X_18522_ _05651_ _05652_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__nor2_1
XFILLER_46_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15665_ _12717_ _12718_ VGND VGND VPWR VPWR _12719_ sky130_fd_sc_hd__nor2_1
X_18453_ systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[3\] systolic_inst.A_outs\[8\]\[4\]
+ systolic_inst.B_outs\[8\]\[0\] VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__a22o_1
XFILLER_181_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14616_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[15\]\[12\]
+ _11778_ _11780_ VGND VGND VPWR VPWR _11781_ sky130_fd_sc_hd__a211o_1
X_17404_ _04642_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__xor2_1
X_18384_ _05536_ _05539_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__nand2_1
XFILLER_18_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15596_ systolic_inst.A_outs\[13\]\[3\] systolic_inst.A_outs\[13\]\[4\] systolic_inst.B_outs\[13\]\[6\]
+ systolic_inst.B_outs\[13\]\[7\] VGND VGND VPWR VPWR _12652_ sky130_fd_sc_hd__and4b_1
XFILLER_57_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17335_ _04563_ _04591_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__xnor2_1
X_14547_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[15\]\[3\]
+ VGND VGND VPWR VPWR _11722_ sky130_fd_sc_hd__or2_1
XFILLER_230_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17266_ _04504_ _04524_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__xnor2_1
X_14478_ _11593_ _11658_ VGND VGND VPWR VPWR _11659_ sky130_fd_sc_hd__nand2_1
XFILLER_105_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload103 clknet_leaf_269_clk VGND VGND VPWR VPWR clkload103/Y sky130_fd_sc_hd__inv_6
XFILLER_31_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload114 clknet_leaf_274_clk VGND VGND VPWR VPWR clkload114/Y sky130_fd_sc_hd__clkinv_2
X_16217_ _03598_ _03599_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__nor2_1
X_19005_ _06091_ _06094_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__or2_1
Xclkload125 clknet_leaf_259_clk VGND VGND VPWR VPWR clkload125/X sky130_fd_sc_hd__clkbuf_8
X_13429_ deser_A.bit_idx\[3\] _11312_ _11314_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17197_ _04460_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__inv_2
Xclkload136 clknet_leaf_248_clk VGND VGND VPWR VPWR clkload136/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_77_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload147 clknet_leaf_227_clk VGND VGND VPWR VPWR clkload147/Y sky130_fd_sc_hd__bufinv_16
Xclkload158 clknet_leaf_214_clk VGND VGND VPWR VPWR clkload158/Y sky130_fd_sc_hd__inv_8
XFILLER_115_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16148_ _03532_ _03531_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__nand2b_1
Xclkload169 clknet_leaf_242_clk VGND VGND VPWR VPWR clkload169/Y sky130_fd_sc_hd__inv_4
XFILLER_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_226_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_226_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16079_ _13062_ _13074_ VGND VGND VPWR VPWR _13075_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19907_ _06895_ _06903_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_239_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19838_ _06829_ _06837_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_32_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 A_in_frame_sync VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_235_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19769_ _06768_ _06769_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_3_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_48_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_232_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21800_ _08551_ _08603_ VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__xor2_1
XFILLER_37_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22780_ _09429_ _09461_ _09462_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__o21a_1
XFILLER_25_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21731_ _08537_ _08536_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__nand2b_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24450_ net114 ser_C.shift_reg\[53\] VGND VGND VPWR VPWR _10695_ sky130_fd_sc_hd__and2_1
X_21662_ _08439_ _08469_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__xor2_1
XFILLER_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23401_ systolic_inst.A_outs\[0\]\[2\] systolic_inst.B_outs\[0\]\[5\] _10025_ VGND
+ VGND VPWR VPWR _10027_ sky130_fd_sc_hd__nand3_1
X_20613_ _07465_ _07530_ _07528_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__a21oi_1
XFILLER_240_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24381_ C_out\[17\] net104 _10643_ ser_C.shift_reg\[17\] _10660_ VGND VGND VPWR VPWR
+ _02267_ sky130_fd_sc_hd__a221o_1
X_21593_ _08373_ _08376_ _08378_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__a21oi_1
XFILLER_165_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26120_ deser_B.serial_word\[75\] deser_B.shift_reg\[75\] net55 VGND VGND VPWR VPWR
+ _03422_ sky130_fd_sc_hd__mux2_1
X_23332_ _09959_ _09960_ VGND VGND VPWR VPWR _09961_ sky130_fd_sc_hd__nor2_1
XFILLER_137_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20544_ _07442_ _07444_ _07475_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__nand3_1
XFILLER_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26051_ deser_B.serial_word\[6\] deser_B.shift_reg\[6\] net55 VGND VGND VPWR VPWR
+ _03353_ sky130_fd_sc_hd__mux2_1
X_23263_ _09904_ _09906_ VGND VGND VPWR VPWR _09907_ sky130_fd_sc_hd__xnor2_1
X_20475_ _07400_ _07408_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__or2_1
XFILLER_118_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25002_ net111 ser_C.shift_reg\[329\] VGND VGND VPWR VPWR _10971_ sky130_fd_sc_hd__and2_1
X_22214_ systolic_inst.A_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[5\] VGND VGND VPWR
+ VPWR _08960_ sky130_fd_sc_hd__nand2_1
XFILLER_152_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23194_ _09846_ _09848_ VGND VGND VPWR VPWR _09849_ sky130_fd_sc_hd__xor2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22145_ systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[5\]
+ systolic_inst.B_outs\[2\]\[0\] VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__a22oi_1
XFILLER_105_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22076_ _08840_ _08843_ _08844_ net60 VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__a31o_1
XFILLER_47_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26953_ clknet_leaf_27_A_in_serial_clk _00751_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25904_ systolic_inst.acc_wires\[11\]\[28\] C_out\[380\] net40 VGND VGND VPWR VPWR
+ _03206_ sky130_fd_sc_hd__mux2_1
X_21027_ _07882_ _07898_ VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__and2_1
X_29672_ clknet_leaf_29_B_in_serial_clk _03467_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_26884_ clknet_leaf_9_A_in_serial_clk _00682_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28623_ clknet_leaf_142_clk _02421_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[171\]
+ sky130_fd_sc_hd__dfrtp_1
X_25835_ systolic_inst.acc_wires\[9\]\[23\] C_out\[311\] net13 VGND VGND VPWR VPWR
+ _03137_ sky130_fd_sc_hd__mux2_1
XFILLER_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_210_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28554_ clknet_leaf_172_clk _02352_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_25766_ systolic_inst.acc_wires\[7\]\[18\] C_out\[242\] net44 VGND VGND VPWR VPWR
+ _03068_ sky130_fd_sc_hd__mux2_1
X_13780_ B_in\[87\] deser_B.word_buffer\[87\] net89 VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__mux2_1
X_22978_ _09653_ _09654_ VGND VGND VPWR VPWR _09655_ sky130_fd_sc_hd__nand2_2
XFILLER_142_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24717_ C_out\[185\] net99 net79 ser_C.shift_reg\[185\] _10828_ VGND VGND VPWR VPWR
+ _02435_ sky130_fd_sc_hd__a221o_1
X_27505_ clknet_leaf_228_clk _01303_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_28485_ clknet_leaf_108_clk _02283_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_21929_ _08718_ _08719_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__and2_1
XFILLER_16_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25697_ systolic_inst.acc_wires\[5\]\[13\] C_out\[173\] net31 VGND VGND VPWR VPWR
+ _02999_ sky130_fd_sc_hd__mux2_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15450_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[5\]
+ systolic_inst.A_outs\[13\]\[6\] VGND VGND VPWR VPWR _12510_ sky130_fd_sc_hd__and4_1
X_27436_ clknet_leaf_248_clk _01234_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24648_ net7 ser_C.shift_reg\[152\] VGND VGND VPWR VPWR _10794_ sky130_fd_sc_hd__and2_1
XFILLER_71_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14401_ _11583_ _11584_ VGND VGND VPWR VPWR _11585_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27367_ clknet_leaf_339_clk _01165_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15381_ _12443_ _12444_ VGND VGND VPWR VPWR _12445_ sky130_fd_sc_hd__or2_1
X_24579_ C_out\[116\] net100 net82 ser_C.shift_reg\[116\] _10759_ VGND VGND VPWR VPWR
+ _02366_ sky130_fd_sc_hd__a221o_1
X_17120_ _04409_ _04410_ _04408_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__o21ai_1
X_29106_ clknet_leaf_162_clk _02904_ net150 VGND VGND VPWR VPWR C_out\[78\] sky130_fd_sc_hd__dfrtp_1
XFILLER_180_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26318_ clknet_leaf_29_A_in_serial_clk _00126_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_14332_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[7\]
+ VGND VGND VPWR VPWR _11517_ sky130_fd_sc_hd__o21a_1
XFILLER_204_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27298_ clknet_leaf_290_clk _01096_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_141_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_208_Left_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29037_ clknet_leaf_124_clk _02835_ net153 VGND VGND VPWR VPWR C_out\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17051_ _04349_ _04350_ _04351_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_169_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _11448_ _11449_ VGND VGND VPWR VPWR _11450_ sky130_fd_sc_hd__or2_1
X_26249_ clknet_leaf_11_A_in_serial_clk _00057_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16002_ _12978_ _12985_ _12987_ VGND VGND VPWR VPWR _13001_ sky130_fd_sc_hd__a21bo_1
X_13214_ deser_A.word_buffer\[52\] deser_A.serial_word\[52\] net128 VGND VGND VPWR
+ VPWR _00062_ sky130_fd_sc_hd__mux2_1
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14194_ _11382_ _11379_ VGND VGND VPWR VPWR _11383_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_111_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13145_ _11297_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__inv_2
XFILLER_112_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17953_ _05081_ _05117_ _05115_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__a21o_1
XFILLER_215_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_221_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16904_ _04219_ _04220_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__or2_1
XFILLER_238_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17884_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[3\] _05062_ _05061_
+ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__a31o_1
XFILLER_65_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_217_Left_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19623_ systolic_inst.B_outs\[5\]\[3\] systolic_inst.B_outs\[1\]\[3\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16835_ _04092_ _04119_ _04118_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_109_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19554_ _06587_ _06588_ _06586_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13978_ deser_B.shift_reg\[12\] deser_B.shift_reg\[13\] net125 VGND VGND VPWR VPWR
+ _00804_ sky130_fd_sc_hd__mux2_1
X_16766_ _04084_ _04085_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__xor2_1
XFILLER_207_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18505_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[4\] _05633_ _05634_
+ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__a22o_1
X_15717_ _12739_ _12744_ _12768_ VGND VGND VPWR VPWR _12770_ sky130_fd_sc_hd__o21ai_1
X_19485_ _06529_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__inv_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16697_ _03995_ _03997_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__nand2_1
XFILLER_146_1236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18436_ _05568_ _05569_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__nor2_1
XFILLER_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15648_ _12702_ _12701_ VGND VGND VPWR VPWR _12703_ sky130_fd_sc_hd__and2b_1
XFILLER_194_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18367_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[26\]
+ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__nand2_1
XFILLER_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15579_ _12633_ _12634_ VGND VGND VPWR VPWR _12636_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17318_ _04572_ _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18298_ _05454_ _05459_ _05464_ _05458_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_228_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_228_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17249_ _04508_ _04505_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__nand2b_1
XFILLER_179_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20260_ _07199_ _07200_ _07190_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__a21o_1
XFILLER_31_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20191_ _07149_ _07151_ _07157_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__a21o_1
XFILLER_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23950_ systolic_inst.B_shift\[14\]\[7\] B_in\[23\] net59 VGND VGND VPWR VPWR _10504_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22901_ _09541_ _09543_ _09579_ VGND VGND VPWR VPWR _09581_ sky130_fd_sc_hd__nand3_1
XFILLER_217_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23881_ _10462_ _10465_ _10464_ VGND VGND VPWR VPWR _10469_ sky130_fd_sc_hd__o21a_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25620_ systolic_inst.acc_wires\[3\]\[0\] C_out\[96\] net48 VGND VGND VPWR VPWR _02922_
+ sky130_fd_sc_hd__mux2_1
X_22832_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.A_outs\[1\]\[7\] _09482_ _09481_
+ VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__a31o_1
XFILLER_72_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25551_ systolic_inst.acc_wires\[0\]\[27\] C_out\[27\] net53 VGND VGND VPWR VPWR
+ _02853_ sky130_fd_sc_hd__mux2_1
XFILLER_225_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22763_ _09444_ _09445_ net122 VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__o21a_1
XFILLER_38_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24502_ net113 ser_C.shift_reg\[79\] VGND VGND VPWR VPWR _10721_ sky130_fd_sc_hd__and2_1
XFILLER_13_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21714_ _08485_ _08520_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__xor2_1
X_28270_ clknet_leaf_45_clk _02068_ VGND VGND VPWR VPWR systolic_inst.B_shift\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25482_ systolic_inst.cycle_cnt\[16\] _11217_ _11218_ VGND VGND VPWR VPWR _02810_
+ sky130_fd_sc_hd__o21ai_1
X_22694_ _09381_ _09379_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[1\]
+ _11258_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27221_ clknet_leaf_291_clk _01019_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_213_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24433_ C_out\[43\] _11302_ net81 ser_C.shift_reg\[43\] _10686_ VGND VGND VPWR VPWR
+ _02293_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_213_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21645_ systolic_inst.A_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[2\] systolic_inst.B_outs\[3\]\[6\]
+ systolic_inst.B_outs\[3\]\[7\] VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__and4b_1
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27152_ clknet_leaf_277_clk _00950_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_24364_ net7 ser_C.shift_reg\[10\] VGND VGND VPWR VPWR _10652_ sky130_fd_sc_hd__and2_1
XFILLER_165_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21576_ systolic_inst.A_outs\[3\]\[1\] systolic_inst.B_outs\[3\]\[6\] VGND VGND VPWR
+ VPWR _08387_ sky130_fd_sc_hd__nand2_1
XFILLER_162_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26103_ deser_B.serial_word\[58\] deser_B.shift_reg\[58\] net56 VGND VGND VPWR VPWR
+ _03405_ sky130_fd_sc_hd__mux2_1
X_23315_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[4\] VGND VGND VPWR
+ VPWR _09944_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20527_ _07460_ _07459_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[11\]
+ net109 VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__a2bb2o_1
X_27083_ clknet_leaf_30_B_in_serial_clk _00881_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_24295_ systolic_inst.A_shift\[12\]\[3\] A_in\[51\] net59 VGND VGND VPWR VPWR _10621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_165_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26034_ systolic_inst.acc_wires\[15\]\[30\] ser_C.parallel_data\[510\] net38 VGND
+ VGND VPWR VPWR _03336_ sky130_fd_sc_hd__mux2_1
X_23246_ _09890_ _09892_ VGND VGND VPWR VPWR _09893_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20458_ _07364_ _07365_ _07366_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__o21ba_1
XFILLER_134_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23177_ _09821_ _09828_ _09829_ VGND VGND VPWR VPWR _09834_ sky130_fd_sc_hd__o21ba_1
XFILLER_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20389_ _07321_ _07324_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22128_ systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[3\] systolic_inst.A_outs\[2\]\[4\]
+ systolic_inst.B_outs\[2\]\[0\] VGND VGND VPWR VPWR _08877_ sky130_fd_sc_hd__a22o_1
XFILLER_171_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27985_ clknet_leaf_151_clk _01783_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_160_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14950_ _12037_ _12039_ _12036_ VGND VGND VPWR VPWR _12071_ sky130_fd_sc_hd__o21ba_1
X_22059_ _08825_ _08827_ _08830_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__a21oi_1
XFILLER_212_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26936_ clknet_leaf_21_A_in_serial_clk _00734_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13901_ deser_A.serial_word\[62\] deser_A.shift_reg\[62\] _00002_ VGND VGND VPWR
+ VPWR _00727_ sky130_fd_sc_hd__mux2_1
X_29655_ clknet_leaf_7_B_in_serial_clk _03450_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_169_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14881_ _12002_ _12003_ VGND VGND VPWR VPWR _12004_ sky130_fd_sc_hd__or2_1
X_26867_ clknet_leaf_14_A_in_serial_clk _00665_ net143 VGND VGND VPWR VPWR deser_A.serial_word\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13832_ deser_B.bit_idx\[3\] deser_B.bit_idx\[2\] _11320_ deser_B.bit_idx\[4\] VGND
+ VGND VPWR VPWR _11326_ sky130_fd_sc_hd__a31o_1
X_28606_ clknet_leaf_135_clk _02404_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[154\]
+ sky130_fd_sc_hd__dfrtp_1
X_16620_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.A_outs\[11\]\[1\] systolic_inst.B_outs\[11\]\[3\]
+ systolic_inst.B_outs\[11\]\[4\] VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__nand4_1
XFILLER_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25818_ systolic_inst.acc_wires\[9\]\[6\] C_out\[294\] net14 VGND VGND VPWR VPWR
+ _03120_ sky130_fd_sc_hd__mux2_1
X_26798_ clknet_leaf_87_clk _00600_ net153 VGND VGND VPWR VPWR B_in\[70\] sky130_fd_sc_hd__dfrtp_1
X_29586_ clknet_leaf_11_B_in_serial_clk _03381_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[34\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap30 net32 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_6
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap41 net42 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_3_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap52 net53 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_8
XFILLER_204_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16551_ net61 _03900_ net108 systolic_inst.acc_wires\[12\]\[27\] VGND VGND VPWR VPWR
+ _01197_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_104_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28537_ clknet_leaf_158_clk _02335_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[85\]
+ sky130_fd_sc_hd__dfrtp_1
X_13763_ B_in\[70\] deser_B.word_buffer\[70\] net87 VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__mux2_1
X_25749_ systolic_inst.acc_wires\[7\]\[1\] C_out\[225\] net42 VGND VGND VPWR VPWR
+ _03051_ sky130_fd_sc_hd__mux2_1
Xmax_cap63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_12
XFILLER_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap74 net76 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_12
XFILLER_188_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap85 net88 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_8
Xmax_cap96 _00003_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_8
X_15502_ _12523_ _12559_ VGND VGND VPWR VPWR _12561_ sky130_fd_sc_hd__and2_1
X_19270_ _06331_ _06332_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__nand2_1
X_16482_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[16\]
+ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28468_ clknet_leaf_101_clk _02266_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13694_ B_in\[1\] deser_B.word_buffer\[1\] net88 VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_0__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_75_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15433_ _12492_ _12493_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[5\]
+ VGND VGND VPWR VPWR _12494_ sky130_fd_sc_hd__and4bb_1
X_18221_ net66 _05399_ _05401_ systolic_inst.acc_wires\[9\]\[4\] net107 VGND VGND
+ VPWR VPWR _01366_ sky130_fd_sc_hd__a32o_1
XFILLER_176_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27419_ clknet_leaf_215_clk _01217_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_117_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28399_ clknet_leaf_32_clk _02197_ VGND VGND VPWR VPWR systolic_inst.A_shift\[16\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[8\]\[0\] net115 VGND
+ VGND VPWR VPWR _01082_ sky130_fd_sc_hd__mux2_1
X_18152_ _05290_ _05339_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17103_ _04394_ _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__and2_1
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14315_ _11482_ _11499_ VGND VGND VPWR VPWR _11501_ sky130_fd_sc_hd__xor2_1
XFILLER_102_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18083_ _05233_ _05235_ _05272_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__a21o_1
XFILLER_106_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15295_ _12385_ _12386_ VGND VGND VPWR VPWR _12387_ sky130_fd_sc_hd__and2_1
XFILLER_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17034_ _04335_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__and2_1
X_14246_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[6\] _11433_ net118
+ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__mux2_1
XFILLER_172_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14177_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\]
+ systolic_inst.A_outs\[15\]\[0\] VGND VGND VPWR VPWR _11367_ sky130_fd_sc_hd__a22o_1
XFILLER_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13128_ deser_A.bit_idx\[6\] _11281_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__and2_4
XFILLER_124_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18985_ net108 systolic_inst.acc_wires\[8\]\[27\] net66 _06078_ VGND VGND VPWR VPWR
+ _01453_ sky130_fd_sc_hd__a22o_1
XFILLER_61_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17936_ _05123_ _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__nor2_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17867_ _05061_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_17_B_in_serial_clk clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_17_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_19606_ _06628_ _06631_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16818_ systolic_inst.A_outs\[11\]\[4\] systolic_inst.B_outs\[11\]\[6\] _11262_ systolic_inst.A_outs\[11\]\[3\]
+ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17798_ systolic_inst.B_outs\[8\]\[5\] systolic_inst.B_outs\[4\]\[5\] net121 VGND
+ VGND VPWR VPWR _01343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_217_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19537_ _06572_ _06573_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__and2_1
XFILLER_19_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16749_ _04068_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__and2b_1
XFILLER_98_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19468_ _06513_ _06514_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__and2_1
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18419_ net115 systolic_inst.B_outs\[8\]\[0\] systolic_inst.A_outs\[8\]\[0\] VGND
+ VGND VPWR VPWR _05556_ sky130_fd_sc_hd__and3_1
XFILLER_210_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19399_ _06453_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21430_ _08267_ _08268_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__nand2_1
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21361_ _08198_ _08204_ _08205_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__o21ba_1
XFILLER_238_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23100_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[1\]\[5\]
+ VGND VGND VPWR VPWR _09768_ sky130_fd_sc_hd__or2_1
XFILLER_200_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20312_ _07250_ _07251_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__nand2_1
XFILLER_107_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24080_ systolic_inst.B_shift\[3\]\[7\] _11332_ net83 systolic_inst.B_shift\[7\]\[7\]
+ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__a22o_1
XFILLER_238_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21292_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[4\]\[6\]
+ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__or2_1
XFILLER_200_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23031_ _09672_ _09675_ _09705_ VGND VGND VPWR VPWR _09707_ sky130_fd_sc_hd__nor3_1
XFILLER_116_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20243_ net116 _07186_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20174_ systolic_inst.acc_wires\[6\]\[20\] systolic_inst.acc_wires\[6\]\[21\] systolic_inst.acc_wires\[6\]\[22\]
+ systolic_inst.acc_wires\[6\]\[23\] systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__o41a_1
XFILLER_131_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_206_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_206_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27770_ clknet_leaf_183_clk _01568_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24982_ net111 ser_C.shift_reg\[319\] VGND VGND VPWR VPWR _10961_ sky130_fd_sc_hd__and2_1
XFILLER_44_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26721_ clknet_leaf_31_B_in_serial_clk _00524_ net134 VGND VGND VPWR VPWR deser_B.word_buffer\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_23933_ systolic_inst.A_shift\[3\]\[5\] net72 _11333_ A_in\[29\] VGND VGND VPWR VPWR
+ _01983_ sky130_fd_sc_hd__a22o_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26652_ clknet_leaf_23_B_in_serial_clk _00455_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_29440_ clknet_leaf_332_clk _03238_ net131 VGND VGND VPWR VPWR C_out\[412\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23864_ _10446_ _10448_ _10454_ VGND VGND VPWR VPWR _10455_ sky130_fd_sc_hd__a21o_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25603_ systolic_inst.acc_wires\[2\]\[15\] C_out\[79\] net51 VGND VGND VPWR VPWR
+ _02905_ sky130_fd_sc_hd__mux2_1
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22815_ _09493_ _09496_ VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__nand2_1
X_26583_ clknet_leaf_28_A_in_serial_clk _00386_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_29371_ clknet_leaf_232_clk _03169_ net147 VGND VGND VPWR VPWR C_out\[343\] sky130_fd_sc_hd__dfrtp_1
X_23795_ _10388_ _10393_ _10394_ _10395_ VGND VGND VPWR VPWR _10397_ sky130_fd_sc_hd__a211o_1
XFILLER_38_1103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25534_ systolic_inst.acc_wires\[0\]\[10\] C_out\[10\] net33 VGND VGND VPWR VPWR
+ _02836_ sky130_fd_sc_hd__mux2_1
X_28322_ clknet_leaf_348_clk _02120_ VGND VGND VPWR VPWR systolic_inst.A_shift\[28\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_22746_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[3\] VGND VGND VPWR
+ VPWR _09430_ sky130_fd_sc_hd__nand2_1
XFILLER_164_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28253_ clknet_leaf_51_clk _02051_ VGND VGND VPWR VPWR systolic_inst.B_shift\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25465_ systolic_inst.ce_local _11206_ VGND VGND VPWR VPWR _11207_ sky130_fd_sc_hd__and2_1
XFILLER_201_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22677_ systolic_inst.A_outs\[1\]\[4\] systolic_inst.A_outs\[0\]\[4\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__mux2_1
XFILLER_179_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27204_ clknet_leaf_259_clk _01002_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_24416_ net114 ser_C.shift_reg\[36\] VGND VGND VPWR VPWR _10678_ sky130_fd_sc_hd__and2_1
XFILLER_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21628_ _08397_ _08400_ _08436_ net122 VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__o31a_1
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28184_ clknet_leaf_64_clk _01982_ VGND VGND VPWR VPWR systolic_inst.A_shift\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25396_ _11167_ systolic_inst.A_shift\[2\]\[5\] net71 VGND VGND VPWR VPWR _02775_
+ sky130_fd_sc_hd__mux2_1
XFILLER_225_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27135_ clknet_leaf_86_clk _00933_ VGND VGND VPWR VPWR systolic_inst.B_shift\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_24347_ C_out\[0\] net104 _10643_ ser_C.shift_reg\[0\] _10642_ VGND VGND VPWR VPWR
+ _02250_ sky130_fd_sc_hd__a221o_1
X_21559_ _08339_ _08342_ _08369_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__or3_1
XFILLER_201_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14100_ systolic_inst.A_shift\[12\]\[0\] net71 _11333_ A_in\[56\] VGND VGND VPWR
+ VPWR _00922_ sky130_fd_sc_hd__a22o_1
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27066_ clknet_leaf_8_B_in_serial_clk _00864_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_15080_ _12105_ _12164_ _12162_ VGND VGND VPWR VPWR _12198_ sky130_fd_sc_hd__a21oi_1
XFILLER_165_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24278_ _10612_ systolic_inst.B_shift\[23\]\[2\] net71 VGND VGND VPWR VPWR _02212_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14031_ deser_B.shift_reg\[65\] deser_B.shift_reg\[66\] net126 VGND VGND VPWR VPWR
+ _00857_ sky130_fd_sc_hd__mux2_1
XFILLER_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26017_ systolic_inst.acc_wires\[15\]\[13\] ser_C.parallel_data\[493\] net37 VGND
+ VGND VPWR VPWR _03319_ sky130_fd_sc_hd__mux2_1
X_23229_ systolic_inst.acc_wires\[1\]\[20\] systolic_inst.acc_wires\[1\]\[21\] systolic_inst.acc_wires\[1\]\[22\]
+ systolic_inst.acc_wires\[1\]\[23\] systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09878_ sky130_fd_sc_hd__o41a_1
XFILLER_180_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_270_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_270_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18770_ systolic_inst.B_outs\[8\]\[5\] systolic_inst.B_outs\[8\]\[6\] systolic_inst.A_outs\[8\]\[7\]
+ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__nand3_1
X_27968_ clknet_leaf_165_clk _01766_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_15982_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.A_outs\[12\]\[2\] VGND VGND
+ VPWR VPWR _12982_ sky130_fd_sc_hd__nand2_1
XFILLER_209_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17721_ _04948_ _04947_ systolic_inst.acc_wires\[10\]\[21\] net106 VGND VGND VPWR
+ VPWR _01319_ sky130_fd_sc_hd__a2bb2o_1
X_14933_ _12000_ _12015_ _12014_ VGND VGND VPWR VPWR _12055_ sky130_fd_sc_hd__o21a_1
X_26919_ clknet_leaf_4_A_in_serial_clk _00717_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27899_ clknet_leaf_43_clk _01697_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29638_ clknet_leaf_28_B_in_serial_clk _03433_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _04878_ _04884_ _04885_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__nand3_1
XFILLER_169_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14864_ _11959_ _11985_ _11986_ VGND VGND VPWR VPWR _11988_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_67_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16603_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[2\] _03929_ VGND
+ VGND VPWR VPWR _03930_ sky130_fd_sc_hd__nand3_1
XFILLER_217_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13815_ B_in\[122\] deser_B.word_buffer\[122\] net89 VGND VGND VPWR VPWR _00652_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29569_ clknet_leaf_17_B_in_serial_clk _03364_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14795_ _11902_ _11919_ _11920_ VGND VGND VPWR VPWR _11921_ sky130_fd_sc_hd__a21oi_1
X_17583_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[10\]\[0\]
+ _04827_ _04828_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__a22o_1
XFILLER_189_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19322_ _06382_ _06381_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__nand2b_1
X_13746_ B_in\[53\] deser_B.word_buffer\[53\] net85 VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__mux2_1
X_16534_ _03884_ _03885_ net61 VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a21o_1
XFILLER_1_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19253_ _06314_ _06315_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__nor2_1
XFILLER_182_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13677_ deser_B.word_buffer\[113\] deser_B.serial_word\[113\] net123 VGND VGND VPWR
+ VPWR _00514_ sky130_fd_sc_hd__mux2_1
X_16465_ _03820_ _03822_ _03826_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__a21o_1
XFILLER_31_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18204_ _05385_ _05386_ _05378_ _05381_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__a211o_1
X_15416_ _12475_ _12476_ _12455_ _12458_ VGND VGND VPWR VPWR _12478_ sky130_fd_sc_hd__o211ai_2
X_19184_ systolic_inst.A_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[6\]
+ systolic_inst.B_outs\[7\]\[7\] VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__and4b_1
X_16396_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[12\]\[5\]
+ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__nand2_1
XFILLER_19_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15347_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[30\]
+ VGND VGND VPWR VPWR _12431_ sky130_fd_sc_hd__or2_1
X_18135_ _05320_ _05321_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__nor2_1
XFILLER_145_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15278_ net107 systolic_inst.acc_wires\[14\]\[19\] _11712_ _12372_ VGND VGND VPWR
+ VPWR _01061_ sky130_fd_sc_hd__a22o_1
X_18066_ systolic_inst.A_outs\[9\]\[6\] _05224_ _05225_ _05191_ VGND VGND VPWR VPWR
+ _05256_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14229_ systolic_inst.A_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[5\]
+ systolic_inst.B_outs\[15\]\[6\] VGND VGND VPWR VPWR _11417_ sky130_fd_sc_hd__and4_1
XFILLER_67_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17017_ _04320_ _04321_ _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__a21o_1
XFILLER_171_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_242_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_261_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_261_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ _06059_ _06061_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_52_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_219_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17919_ _05111_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__nand2_1
XFILLER_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18899_ _06002_ _06004_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__or2_1
XFILLER_187_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20930_ systolic_inst.A_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[3\]
+ systolic_inst.B_outs\[4\]\[4\] VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__and4_1
XFILLER_226_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20861_ _07737_ _07738_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__and2_1
XFILLER_241_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22600_ _09299_ _09304_ _09309_ _09313_ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__or4_1
XFILLER_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23580_ _10199_ _10200_ VGND VGND VPWR VPWR _10202_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_18_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20792_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[26\]
+ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22531_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[2\]\[10\]
+ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__nand2_1
XFILLER_210_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25250_ net111 ser_C.shift_reg\[453\] VGND VGND VPWR VPWR _11095_ sky130_fd_sc_hd__and2_1
XFILLER_195_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22462_ _09126_ _09187_ _09185_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24201_ systolic_inst.A_shift\[21\]\[0\] A_in\[80\] net59 VGND VGND VPWR VPWR _10586_
+ sky130_fd_sc_hd__mux2_1
X_21413_ net63 _08253_ _08254_ systolic_inst.acc_wires\[4\]\[23\] _11258_ VGND VGND
+ VPWR VPWR _01705_ sky130_fd_sc_hd__a32o_1
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25181_ C_out\[417\] net103 net75 ser_C.shift_reg\[417\] _11060_ VGND VGND VPWR VPWR
+ _02667_ sky130_fd_sc_hd__a221o_1
X_22393_ _09133_ _09132_ VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__nand2b_1
XFILLER_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24132_ _10567_ systolic_inst.A_shift\[29\]\[5\] net71 VGND VGND VPWR VPWR _02111_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_187_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21344_ _08188_ _08193_ _08195_ net63 VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_187_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_208_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_208_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24063_ systolic_inst.B_shift\[19\]\[3\] B_in\[27\] net59 VGND VGND VPWR VPWR _10549_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28940_ clknet_leaf_256_clk _02738_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[488\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21275_ net63 _08134_ _08136_ systolic_inst.acc_wires\[4\]\[3\] net108 VGND VGND
+ VPWR VPWR _01685_ sky130_fd_sc_hd__a32o_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23014_ _09660_ _09688_ VGND VGND VPWR VPWR _09690_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20226_ systolic_inst.A_outs\[5\]\[3\] systolic_inst.A_outs\[4\]\[3\] net116 VGND
+ VGND VPWR VPWR _01589_ sky130_fd_sc_hd__mux2_1
XFILLER_46_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28871_ clknet_leaf_296_clk _02669_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[419\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_231_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_252_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_252_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27822_ clknet_leaf_218_clk _01620_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20157_ _07119_ _07125_ _07126_ net60 VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__a31o_1
XFILLER_77_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27753_ clknet_leaf_208_clk _01551_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24965_ C_out\[309\] net103 net76 ser_C.shift_reg\[309\] _10952_ VGND VGND VPWR VPWR
+ _02559_ sky130_fd_sc_hd__a221o_1
XFILLER_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20088_ _07068_ _07069_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26704_ clknet_leaf_8_B_in_serial_clk _00507_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_23916_ systolic_inst.B_shift\[22\]\[2\] B_in\[82\] _00008_ VGND VGND VPWR VPWR _10491_
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27684_ clknet_leaf_198_clk _01482_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24896_ net110 ser_C.shift_reg\[276\] VGND VGND VPWR VPWR _10918_ sky130_fd_sc_hd__and2_1
XFILLER_175_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29423_ clknet_leaf_338_clk _03221_ net131 VGND VGND VPWR VPWR C_out\[395\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23847_ _10399_ _10400_ _10420_ _10439_ VGND VGND VPWR VPWR _10440_ sky130_fd_sc_hd__a211o_1
X_26635_ clknet_leaf_12_B_in_serial_clk _00438_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13600_ deser_B.word_buffer\[36\] deser_B.serial_word\[36\] net123 VGND VGND VPWR
+ VPWR _00437_ sky130_fd_sc_hd__mux2_1
XFILLER_14_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _11746_ _11747_ _11745_ VGND VGND VPWR VPWR _11750_ sky130_fd_sc_hd__a21bo_1
X_29354_ clknet_leaf_229_clk _03152_ net140 VGND VGND VPWR VPWR C_out\[326\] sky130_fd_sc_hd__dfrtp_1
XFILLER_214_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23778_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[0\]\[12\]
+ _10379_ _10381_ VGND VGND VPWR VPWR _10382_ sky130_fd_sc_hd__a211o_1
XFILLER_60_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26566_ clknet_leaf_23_A_in_serial_clk _00369_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_220_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28305_ clknet_leaf_69_clk _02103_ VGND VGND VPWR VPWR systolic_inst.B_shift\[27\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13531_ deser_A.shift_reg\[95\] deser_A.shift_reg\[96\] net129 VGND VGND VPWR VPWR
+ _00368_ sky130_fd_sc_hd__mux2_1
X_25517_ _11239_ _11240_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__nor2_1
X_22729_ _09393_ _09411_ _09412_ VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__nor3_1
XFILLER_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26497_ clknet_leaf_7_A_in_serial_clk _00300_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29285_ clknet_leaf_323_clk _03083_ net136 VGND VGND VPWR VPWR C_out\[257\] sky130_fd_sc_hd__dfrtp_1
XFILLER_186_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1094 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16250_ _03560_ _03631_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__xnor2_4
X_25448_ systolic_inst.ce_local _11195_ VGND VGND VPWR VPWR _11196_ sky130_fd_sc_hd__and2_1
X_28236_ clknet_leaf_123_clk _02034_ VGND VGND VPWR VPWR systolic_inst.B_shift\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13462_ deser_A.shift_reg\[26\] deser_A.shift_reg\[27\] deser_A.receiving VGND VGND
+ VPWR VPWR _00299_ sky130_fd_sc_hd__mux2_1
XFILLER_51_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15201_ _12302_ _12306_ VGND VGND VPWR VPWR _12307_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_209_Right_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16181_ systolic_inst.A_outs\[12\]\[4\] systolic_inst.B_outs\[12\]\[5\] VGND VGND
+ VPWR VPWR _03565_ sky130_fd_sc_hd__nand2_1
X_28167_ clknet_leaf_94_clk _01965_ VGND VGND VPWR VPWR systolic_inst.B_shift\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25379_ systolic_inst.B_shift\[18\]\[5\] B_in\[53\] net59 VGND VGND VPWR VPWR _11159_
+ sky130_fd_sc_hd__mux2_1
X_13393_ A_in\[102\] deser_A.word_buffer\[102\] net96 VGND VGND VPWR VPWR _00241_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15132_ _12247_ _12246_ VGND VGND VPWR VPWR _12248_ sky130_fd_sc_hd__and2b_1
X_27118_ clknet_leaf_32_B_in_serial_clk _00916_ net134 VGND VGND VPWR VPWR deser_B.shift_reg\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_28098_ clknet_leaf_109_clk _01896_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_153_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19940_ _06924_ _06936_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__xnor2_1
X_27049_ clknet_leaf_24_B_in_serial_clk _00847_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15063_ systolic_inst.B_outs\[14\]\[5\] systolic_inst.A_outs\[14\]\[7\] VGND VGND
+ VPWR VPWR _12181_ sky130_fd_sc_hd__nand2_1
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14014_ deser_B.shift_reg\[48\] deser_B.shift_reg\[49\] net125 VGND VGND VPWR VPWR
+ _00840_ sky130_fd_sc_hd__mux2_1
XFILLER_135_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19871_ _06860_ _06868_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__or2_1
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_243_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_243_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_214_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18822_ net63 _05937_ _05939_ systolic_inst.acc_wires\[8\]\[3\] net108 VGND VGND
+ VPWR VPWR _01429_ sky130_fd_sc_hd__a32o_1
XFILLER_95_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_158_Left_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18753_ _05875_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__nand2b_1
XFILLER_49_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15965_ systolic_inst.A_outs\[12\]\[6\] systolic_inst.A_shift\[24\]\[6\] net115 VGND
+ VGND VPWR VPWR _01144_ sky130_fd_sc_hd__mux2_1
XFILLER_62_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17704_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[19\]
+ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14916_ _12036_ _12037_ VGND VGND VPWR VPWR _12038_ sky130_fd_sc_hd__nor2_1
X_18684_ _05808_ _05809_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__or2_1
X_15896_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[22\]
+ VGND VGND VPWR VPWR _12924_ sky130_fd_sc_hd__or2_1
XFILLER_97_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17635_ net60 _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__nor2_1
XFILLER_91_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14847_ systolic_inst.B_outs\[14\]\[3\] systolic_inst.A_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\]
+ systolic_inst.A_outs\[14\]\[2\] VGND VGND VPWR VPWR _11971_ sky130_fd_sc_hd__a22oi_1
XFILLER_17_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17566_ _04813_ _04815_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__xor2_1
X_14778_ _11893_ _11903_ _11904_ VGND VGND VPWR VPWR _11905_ sky130_fd_sc_hd__nand3_1
XFILLER_56_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19305_ _06329_ _06331_ _06366_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__and3_1
XFILLER_182_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16517_ _03870_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__and2_1
XFILLER_232_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13729_ B_in\[36\] deser_B.word_buffer\[36\] net90 VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__mux2_1
XFILLER_189_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Left_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17497_ _04749_ _04748_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__nand2b_1
XFILLER_225_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19236_ _06263_ _06265_ _06298_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__nand3_1
XFILLER_149_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16448_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[12\]\[12\]
+ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__nand2_1
XFILLER_165_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19167_ _06231_ _06232_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__xor2_1
XFILLER_121_1323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16379_ _03745_ _03747_ _03750_ _03752_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__o211a_1
XFILLER_121_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18118_ _05306_ _05305_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__and2b_1
XFILLER_173_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19098_ _06164_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__nand2_1
X_18049_ _05237_ _05238_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__xor2_1
XFILLER_236_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21060_ systolic_inst.A_outs\[4\]\[2\] systolic_inst.B_outs\[4\]\[6\] _07891_ _07890_
+ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__a31o_1
XFILLER_235_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20011_ net119 _06994_ _07004_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__and3_1
XFILLER_154_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_234_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_234_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_28_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24750_ net113 ser_C.shift_reg\[203\] VGND VGND VPWR VPWR _10845_ sky130_fd_sc_hd__and2_1
XFILLER_41_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21962_ _08747_ _08748_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__nand2_1
XFILLER_215_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23701_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[0\]\[2\]
+ VGND VGND VPWR VPWR _10316_ sky130_fd_sc_hd__nand2_1
XFILLER_66_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20913_ _07786_ _07787_ _07779_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__a21o_1
X_24681_ C_out\[167\] net103 net76 ser_C.shift_reg\[167\] _10810_ VGND VGND VPWR VPWR
+ _02417_ sky130_fd_sc_hd__a221o_1
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21893_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[3\]\[4\]
+ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__or2_1
XFILLER_82_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23632_ _10178_ _10182_ _10215_ _10217_ _10251_ VGND VGND VPWR VPWR _10253_ sky130_fd_sc_hd__o311a_1
X_26420_ clknet_leaf_13_clk _00227_ net133 VGND VGND VPWR VPWR A_in\[88\] sky130_fd_sc_hd__dfrtp_1
X_20844_ net108 systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[0\] _07724_
+ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__a21o_1
XFILLER_70_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26351_ clknet_leaf_65_clk _00158_ net135 VGND VGND VPWR VPWR A_in\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_126_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23563_ systolic_inst.A_outs\[0\]\[6\] _10154_ _10156_ VGND VGND VPWR VPWR _10185_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_23_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20775_ _07672_ _07676_ _07679_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__a21o_1
XFILLER_204_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_A_in_serial_clk clknet_2_1__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_23_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_167_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25302_ net111 ser_C.shift_reg\[479\] VGND VGND VPWR VPWR _11121_ sky130_fd_sc_hd__and2_1
X_22514_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[2\]\[7\]
+ VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__or2_1
X_29070_ clknet_leaf_118_clk _02868_ net152 VGND VGND VPWR VPWR C_out\[42\] sky130_fd_sc_hd__dfrtp_1
X_26282_ clknet_leaf_19_A_in_serial_clk _00090_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_210_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_189_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23494_ _10114_ _10117_ VGND VGND VPWR VPWR _10118_ sky130_fd_sc_hd__xor2_1
XFILLER_50_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_189_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28021_ clknet_leaf_154_clk _01819_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25233_ ser_C.parallel_data\[443\] net102 net74 ser_C.shift_reg\[443\] _11086_ VGND
+ VGND VPWR VPWR _02693_ sky130_fd_sc_hd__a221o_1
X_22445_ _09182_ _09183_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__nand2_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25164_ net110 ser_C.shift_reg\[410\] VGND VGND VPWR VPWR _11052_ sky130_fd_sc_hd__and2_1
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22376_ _09079_ _09081_ _09115_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24115_ systolic_inst.B_shift\[27\]\[2\] net72 _11333_ B_in\[122\] VGND VGND VPWR
+ VPWR _02100_ sky130_fd_sc_hd__a22o_1
XFILLER_151_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21327_ _08172_ _08177_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__nor2_1
X_25095_ C_out\[374\] net98 net78 ser_C.shift_reg\[374\] _11017_ VGND VGND VPWR VPWR
+ _02624_ sky130_fd_sc_hd__a221o_1
XFILLER_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24046_ _10540_ systolic_inst.B_shift\[0\]\[2\] _11332_ VGND VGND VPWR VPWR _02052_
+ sky130_fd_sc_hd__mux2_1
X_28923_ clknet_leaf_268_clk _02721_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[471\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21258_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[4\]\[0\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__and4_1
XFILLER_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_225_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_225_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20209_ _07170_ _07172_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28854_ clknet_leaf_345_clk _02652_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[402\]
+ sky130_fd_sc_hd__dfrtp_1
X_21189_ _08055_ _08056_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__nor2_1
XFILLER_77_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27805_ clknet_leaf_139_clk _01603_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28785_ clknet_leaf_231_clk _02583_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[333\]
+ sky130_fd_sc_hd__dfrtp_1
X_25997_ systolic_inst.acc_wires\[14\]\[25\] ser_C.parallel_data\[473\] net25 VGND
+ VGND VPWR VPWR _03299_ sky130_fd_sc_hd__mux2_1
X_27736_ clknet_leaf_132_clk _01534_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15750_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[13\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _12800_ sky130_fd_sc_hd__a21o_1
X_24948_ net111 ser_C.shift_reg\[302\] VGND VGND VPWR VPWR _10944_ sky130_fd_sc_hd__and2_1
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14701_ _11847_ _11850_ _11852_ VGND VGND VPWR VPWR _11854_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27667_ clknet_leaf_204_clk _01465_ net147 VGND VGND VPWR VPWR systolic_inst.A_outs\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_15681_ _12682_ _12734_ VGND VGND VPWR VPWR _12735_ sky130_fd_sc_hd__and2b_1
XFILLER_205_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24879_ C_out\[266\] net101 net73 ser_C.shift_reg\[266\] _10909_ VGND VGND VPWR VPWR
+ _02516_ sky130_fd_sc_hd__a221o_1
XFILLER_234_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29406_ clknet_leaf_194_clk _03204_ net146 VGND VGND VPWR VPWR C_out\[378\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17420_ systolic_inst.B_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[6\] systolic_inst.A_outs\[10\]\[7\]
+ systolic_inst.B_outs\[10\]\[3\] VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a22o_1
X_26618_ clknet_leaf_21_B_in_serial_clk _00421_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14632_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[15\]
+ VGND VGND VPWR VPWR _11795_ sky130_fd_sc_hd__and2_1
XFILLER_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27598_ clknet_leaf_33_clk _01396_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_199_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29337_ clknet_leaf_215_clk _03135_ net149 VGND VGND VPWR VPWR C_out\[309\] sky130_fd_sc_hd__dfrtp_1
XFILLER_18_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14563_ _11733_ _11734_ _11735_ VGND VGND VPWR VPWR _11736_ sky130_fd_sc_hd__a21o_1
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17351_ systolic_inst.B_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[5\]
+ systolic_inst.B_outs\[10\]\[3\] VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_81_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26549_ clknet_leaf_19_A_in_serial_clk _00352_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_220_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16302_ _03681_ _03682_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__nor2_1
X_13514_ deser_A.shift_reg\[78\] deser_A.shift_reg\[79\] net129 VGND VGND VPWR VPWR
+ _00351_ sky130_fd_sc_hd__mux2_1
X_29268_ clknet_leaf_194_clk _03066_ net146 VGND VGND VPWR VPWR C_out\[240\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14494_ _11673_ _11674_ VGND VGND VPWR VPWR _11675_ sky130_fd_sc_hd__xnor2_1
X_17282_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[4\] _04538_ _04539_
+ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__a22o_1
X_19021_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.B_outs\[2\]\[2\] net119 VGND
+ VGND VPWR VPWR _01468_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28219_ clknet_leaf_81_clk _02017_ VGND VGND VPWR VPWR systolic_inst.B_shift\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13445_ deser_A.shift_reg\[9\] deser_A.shift_reg\[10\] deser_A.receiving VGND VGND
+ VPWR VPWR _00282_ sky130_fd_sc_hd__mux2_1
X_16233_ _03557_ _03614_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29199_ clknet_leaf_142_clk _02997_ net149 VGND VGND VPWR VPWR C_out\[171\] sky130_fd_sc_hd__dfrtp_1
Xclkload307 clknet_leaf_117_clk VGND VGND VPWR VPWR clkload307/Y sky130_fd_sc_hd__bufinv_16
XFILLER_186_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload318 clknet_leaf_113_clk VGND VGND VPWR VPWR clkload318/Y sky130_fd_sc_hd__clkinv_4
Xclkload15 clknet_5_17__leaf_clk VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload26 clknet_5_31__leaf_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinv_8
Xclkload329 clknet_leaf_173_clk VGND VGND VPWR VPWR clkload329/Y sky130_fd_sc_hd__inv_6
XFILLER_139_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16164_ _03545_ _03546_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__and2_1
Xclkload37 clknet_leaf_320_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__clkinv_4
X_13376_ A_in\[85\] deser_A.word_buffer\[85\] net95 VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload48 clknet_leaf_330_clk VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__clkinv_2
Xclkload59 clknet_leaf_324_clk VGND VGND VPWR VPWR clkload59/Y sky130_fd_sc_hd__inv_8
XFILLER_115_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15115_ systolic_inst.B_outs\[14\]\[5\] systolic_inst.A_outs\[14\]\[7\] _12209_ _12208_
+ VGND VGND VPWR VPWR _12231_ sky130_fd_sc_hd__a31o_1
X_16095_ _11260_ _13089_ VGND VGND VPWR VPWR _13090_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_90_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_192_Right_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19923_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[7\] _06893_ _06858_
+ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__a31o_1
X_15046_ _12105_ _12164_ VGND VGND VPWR VPWR _12165_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_216_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_216_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19854_ _06825_ _06826_ _06827_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__o21ba_1
XFILLER_218_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18805_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[8\]\[0\]
+ _05923_ _05924_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__and4_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19785_ _06781_ _06784_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16997_ _04302_ _04303_ _04304_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__and3_1
XFILLER_84_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18736_ _05792_ _05797_ _05827_ _05859_ _05825_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_88_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ _12958_ _12961_ _12964_ _12967_ VGND VGND VPWR VPWR _12968_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_88_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_237_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_237_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18667_ _05792_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__or2_1
XFILLER_110_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15879_ _12905_ _12907_ _12904_ VGND VGND VPWR VPWR _12910_ sky130_fd_sc_hd__o21ai_1
XFILLER_97_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17618_ _04860_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__inv_2
XFILLER_97_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_233_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18598_ _05725_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__nand2_1
XFILLER_240_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17549_ _04714_ _04798_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__nand2_1
XFILLER_36_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20560_ _07491_ _07492_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__nor2_1
XFILLER_165_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload9 clknet_5_10__leaf_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__clkinvlp_4
X_19219_ systolic_inst.A_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[6\]
+ systolic_inst.B_outs\[7\]\[7\] VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__and4b_1
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20491_ _07387_ _07424_ _07425_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__and3_1
XFILLER_121_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22230_ _08946_ _08974_ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_184_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22161_ _08884_ _08907_ VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__xor2_1
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21112_ _07980_ _07981_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_7_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22092_ systolic_inst.B_outs\[1\]\[6\] systolic_inst.B_shift\[1\]\[6\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__mux2_1
XFILLER_160_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_207_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_207_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21043_ _07914_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__inv_2
X_25920_ systolic_inst.acc_wires\[12\]\[12\] C_out\[396\] net18 VGND VGND VPWR VPWR
+ _03222_ sky130_fd_sc_hd__mux2_1
XFILLER_115_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25851_ systolic_inst.acc_wires\[10\]\[7\] C_out\[327\] net12 VGND VGND VPWR VPWR
+ _03153_ sky130_fd_sc_hd__mux2_1
X_24802_ net113 ser_C.shift_reg\[229\] VGND VGND VPWR VPWR _10871_ sky130_fd_sc_hd__and2_1
XFILLER_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28570_ clknet_leaf_175_clk _02368_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_234_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22994_ _09624_ _09640_ _09638_ VGND VGND VPWR VPWR _09671_ sky130_fd_sc_hd__o21a_1
X_25782_ systolic_inst.acc_wires\[8\]\[2\] C_out\[258\] net22 VGND VGND VPWR VPWR
+ _03084_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27521_ clknet_leaf_232_clk _01319_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21945_ _08710_ _08713_ _08714_ _08732_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__or4b_1
X_24733_ C_out\[193\] net100 net80 ser_C.shift_reg\[193\] _10836_ VGND VGND VPWR VPWR
+ _02443_ sky130_fd_sc_hd__a221o_1
XFILLER_215_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24664_ net7 ser_C.shift_reg\[160\] VGND VGND VPWR VPWR _10802_ sky130_fd_sc_hd__and2_1
XFILLER_70_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27452_ clknet_leaf_239_clk _01250_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_242_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21876_ net68 _08674_ _08675_ systolic_inst.acc_wires\[3\]\[1\] net106 VGND VGND
+ VPWR VPWR _01747_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_137_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23615_ systolic_inst.A_outs\[0\]\[6\] _10195_ _10235_ VGND VGND VPWR VPWR _10236_
+ sky130_fd_sc_hd__a21o_1
X_26403_ clknet_leaf_31_clk _00210_ net133 VGND VGND VPWR VPWR A_in\[71\] sky130_fd_sc_hd__dfrtp_1
X_20827_ systolic_inst.A_outs\[4\]\[0\] systolic_inst.A_shift\[8\]\[0\] net121 VGND
+ VGND VPWR VPWR _01650_ sky130_fd_sc_hd__mux2_1
XFILLER_208_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24595_ C_out\[124\] net99 net80 ser_C.shift_reg\[124\] _10767_ VGND VGND VPWR VPWR
+ _02374_ sky130_fd_sc_hd__a221o_1
X_27383_ clknet_leaf_339_clk _01181_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29122_ clknet_leaf_164_clk _02920_ net150 VGND VGND VPWR VPWR C_out\[94\] sky130_fd_sc_hd__dfrtp_1
X_23546_ _10167_ _10168_ VGND VGND VPWR VPWR _10169_ sky130_fd_sc_hd__or2_1
X_26334_ clknet_leaf_59_clk _00141_ net137 VGND VGND VPWR VPWR A_in\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20758_ net68 _07665_ _07666_ systolic_inst.acc_wires\[5\]\[20\] net106 VGND VGND
+ VPWR VPWR _01638_ sky130_fd_sc_hd__a32o_1
XFILLER_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29053_ clknet_leaf_106_clk _02851_ net151 VGND VGND VPWR VPWR C_out\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_196_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26265_ clknet_leaf_3_A_in_serial_clk _00073_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_210_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23477_ _10058_ _10061_ _10100_ _10101_ VGND VGND VPWR VPWR _10102_ sky130_fd_sc_hd__o211a_1
XFILLER_17_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20689_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[5\]\[11\]
+ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__nor2_1
XFILLER_149_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28004_ clknet_leaf_153_clk _01802_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25216_ net110 ser_C.shift_reg\[436\] VGND VGND VPWR VPWR _11078_ sky130_fd_sc_hd__and2_1
X_13230_ deser_A.word_buffer\[68\] deser_A.serial_word\[68\] net127 VGND VGND VPWR
+ VPWR _00078_ sky130_fd_sc_hd__mux2_1
X_22428_ _09126_ _09167_ VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26196_ systolic_inst.A_shift\[30\]\[2\] net71 _11333_ A_in\[122\] VGND VGND VPWR
+ VPWR _03486_ sky130_fd_sc_hd__a22o_1
XFILLER_164_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13161_ _00000_ _11307_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__nor2_1
XFILLER_124_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25147_ C_out\[400\] net101 net73 ser_C.shift_reg\[400\] _11043_ VGND VGND VPWR VPWR
+ _02650_ sky130_fd_sc_hd__a221o_1
X_22359_ _09097_ _09100_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__xor2_1
XFILLER_87_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25078_ net112 ser_C.shift_reg\[367\] VGND VGND VPWR VPWR _11009_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_167_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24029_ systolic_inst.B_shift\[8\]\[2\] B_in\[34\] _00008_ VGND VGND VPWR VPWR _10532_
+ sky130_fd_sc_hd__mux2_1
X_28906_ clknet_leaf_271_clk _02704_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[454\]
+ sky130_fd_sc_hd__dfrtp_1
X_16920_ _04169_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__nand2_1
XFILLER_172_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1092 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28837_ clknet_leaf_329_clk _02635_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[385\]
+ sky130_fd_sc_hd__dfrtp_1
X_16851_ _04097_ _04168_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__xnor2_4
XFILLER_120_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15802_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[13\]\[8\]
+ VGND VGND VPWR VPWR _12844_ sky130_fd_sc_hd__xor2_1
X_19570_ _06596_ _06598_ _06601_ net60 VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__a31o_1
XFILLER_93_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28768_ clknet_leaf_212_clk _02566_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[316\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16782_ systolic_inst.A_outs\[11\]\[4\] systolic_inst.B_outs\[11\]\[5\] VGND VGND
+ VPWR VPWR _04102_ sky130_fd_sc_hd__nand2_1
X_13994_ deser_B.shift_reg\[28\] deser_B.shift_reg\[29\] net125 VGND VGND VPWR VPWR
+ _00820_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18521_ _05649_ _05650_ _05617_ _05619_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__o211a_1
XFILLER_74_951 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27719_ clknet_leaf_187_clk _01517_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_15733_ _12783_ _12784_ VGND VGND VPWR VPWR _12785_ sky130_fd_sc_hd__nor2_1
XFILLER_80_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28699_ clknet_leaf_189_clk _02497_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18452_ _05581_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__xnor2_1
XFILLER_234_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15664_ systolic_inst.A_outs\[13\]\[5\] systolic_inst.B_outs\[13\]\[6\] systolic_inst.A_outs\[13\]\[6\]
+ systolic_inst.B_outs\[13\]\[7\] VGND VGND VPWR VPWR _12718_ sky130_fd_sc_hd__and4b_1
XFILLER_146_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17403_ _04657_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__nand2_1
X_14615_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[15\]\[13\]
+ VGND VGND VPWR VPWR _11780_ sky130_fd_sc_hd__xor2_1
X_18383_ _05536_ _05539_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__or2_1
X_15595_ systolic_inst.B_outs\[13\]\[5\] systolic_inst.A_outs\[13\]\[5\] VGND VGND
+ VPWR VPWR _12651_ sky130_fd_sc_hd__nand2_1
XFILLER_159_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17334_ _04563_ _04591_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__and2b_1
XFILLER_222_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14546_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[15\]\[3\]
+ VGND VGND VPWR VPWR _11721_ sky130_fd_sc_hd__nand2_1
XFILLER_230_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17265_ _04504_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__nand2b_1
XFILLER_197_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14477_ _11655_ _11656_ VGND VGND VPWR VPWR _11658_ sky130_fd_sc_hd__xnor2_1
Xclkload104 clknet_leaf_270_clk VGND VGND VPWR VPWR clkload104/Y sky130_fd_sc_hd__inv_8
X_19004_ _06091_ _06094_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__nand2_1
X_16216_ systolic_inst.A_outs\[12\]\[4\] systolic_inst.B_outs\[12\]\[6\] _11260_ systolic_inst.A_outs\[12\]\[3\]
+ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__o2bb2a_1
Xclkload115 clknet_leaf_275_clk VGND VGND VPWR VPWR clkload115/Y sky130_fd_sc_hd__bufinv_16
X_13428_ deser_A.bit_idx\[3\] _11312_ _11310_ VGND VGND VPWR VPWR _11314_ sky130_fd_sc_hd__o21ai_1
Xclkload126 clknet_leaf_260_clk VGND VGND VPWR VPWR clkload126/X sky130_fd_sc_hd__clkbuf_4
X_17196_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.A_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\]
+ systolic_inst.A_outs\[10\]\[1\] VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__and4_1
Xclkload137 clknet_leaf_250_clk VGND VGND VPWR VPWR clkload137/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload148 clknet_leaf_231_clk VGND VGND VPWR VPWR clkload148/X sky130_fd_sc_hd__clkbuf_4
Xclkload159 clknet_leaf_216_clk VGND VGND VPWR VPWR clkload159/Y sky130_fd_sc_hd__clkinv_8
X_16147_ systolic_inst.A_outs\[12\]\[2\] systolic_inst.B_outs\[12\]\[5\] _03494_ _03493_
+ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__a31oi_1
X_13359_ A_in\[68\] deser_A.word_buffer\[68\] net96 VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16078_ _13041_ _13073_ VGND VGND VPWR VPWR _13074_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19906_ _06895_ _06903_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15029_ systolic_inst.A_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[5\] systolic_inst.B_outs\[14\]\[6\]
+ systolic_inst.B_outs\[14\]\[7\] VGND VGND VPWR VPWR _12148_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_36_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19837_ _06834_ _06835_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19768_ _06769_ _06768_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__nand2b_1
Xinput2 A_in_serial_data VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_216_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18719_ _05806_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__xnor2_1
XFILLER_232_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19699_ _06692_ _06700_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__xor2_1
XFILLER_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21730_ _08484_ _08501_ _08499_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__o21a_1
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21661_ _08469_ _08439_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__nand2b_1
XFILLER_240_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23400_ systolic_inst.A_outs\[0\]\[2\] systolic_inst.B_outs\[0\]\[5\] _10025_ VGND
+ VGND VPWR VPWR _10026_ sky130_fd_sc_hd__a21o_1
X_20612_ _07323_ _07461_ _07535_ _07533_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__a31o_1
X_24380_ net7 ser_C.shift_reg\[18\] VGND VGND VPWR VPWR _10660_ sky130_fd_sc_hd__and2_1
XFILLER_127_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21592_ _08363_ _08393_ _08395_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__o21ba_1
XFILLER_177_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23331_ _09957_ _09958_ _09937_ VGND VGND VPWR VPWR _09960_ sky130_fd_sc_hd__a21oi_1
X_20543_ _07442_ _07444_ _07475_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__a21o_1
XFILLER_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26050_ deser_B.serial_word\[5\] deser_B.shift_reg\[5\] net55 VGND VGND VPWR VPWR
+ _03352_ sky130_fd_sc_hd__mux2_1
X_23262_ _09899_ _09902_ _09901_ VGND VGND VPWR VPWR _09906_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_211_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20474_ _07400_ _07408_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_104_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25001_ C_out\[327\] net97 net80 ser_C.shift_reg\[327\] _10970_ VGND VGND VPWR VPWR
+ _02577_ sky130_fd_sc_hd__a221o_1
X_22213_ _08955_ _08958_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23193_ _09838_ _09840_ _09847_ VGND VGND VPWR VPWR _09848_ sky130_fd_sc_hd__a21oi_1
XFILLER_180_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22144_ _08872_ _08874_ _08873_ VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__a21bo_1
XFILLER_133_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22075_ _08840_ _08843_ _08844_ VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__a21oi_1
X_26952_ clknet_leaf_27_A_in_serial_clk _00750_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25903_ systolic_inst.acc_wires\[11\]\[27\] C_out\[379\] net42 VGND VGND VPWR VPWR
+ _03205_ sky130_fd_sc_hd__mux2_1
X_21026_ _07882_ _07898_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_162_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29671_ clknet_leaf_29_B_in_serial_clk _03466_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_26883_ clknet_leaf_9_A_in_serial_clk _00681_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28622_ clknet_leaf_141_clk _02420_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_1399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25834_ systolic_inst.acc_wires\[9\]\[22\] C_out\[310\] net13 VGND VGND VPWR VPWR
+ _03136_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_113_Left_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28553_ clknet_leaf_172_clk _02351_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_22977_ _09516_ _09652_ VGND VGND VPWR VPWR _09654_ sky130_fd_sc_hd__nand2_2
X_25765_ systolic_inst.acc_wires\[7\]\[17\] C_out\[241\] net41 VGND VGND VPWR VPWR
+ _03067_ sky130_fd_sc_hd__mux2_1
XFILLER_16_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27504_ clknet_leaf_228_clk _01302_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24716_ net113 ser_C.shift_reg\[186\] VGND VGND VPWR VPWR _10828_ sky130_fd_sc_hd__and2_1
X_28484_ clknet_leaf_108_clk _02282_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_21928_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[3\]\[10\]
+ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__or2_1
XFILLER_167_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25696_ systolic_inst.acc_wires\[5\]\[12\] C_out\[172\] net31 VGND VGND VPWR VPWR
+ _02998_ sky130_fd_sc_hd__mux2_1
XFILLER_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27435_ clknet_leaf_235_clk _01233_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_21859_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[14\] _08661_ net122
+ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__mux2_1
X_24647_ C_out\[150\] net104 net76 ser_C.shift_reg\[150\] _10793_ VGND VGND VPWR VPWR
+ _02400_ sky130_fd_sc_hd__a221o_1
XFILLER_54_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14400_ _11580_ _11581_ _11582_ VGND VGND VPWR VPWR _11584_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_156_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27366_ clknet_leaf_339_clk _01164_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15380_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[1\]
+ systolic_inst.A_outs\[13\]\[2\] VGND VGND VPWR VPWR _12444_ sky130_fd_sc_hd__and4_1
X_24578_ net114 ser_C.shift_reg\[117\] VGND VGND VPWR VPWR _10759_ sky130_fd_sc_hd__and2_1
Xclkbuf_5_19__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_19__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_230_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29105_ clknet_leaf_161_clk _02903_ net150 VGND VGND VPWR VPWR C_out\[77\] sky130_fd_sc_hd__dfrtp_1
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26317_ clknet_leaf_29_A_in_serial_clk _00125_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_14331_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\] VGND VGND
+ VPWR VPWR _11516_ sky130_fd_sc_hd__nand2_1
XFILLER_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23529_ _10150_ _10151_ VGND VGND VPWR VPWR _10152_ sky130_fd_sc_hd__nand2_1
XFILLER_180_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27297_ clknet_leaf_293_clk _01095_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_29036_ clknet_leaf_97_clk _02834_ net153 VGND VGND VPWR VPWR C_out\[8\] sky130_fd_sc_hd__dfrtp_1
X_14262_ systolic_inst.A_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[4\]
+ systolic_inst.B_outs\[15\]\[3\] VGND VGND VPWR VPWR _11449_ sky130_fd_sc_hd__a22oi_1
X_17050_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[11\]\[12\]
+ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_169_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26248_ clknet_leaf_11_A_in_serial_clk _00056_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16001_ _12992_ _12998_ VGND VGND VPWR VPWR _13000_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13213_ deser_A.word_buffer\[51\] deser_A.serial_word\[51\] net128 VGND VGND VPWR
+ VPWR _00061_ sky130_fd_sc_hd__mux2_1
XFILLER_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14193_ _11380_ _11381_ VGND VGND VPWR VPWR _11382_ sky130_fd_sc_hd__or2_1
X_26179_ _11247_ _11248_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__nor2_1
XFILLER_139_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13144_ _11288_ _11290_ _11296_ systolic_inst.ce_local VGND VGND VPWR VPWR _11297_
+ sky130_fd_sc_hd__o31ai_2
XFILLER_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_B_in_serial_clk clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_25_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_140_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17952_ net107 _05143_ _05144_ _05145_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__o31ai_1
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_221_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_221_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16903_ _04128_ _04187_ _04185_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__a21oi_1
XFILLER_215_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Left_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17883_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[5\] _05077_
+ _05078_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__a22o_1
XFILLER_211_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19622_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.B_outs\[1\]\[2\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__mux2_1
XFILLER_113_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16834_ _04094_ _04151_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_109_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19553_ _06579_ _06580_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__nor2_1
XFILLER_150_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16765_ _04084_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__or2_1
X_13977_ deser_B.shift_reg\[11\] deser_B.shift_reg\[12\] net125 VGND VGND VPWR VPWR
+ _00803_ sky130_fd_sc_hd__mux2_1
XFILLER_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18504_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[4\] _05633_ _05634_
+ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__nand4_2
XFILLER_206_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15716_ _12739_ _12744_ _12768_ VGND VGND VPWR VPWR _12769_ sky130_fd_sc_hd__or3_1
XFILLER_111_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19484_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[7\]\[12\]
+ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16696_ _03966_ _03993_ _03992_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__a21oi_1
XFILLER_146_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18435_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.A_outs\[8\]\[1\] systolic_inst.B_outs\[8\]\[2\]
+ systolic_inst.B_outs\[8\]\[3\] VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__and4_1
XFILLER_221_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15647_ _12646_ _12664_ _12663_ VGND VGND VPWR VPWR _12702_ sky130_fd_sc_hd__o21a_1
XFILLER_59_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18366_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[26\]
+ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_140_Left_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15578_ _12634_ _12633_ VGND VGND VPWR VPWR _12635_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_25_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17317_ _04573_ _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__or2_1
X_14529_ net118 _11705_ _11706_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__a21oi_1
X_18297_ _05466_ _05465_ systolic_inst.acc_wires\[9\]\[15\] net107 VGND VGND VPWR
+ VPWR _01377_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_228_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_228_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17248_ _04506_ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_228_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17179_ systolic_inst.A_outs\[10\]\[1\] systolic_inst.A_outs\[9\]\[1\] net120 VGND
+ VGND VPWR VPWR _01267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20190_ systolic_inst.acc_wires\[6\]\[24\] systolic_inst.acc_wires\[6\]\[25\] systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__o21a_1
XFILLER_116_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22900_ _09541_ _09543_ _09579_ VGND VGND VPWR VPWR _09580_ sky130_fd_sc_hd__a21o_1
X_23880_ _10467_ VGND VGND VPWR VPWR _10468_ sky130_fd_sc_hd__inv_2
X_22831_ _09451_ _09486_ _09485_ VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__a21oi_1
XFILLER_77_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25550_ systolic_inst.acc_wires\[0\]\[26\] C_out\[26\] net53 VGND VGND VPWR VPWR
+ _02852_ sky130_fd_sc_hd__mux2_1
X_22762_ _09444_ _09445_ VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__nand2_1
XFILLER_77_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24501_ C_out\[77\] net100 net80 ser_C.shift_reg\[77\] _10720_ VGND VGND VPWR VPWR
+ _02327_ sky130_fd_sc_hd__a221o_1
X_21713_ systolic_inst.A_outs\[3\]\[6\] _08519_ _08518_ VGND VGND VPWR VPWR _08520_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25481_ _00008_ _11216_ systolic_inst.cycle_cnt\[16\] VGND VGND VPWR VPWR _11218_
+ sky130_fd_sc_hd__or3b_1
XFILLER_213_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ net122 _09380_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__nand2_1
XFILLER_201_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27220_ clknet_leaf_291_clk _01018_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_24432_ net114 ser_C.shift_reg\[44\] VGND VGND VPWR VPWR _10686_ sky130_fd_sc_hd__and2_1
X_21644_ systolic_inst.A_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[5\] VGND VGND VPWR
+ VPWR _08453_ sky130_fd_sc_hd__nand2_1
XFILLER_240_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24363_ C_out\[8\] net104 _10643_ ser_C.shift_reg\[8\] _10651_ VGND VGND VPWR VPWR
+ _02258_ sky130_fd_sc_hd__a221o_1
XFILLER_177_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27151_ clknet_leaf_251_clk _00949_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_40 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ systolic_inst.A_outs\[3\]\[1\] systolic_inst.B_outs\[3\]\[5\] systolic_inst.B_outs\[3\]\[6\]
+ systolic_inst.A_outs\[3\]\[0\] VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__a22oi_1
XFILLER_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23314_ net121 _09941_ _09942_ _09943_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_151_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26102_ deser_B.serial_word\[57\] deser_B.shift_reg\[57\] net56 VGND VGND VPWR VPWR
+ _03404_ sky130_fd_sc_hd__mux2_1
XFILLER_20_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20526_ _07422_ _07427_ _07458_ net109 VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_151_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27082_ clknet_leaf_29_B_in_serial_clk _00880_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_24294_ _10620_ systolic_inst.A_shift\[11\]\[2\] net71 VGND VGND VPWR VPWR _02220_
+ sky130_fd_sc_hd__mux2_1
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23245_ _09883_ _09885_ _09891_ VGND VGND VPWR VPWR _09892_ sky130_fd_sc_hd__a21o_1
XFILLER_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26033_ systolic_inst.acc_wires\[15\]\[29\] ser_C.parallel_data\[509\] net38 VGND
+ VGND VPWR VPWR _03335_ sky130_fd_sc_hd__mux2_1
XFILLER_101_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20457_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[9\] _07392_ net120
+ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__mux2_1
XFILLER_106_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23176_ _09817_ _09824_ _09830_ _09823_ VGND VGND VPWR VPWR _09833_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_164_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20388_ _07324_ _07321_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__and2b_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22127_ _08872_ _08875_ VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27984_ clknet_leaf_151_clk _01782_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_160_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22058_ _08825_ _08827_ _08830_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__and3_1
X_26935_ clknet_leaf_21_A_in_serial_clk _00733_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13900_ deser_A.serial_word\[61\] deser_A.shift_reg\[61\] _00002_ VGND VGND VPWR
+ VPWR _00726_ sky130_fd_sc_hd__mux2_1
X_21009_ _07873_ _07881_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__xnor2_1
X_29654_ clknet_leaf_6_B_in_serial_clk _03449_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_26866_ clknet_leaf_94_clk net84 net151 VGND VGND VPWR VPWR B_in_valid sky130_fd_sc_hd__dfrtp_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14880_ systolic_inst.A_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[4\]
+ systolic_inst.B_outs\[14\]\[3\] VGND VGND VPWR VPWR _12003_ sky130_fd_sc_hd__a22oi_1
XFILLER_75_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28605_ clknet_leaf_135_clk _02403_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[153\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13831_ deser_B.bit_idx\[3\] _11323_ _11325_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25817_ systolic_inst.acc_wires\[9\]\[5\] C_out\[293\] net14 VGND VGND VPWR VPWR
+ _03119_ sky130_fd_sc_hd__mux2_1
X_29585_ clknet_leaf_19_B_in_serial_clk _03380_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26797_ clknet_leaf_86_clk _00599_ net153 VGND VGND VPWR VPWR B_in\[69\] sky130_fd_sc_hd__dfrtp_1
Xmax_cap20 net21 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_6
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap31 net32 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_6
Xmax_cap42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_3_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28536_ clknet_leaf_160_clk _02334_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[84\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap53 net54 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_8
X_16550_ _03898_ _03899_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13762_ B_in\[69\] deser_B.word_buffer\[69\] net87 VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25748_ systolic_inst.acc_wires\[7\]\[0\] C_out\[224\] net42 VGND VGND VPWR VPWR
+ _03050_ sky130_fd_sc_hd__mux2_1
Xmax_cap64 net66 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_12
XFILLER_44_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap75 net76 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_16
XFILLER_43_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap86 net88 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_8
X_15501_ _12523_ _12559_ VGND VGND VPWR VPWR _12560_ sky130_fd_sc_hd__or2_1
XFILLER_188_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap97 net100 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_12
XFILLER_56_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28467_ clknet_leaf_100_clk _02265_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16481_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[16\]
+ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13693_ B_in\[0\] deser_B.word_buffer\[0\] net85 VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__mux2_1
X_25679_ systolic_inst.acc_wires\[4\]\[27\] C_out\[155\] net30 VGND VGND VPWR VPWR
+ _02981_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18220_ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__inv_2
X_27418_ clknet_leaf_215_clk _01216_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_15432_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[3\] _12489_ _12490_
+ VGND VGND VPWR VPWR _12493_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_117_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28398_ clknet_leaf_33_clk _02196_ VGND VGND VPWR VPWR systolic_inst.A_shift\[16\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18151_ _05337_ _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__nor2_1
XFILLER_200_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27349_ clknet_leaf_233_clk _01147_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_14_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15363_ systolic_inst.A_outs\[13\]\[7\] systolic_inst.A_outs\[12\]\[7\] net115 VGND
+ VGND VPWR VPWR _01081_ sky130_fd_sc_hd__mux2_1
XFILLER_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17102_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[20\]
+ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__nand2_1
XFILLER_200_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ _11482_ _11499_ VGND VGND VPWR VPWR _11500_ sky130_fd_sc_hd__nor2_1
X_18082_ _05262_ _05270_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__xnor2_1
X_15294_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[22\]
+ VGND VGND VPWR VPWR _12386_ sky130_fd_sc_hd__nand2_1
XFILLER_102_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29019_ clknet_leaf_93_clk _02817_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17033_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[11\]\[10\]
+ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__or2_1
X_14245_ _11401_ _11432_ VGND VGND VPWR VPWR _11433_ sky130_fd_sc_hd__xor2_1
XFILLER_109_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_223_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_223_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14176_ systolic_inst.A_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[3\]
+ systolic_inst.B_outs\[15\]\[4\] VGND VGND VPWR VPWR _11366_ sky130_fd_sc_hd__nand4_1
XFILLER_139_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13127_ _11281_ VGND VGND VPWR VPWR _11282_ sky130_fd_sc_hd__inv_2
X_18984_ _06076_ _06077_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17935_ _05094_ _05128_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17866_ systolic_inst.A_outs\[9\]\[2\] systolic_inst.B_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\]
+ systolic_inst.A_outs\[9\]\[1\] VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__a22o_1
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19605_ _06628_ _06631_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__nand2_1
XFILLER_66_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16817_ systolic_inst.A_outs\[11\]\[3\] systolic_inst.A_outs\[11\]\[4\] systolic_inst.B_outs\[11\]\[6\]
+ systolic_inst.B_outs\[11\]\[7\] VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__and4b_1
XFILLER_96_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17797_ systolic_inst.B_outs\[8\]\[4\] systolic_inst.B_outs\[4\]\[4\] net121 VGND
+ VGND VPWR VPWR _01342_ sky130_fd_sc_hd__mux2_1
XFILLER_226_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_217_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19536_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[20\]
+ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_217_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16748_ systolic_inst.A_outs\[11\]\[1\] _11262_ systolic_inst.B_outs\[11\]\[6\] systolic_inst.A_outs\[11\]\[2\]
+ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19467_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[7\]\[10\]
+ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16679_ _03999_ _04001_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__nor2_1
X_18418_ systolic_inst.B_outs\[7\]\[7\] systolic_inst.B_outs\[3\]\[7\] net119 VGND
+ VGND VPWR VPWR _01409_ sky130_fd_sc_hd__mux2_1
XFILLER_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19398_ _06454_ _06455_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18349_ _05503_ _05507_ _05510_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__nand3_1
XFILLER_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21360_ _08195_ _08200_ _08208_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__a21o_1
XFILLER_120_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20311_ _07207_ _07225_ _07224_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__a21bo_1
XFILLER_200_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21291_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[4\]\[6\]
+ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__nand2_1
X_23030_ _09672_ _09675_ _09705_ VGND VGND VPWR VPWR _09706_ sky130_fd_sc_hd__o21a_1
X_20242_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[1\]
+ systolic_inst.B_outs\[5\]\[0\] VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__a22o_1
XFILLER_200_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20173_ _07098_ _07099_ _07121_ _07141_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__a211o_1
XFILLER_143_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24981_ C_out\[317\] net97 net80 ser_C.shift_reg\[317\] _10960_ VGND VGND VPWR VPWR
+ _02567_ sky130_fd_sc_hd__a221o_1
XFILLER_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26720_ clknet_leaf_31_B_in_serial_clk _00523_ net134 VGND VGND VPWR VPWR deser_B.word_buffer\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23932_ systolic_inst.A_shift\[3\]\[4\] net71 _11333_ A_in\[28\] VGND VGND VPWR VPWR
+ _01982_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_198_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26651_ clknet_leaf_25_B_in_serial_clk _00454_ net137 VGND VGND VPWR VPWR deser_B.word_buffer\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23863_ systolic_inst.acc_wires\[0\]\[24\] systolic_inst.acc_wires\[0\]\[25\] systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _10454_ sky130_fd_sc_hd__o21a_1
XFILLER_44_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25602_ systolic_inst.acc_wires\[2\]\[14\] C_out\[78\] net51 VGND VGND VPWR VPWR
+ _02904_ sky130_fd_sc_hd__mux2_1
XFILLER_211_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22814_ _09494_ _09495_ VGND VGND VPWR VPWR _09496_ sky130_fd_sc_hd__and2_1
X_29370_ clknet_leaf_232_clk _03168_ net147 VGND VGND VPWR VPWR C_out\[342\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26582_ clknet_leaf_28_A_in_serial_clk _00385_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23794_ _10394_ _10395_ _10388_ _10393_ VGND VGND VPWR VPWR _10396_ sky130_fd_sc_hd__o211ai_1
XFILLER_198_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28321_ clknet_leaf_0_clk _02119_ VGND VGND VPWR VPWR systolic_inst.A_shift\[28\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25533_ systolic_inst.acc_wires\[0\]\[9\] C_out\[9\] net33 VGND VGND VPWR VPWR _02835_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_1115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_236_Left_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22745_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[5\] VGND VGND VPWR
+ VPWR _09429_ sky130_fd_sc_hd__nand2_1
XFILLER_198_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28252_ clknet_leaf_78_clk _02050_ VGND VGND VPWR VPWR systolic_inst.B_shift\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25464_ systolic_inst.cycle_cnt\[11\] systolic_inst.cycle_cnt\[10\] _11199_ _11202_
+ VGND VGND VPWR VPWR _11206_ sky130_fd_sc_hd__and4_1
X_22676_ systolic_inst.A_outs\[1\]\[3\] systolic_inst.A_outs\[0\]\[3\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27203_ clknet_leaf_259_clk _01001_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_24415_ C_out\[34\] _11302_ net81 ser_C.shift_reg\[34\] _10677_ VGND VGND VPWR VPWR
+ _02284_ sky130_fd_sc_hd__a221o_1
X_21627_ _08397_ _08400_ _08436_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__o21ai_1
XFILLER_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28183_ clknet_leaf_65_clk _01981_ VGND VGND VPWR VPWR systolic_inst.A_shift\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25395_ systolic_inst.A_shift\[3\]\[5\] A_in\[21\] net59 VGND VGND VPWR VPWR _11167_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27134_ clknet_leaf_85_clk _00932_ VGND VGND VPWR VPWR systolic_inst.B_shift\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24346_ net10 net7 VGND VGND VPWR VPWR _10643_ sky130_fd_sc_hd__nor2_8
XFILLER_205_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21558_ _08339_ _08342_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__nor2_1
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20509_ _07440_ _07441_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__xnor2_1
X_27065_ clknet_leaf_8_B_in_serial_clk _00863_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_24277_ systolic_inst.B_shift\[27\]\[2\] B_in\[90\] net59 VGND VGND VPWR VPWR _10612_
+ sky130_fd_sc_hd__mux2_1
X_21489_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[1\]
+ systolic_inst.A_outs\[3\]\[2\] VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__and4_1
X_14030_ deser_B.shift_reg\[64\] deser_B.shift_reg\[65\] net126 VGND VGND VPWR VPWR
+ _00856_ sky130_fd_sc_hd__mux2_1
X_23228_ _09833_ _09834_ _09856_ _09876_ VGND VGND VPWR VPWR _09877_ sky130_fd_sc_hd__a211o_1
X_26016_ systolic_inst.acc_wires\[15\]\[12\] ser_C.parallel_data\[492\] net37 VGND
+ VGND VPWR VPWR _03318_ sky130_fd_sc_hd__mux2_1
XFILLER_181_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23159_ _11713_ _09818_ VGND VGND VPWR VPWR _09819_ sky130_fd_sc_hd__nor2_1
XFILLER_136_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27967_ clknet_leaf_165_clk _01765_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_15981_ systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[1\] VGND VGND
+ VPWR VPWR _12981_ sky130_fd_sc_hd__nand2_1
XFILLER_67_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17720_ _04938_ _04944_ _04945_ net60 VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__a31o_1
XFILLER_76_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14932_ _12035_ _12052_ VGND VGND VPWR VPWR _12054_ sky130_fd_sc_hd__xor2_1
XFILLER_94_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26918_ clknet_leaf_4_A_in_serial_clk _00716_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27898_ clknet_leaf_45_clk _01696_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29637_ clknet_leaf_28_B_in_serial_clk _03432_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _04888_ _04887_ systolic_inst.acc_wires\[10\]\[11\] net105 VGND VGND VPWR
+ VPWR _01309_ sky130_fd_sc_hd__a2bb2o_1
X_26849_ clknet_leaf_66_clk _00651_ net134 VGND VGND VPWR VPWR B_in\[121\] sky130_fd_sc_hd__dfrtp_1
X_14863_ _11985_ _11986_ _11959_ VGND VGND VPWR VPWR _11987_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_67_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16602_ _03921_ _03927_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__xnor2_1
X_13814_ B_in\[121\] deser_B.word_buffer\[121\] net89 VGND VGND VPWR VPWR _00651_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29568_ clknet_leaf_17_B_in_serial_clk _03363_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_17582_ _04829_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__inv_2
X_14794_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[3\]
+ systolic_inst.A_outs\[14\]\[4\] VGND VGND VPWR VPWR _11920_ sky130_fd_sc_hd__and4_1
XFILLER_1_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19321_ _06349_ _06351_ _06350_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__o21ba_1
XFILLER_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28519_ clknet_leaf_155_clk _02317_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_16533_ _03884_ _03885_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13745_ B_in\[52\] deser_B.word_buffer\[52\] net85 VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__mux2_1
X_29499_ clknet_leaf_268_clk _03297_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[471\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19252_ systolic_inst.A_outs\[7\]\[4\] systolic_inst.B_outs\[7\]\[6\] _11261_ systolic_inst.A_outs\[7\]\[3\]
+ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_143_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16464_ _03820_ _03822_ _03826_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__nand3_1
XFILLER_32_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13676_ deser_B.word_buffer\[112\] deser_B.serial_word\[112\] net123 VGND VGND VPWR
+ VPWR _00513_ sky130_fd_sc_hd__mux2_1
XFILLER_188_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18203_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[9\]\[2\]
+ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__or2_1
XFILLER_223_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15415_ _12455_ _12458_ _12475_ _12476_ VGND VGND VPWR VPWR _12477_ sky130_fd_sc_hd__a211o_1
X_19183_ systolic_inst.A_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[5\] VGND VGND VPWR
+ VPWR _06248_ sky130_fd_sc_hd__nand2_1
XFILLER_19_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16395_ net67 _03765_ _03767_ systolic_inst.acc_wires\[12\]\[4\] net108 VGND VGND
+ VPWR VPWR _01174_ sky130_fd_sc_hd__a32o_1
XFILLER_185_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18134_ _05320_ _05321_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__and2_1
X_15346_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[30\]
+ VGND VGND VPWR VPWR _12430_ sky130_fd_sc_hd__nand2_1
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18065_ net116 _05254_ _05255_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__a21oi_1
X_15277_ _12370_ _12371_ VGND VGND VPWR VPWR _12372_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17016_ _04315_ _04316_ _04314_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__a21bo_1
XFILLER_176_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14228_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[6\] VGND VGND
+ VPWR VPWR _11416_ sky130_fd_sc_hd__nand2_1
XFILLER_119_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_242_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ systolic_inst.A_outs\[15\]\[0\] systolic_inst.B_outs\[15\]\[3\] systolic_inst.A_outs\[15\]\[3\]
+ systolic_inst.B_outs\[15\]\[0\] VGND VGND VPWR VPWR _11350_ sky130_fd_sc_hd__a22oi_1
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_242_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _06062_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__or2_1
XFILLER_85_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17918_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[6\]
+ systolic_inst.A_outs\[9\]\[7\] VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__nand4_1
X_18898_ _06002_ _06004_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__nand2_1
XFILLER_26_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17849_ _05021_ _05024_ _05043_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__nand3_1
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20860_ systolic_inst.B_outs\[4\]\[3\] _07729_ VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__nand2_1
XFILLER_214_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19519_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[17\]
+ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__xor2_2
X_20791_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[26\]
+ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22530_ _09253_ _09255_ _09257_ systolic_inst.acc_wires\[2\]\[9\] net109 VGND VGND
+ VPWR VPWR _01819_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_18_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22461_ _08984_ _09122_ _09192_ _09190_ VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__a31oi_1
XFILLER_210_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_951 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24200_ systolic_inst.B_shift\[22\]\[7\] net71 _11333_ B_in\[119\] VGND VGND VPWR
+ VPWR _02161_ sky130_fd_sc_hd__a22o_1
X_21412_ _08245_ _08249_ _08252_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__a21o_1
XFILLER_148_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25180_ net111 ser_C.shift_reg\[418\] VGND VGND VPWR VPWR _11060_ sky130_fd_sc_hd__and2_1
X_22392_ _09097_ _09099_ _09098_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__o21ba_1
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24131_ systolic_inst.A_shift\[30\]\[5\] A_in\[117\] net59 VGND VGND VPWR VPWR _10567_
+ sky130_fd_sc_hd__mux2_1
X_21343_ _08182_ _08185_ _08189_ _08193_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__a211o_1
XFILLER_194_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_208_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24062_ _10548_ systolic_inst.B_shift\[15\]\[2\] net70 VGND VGND VPWR VPWR _02060_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21274_ _08135_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__inv_2
XFILLER_116_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23013_ _09660_ _09688_ VGND VGND VPWR VPWR _09689_ sky130_fd_sc_hd__nand2b_1
XFILLER_116_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20225_ systolic_inst.A_outs\[5\]\[2\] systolic_inst.A_outs\[4\]\[2\] net116 VGND
+ VGND VPWR VPWR _01588_ sky130_fd_sc_hd__mux2_1
X_28870_ clknet_leaf_300_clk _02668_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[418\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_146_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27821_ clknet_leaf_307_clk _01619_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_104_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20156_ _07119_ _07125_ _07126_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_142_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27752_ clknet_leaf_208_clk _01550_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20087_ _07061_ _07063_ _07059_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__a21bo_1
X_24964_ net111 ser_C.shift_reg\[310\] VGND VGND VPWR VPWR _10952_ sky130_fd_sc_hd__and2_1
XFILLER_131_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26703_ clknet_leaf_7_B_in_serial_clk _00506_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_23915_ _10490_ systolic_inst.B_shift\[18\]\[1\] _11332_ VGND VGND VPWR VPWR _01971_
+ sky130_fd_sc_hd__mux2_1
X_27683_ clknet_leaf_197_clk _01481_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_217_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24895_ C_out\[274\] net101 net73 ser_C.shift_reg\[274\] _10917_ VGND VGND VPWR VPWR
+ _02524_ sky130_fd_sc_hd__a221o_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29422_ clknet_leaf_340_clk _03220_ net131 VGND VGND VPWR VPWR C_out\[394\] sky130_fd_sc_hd__dfrtp_1
XFILLER_217_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26634_ clknet_leaf_12_B_in_serial_clk _00437_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_23846_ _10419_ _10425_ _10430_ _10436_ VGND VGND VPWR VPWR _10439_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_101_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29353_ clknet_leaf_228_clk _03151_ net140 VGND VGND VPWR VPWR C_out\[325\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26565_ clknet_leaf_25_A_in_serial_clk _00368_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_23777_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[0\]\[13\]
+ VGND VGND VPWR VPWR _10381_ sky130_fd_sc_hd__xor2_1
XFILLER_26_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20989_ _07809_ _07821_ _07820_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__o21a_1
XFILLER_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28304_ clknet_leaf_67_clk _02102_ VGND VGND VPWR VPWR systolic_inst.B_shift\[27\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25516_ systolic_inst.cycle_cnt\[29\] _11279_ _11237_ VGND VGND VPWR VPWR _11240_
+ sky130_fd_sc_hd__a21oi_1
X_13530_ deser_A.shift_reg\[94\] deser_A.shift_reg\[95\] net129 VGND VGND VPWR VPWR
+ _00367_ sky130_fd_sc_hd__mux2_1
XFILLER_242_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22728_ _09411_ _09412_ _09393_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__o21ai_1
X_29284_ clknet_leaf_325_clk _03082_ net136 VGND VGND VPWR VPWR C_out\[256\] sky130_fd_sc_hd__dfrtp_1
X_26496_ clknet_leaf_7_A_in_serial_clk _00299_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28235_ clknet_leaf_130_clk _02033_ VGND VGND VPWR VPWR systolic_inst.B_shift\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25447_ systolic_inst.cycle_cnt\[5\] systolic_inst.cycle_cnt\[4\] _11190_ VGND VGND
+ VPWR VPWR _11195_ sky130_fd_sc_hd__and3_1
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13461_ deser_A.shift_reg\[25\] deser_A.shift_reg\[26\] deser_A.receiving VGND VGND
+ VPWR VPWR _00298_ sky130_fd_sc_hd__mux2_1
XFILLER_13_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22659_ _09364_ _09366_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15200_ _12304_ _12305_ VGND VGND VPWR VPWR _12306_ sky130_fd_sc_hd__nor2_1
X_28166_ clknet_leaf_95_clk _01964_ VGND VGND VPWR VPWR systolic_inst.B_shift\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16180_ _03560_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25378_ _11158_ systolic_inst.B_shift\[14\]\[4\] net71 VGND VGND VPWR VPWR _02766_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13392_ A_in\[101\] deser_A.word_buffer\[101\] _00003_ VGND VGND VPWR VPWR _00240_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27117_ clknet_leaf_32_B_in_serial_clk _00915_ net134 VGND VGND VPWR VPWR deser_B.shift_reg\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15131_ _12175_ _12223_ _12222_ VGND VGND VPWR VPWR _12247_ sky130_fd_sc_hd__o21ba_1
X_24329_ systolic_inst.A_shift\[10\]\[4\] A_in\[36\] net59 VGND VGND VPWR VPWR _10638_
+ sky130_fd_sc_hd__mux2_1
X_28097_ clknet_leaf_109_clk _01895_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_182_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27048_ clknet_leaf_24_B_in_serial_clk _00846_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15062_ _12178_ _12179_ VGND VGND VPWR VPWR _12180_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14013_ deser_B.shift_reg\[47\] deser_B.shift_reg\[48\] net125 VGND VGND VPWR VPWR
+ _00839_ sky130_fd_sc_hd__mux2_1
XFILLER_49_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19870_ _06860_ _06868_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__nand2_1
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18821_ _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__inv_2
X_28999_ clknet_leaf_92_clk _02797_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18752_ _05806_ _05843_ _05842_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__a21bo_1
XFILLER_216_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15964_ systolic_inst.A_outs\[12\]\[5\] systolic_inst.A_shift\[24\]\[5\] net115 VGND
+ VGND VPWR VPWR _01143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17703_ net106 systolic_inst.acc_wires\[10\]\[18\] net68 _04933_ VGND VGND VPWR VPWR
+ _01316_ sky130_fd_sc_hd__a22o_1
XFILLER_188_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14915_ systolic_inst.B_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[5\]
+ systolic_inst.B_outs\[14\]\[3\] VGND VGND VPWR VPWR _12037_ sky130_fd_sc_hd__a22oi_1
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18683_ systolic_inst.A_outs\[8\]\[5\] systolic_inst.B_outs\[8\]\[6\] _11259_ systolic_inst.A_outs\[8\]\[4\]
+ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__o2bb2a_1
X_15895_ _12923_ _12922_ systolic_inst.acc_wires\[13\]\[21\] net108 VGND VGND VPWR
+ VPWR _01127_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[10\]\[8\]
+ _04871_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__and3_1
XFILLER_1_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14846_ systolic_inst.A_outs\[14\]\[2\] systolic_inst.B_outs\[14\]\[3\] systolic_inst.A_outs\[14\]\[3\]
+ systolic_inst.B_outs\[14\]\[4\] VGND VGND VPWR VPWR _11970_ sky130_fd_sc_hd__and4_1
XFILLER_236_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17565_ _04813_ _04815_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__nand2_1
XFILLER_205_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14777_ systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[3\]
+ systolic_inst.B_outs\[14\]\[0\] VGND VGND VPWR VPWR _11904_ sky130_fd_sc_hd__a22o_1
XFILLER_44_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19304_ _06306_ _06365_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16516_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[22\]
+ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__nand2_1
XFILLER_220_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13728_ B_in\[35\] deser_B.word_buffer\[35\] net86 VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__mux2_1
XFILLER_32_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17496_ _04715_ _04717_ _04716_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__o21ba_1
XFILLER_108_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19235_ _06263_ _06265_ _06298_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__a21o_1
X_16447_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[12\]\[12\]
+ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__nor2_1
X_13659_ deser_B.word_buffer\[95\] deser_B.serial_word\[95\] net123 VGND VGND VPWR
+ VPWR _00496_ sky130_fd_sc_hd__mux2_1
XFILLER_34_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19166_ _06164_ _06165_ _06196_ _06194_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__a31o_1
X_16378_ _03750_ _03752_ _03745_ _03747_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_41_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18117_ _05259_ _05275_ _05273_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__o21a_1
X_15329_ _12414_ _12415_ VGND VGND VPWR VPWR _12416_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_10_A_in_serial_clk clknet_2_2__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_10_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_144_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19097_ _06123_ _06140_ _06139_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__a21bo_1
XFILLER_195_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18048_ _05237_ _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__nand2b_1
XFILLER_172_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20010_ _07000_ _07003_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_203_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19999_ _06993_ _06992_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__nand2b_1
XFILLER_150_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21961_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[3\]\[14\]
+ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__nand2_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23700_ net63 _10314_ _10315_ systolic_inst.acc_wires\[0\]\[1\] _11258_ VGND VGND
+ VPWR VPWR _01931_ sky130_fd_sc_hd__a32o_1
XFILLER_27_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20912_ _07779_ _07786_ _07787_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__nand3_1
XFILLER_242_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21892_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[3\]\[4\]
+ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__nand2_1
X_24680_ net111 ser_C.shift_reg\[168\] VGND VGND VPWR VPWR _10810_ sky130_fd_sc_hd__and2_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23631_ _10178_ _10182_ _10215_ _10217_ VGND VGND VPWR VPWR _10252_ sky130_fd_sc_hd__o31a_1
XFILLER_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20843_ net117 systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[0\] VGND
+ VGND VPWR VPWR _07724_ sky130_fd_sc_hd__and3_1
XFILLER_42_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26350_ clknet_leaf_65_clk _00157_ net135 VGND VGND VPWR VPWR A_in\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20774_ _07672_ _07676_ _07679_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__nand3_1
X_23562_ _10178_ _10182_ VGND VGND VPWR VPWR _10184_ sky130_fd_sc_hd__nor2_1
XFILLER_35_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25301_ ser_C.parallel_data\[477\] net102 net74 ser_C.shift_reg\[477\] _11120_ VGND
+ VGND VPWR VPWR _02727_ sky130_fd_sc_hd__a221o_1
XFILLER_35_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22513_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[2\]\[7\]
+ VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__nand2_1
XFILLER_126_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23493_ _10115_ _10116_ VGND VGND VPWR VPWR _10117_ sky130_fd_sc_hd__or2_1
X_26281_ clknet_leaf_19_A_in_serial_clk _00089_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_196_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_170_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_170_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_167_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28020_ clknet_leaf_154_clk _01818_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22444_ _09096_ _09181_ VGND VGND VPWR VPWR _09183_ sky130_fd_sc_hd__nand2_1
X_25232_ net111 ser_C.shift_reg\[444\] VGND VGND VPWR VPWR _11086_ sky130_fd_sc_hd__and2_1
XFILLER_136_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22375_ _09116_ VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__inv_2
XFILLER_164_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25163_ C_out\[408\] net101 net73 ser_C.shift_reg\[408\] _11051_ VGND VGND VPWR VPWR
+ _02658_ sky130_fd_sc_hd__a221o_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24114_ systolic_inst.B_shift\[27\]\[1\] net72 _11333_ B_in\[121\] VGND VGND VPWR
+ VPWR _02099_ sky130_fd_sc_hd__a22o_1
X_21326_ net63 _08178_ _08179_ systolic_inst.acc_wires\[4\]\[11\] _11258_ VGND VGND
+ VPWR VPWR _01693_ sky130_fd_sc_hd__a32o_1
XFILLER_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25094_ net113 ser_C.shift_reg\[375\] VGND VGND VPWR VPWR _11017_ sky130_fd_sc_hd__and2_1
XFILLER_159_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28922_ clknet_leaf_268_clk _02720_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[470\]
+ sky130_fd_sc_hd__dfrtp_1
X_24045_ systolic_inst.B_shift\[4\]\[2\] B_in\[2\] _00008_ VGND VGND VPWR VPWR _10540_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21257_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[4\]\[1\]
+ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__or2_1
XFILLER_151_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20208_ _07165_ _07168_ _07167_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__o21a_1
XFILLER_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28853_ clknet_leaf_345_clk _02651_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[401\]
+ sky130_fd_sc_hd__dfrtp_1
X_21188_ _07982_ _07986_ _08022_ _08055_ _08020_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__o311a_1
XFILLER_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27804_ clknet_leaf_41_clk _01602_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_20139_ _07111_ _07113_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__xor2_1
X_28784_ clknet_leaf_231_clk _02582_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[332\]
+ sky130_fd_sc_hd__dfrtp_1
X_25996_ systolic_inst.acc_wires\[14\]\[24\] ser_C.parallel_data\[472\] net25 VGND
+ VGND VPWR VPWR _03298_ sky130_fd_sc_hd__mux2_1
XFILLER_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27735_ clknet_leaf_132_clk _01533_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_20_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24947_ C_out\[300\] net103 net76 ser_C.shift_reg\[300\] _10943_ VGND VGND VPWR VPWR
+ _02550_ sky130_fd_sc_hd__a221o_1
XFILLER_46_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14700_ _11847_ _11850_ _11852_ VGND VGND VPWR VPWR _11853_ sky130_fd_sc_hd__or3_1
XFILLER_234_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_242_Right_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27666_ clknet_leaf_203_clk _01464_ net147 VGND VGND VPWR VPWR systolic_inst.A_outs\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_15680_ _12732_ _12733_ VGND VGND VPWR VPWR _12734_ sky130_fd_sc_hd__nor2_1
XFILLER_218_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24878_ net110 ser_C.shift_reg\[267\] VGND VGND VPWR VPWR _10909_ sky130_fd_sc_hd__and2_1
X_29405_ clknet_leaf_194_clk _03203_ net146 VGND VGND VPWR VPWR C_out\[377\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26617_ clknet_leaf_21_B_in_serial_clk _00420_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14631_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[15\]
+ VGND VGND VPWR VPWR _11794_ sky130_fd_sc_hd__nor2_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23829_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[21\]
+ VGND VGND VPWR VPWR _10425_ sky130_fd_sc_hd__xor2_1
XFILLER_2_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27597_ clknet_leaf_33_clk _01395_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_120_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29336_ clknet_leaf_216_clk _03134_ net140 VGND VGND VPWR VPWR C_out\[308\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ systolic_inst.B_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[4\]
+ systolic_inst.A_outs\[10\]\[5\] VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__and4_1
XFILLER_144_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14562_ _11728_ _11729_ _11727_ VGND VGND VPWR VPWR _11735_ sky130_fd_sc_hd__a21bo_1
X_26548_ clknet_leaf_26_A_in_serial_clk _00351_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _03679_ _03680_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_81_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13513_ deser_A.shift_reg\[77\] deser_A.shift_reg\[78\] net129 VGND VGND VPWR VPWR
+ _00350_ sky130_fd_sc_hd__mux2_1
XFILLER_92_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29267_ clknet_leaf_190_clk _03065_ net146 VGND VGND VPWR VPWR C_out\[239\] sky130_fd_sc_hd__dfrtp_1
X_17281_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[4\] _04538_ _04539_
+ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__nand4_2
Xclkbuf_leaf_161_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_161_clk
+ sky130_fd_sc_hd__clkbuf_8
X_26479_ clknet_leaf_13_A_in_serial_clk _00282_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14493_ _11643_ _11647_ VGND VGND VPWR VPWR _11674_ sky130_fd_sc_hd__nor2_1
XFILLER_158_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19020_ systolic_inst.B_outs\[6\]\[1\] systolic_inst.B_outs\[2\]\[1\] net119 VGND
+ VGND VPWR VPWR _01467_ sky130_fd_sc_hd__mux2_1
X_28218_ clknet_leaf_80_clk _02016_ VGND VGND VPWR VPWR systolic_inst.B_shift\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16232_ _03557_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_133_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13444_ deser_A.shift_reg\[8\] deser_A.shift_reg\[9\] deser_A.receiving VGND VGND
+ VPWR VPWR _00281_ sky130_fd_sc_hd__mux2_1
XFILLER_186_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29198_ clknet_leaf_141_clk _02996_ net149 VGND VGND VPWR VPWR C_out\[170\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload308 clknet_leaf_118_clk VGND VGND VPWR VPWR clkload308/Y sky130_fd_sc_hd__bufinv_16
XFILLER_139_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28149_ clknet_leaf_108_clk _01947_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload319 clknet_leaf_114_clk VGND VGND VPWR VPWR clkload319/Y sky130_fd_sc_hd__inv_8
Xclkload16 clknet_5_18__leaf_clk VGND VGND VPWR VPWR clkload16/X sky130_fd_sc_hd__clkbuf_8
X_16163_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__inv_2
Xclkload27 clknet_leaf_328_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__clkinvlp_4
X_13375_ A_in\[84\] deser_A.word_buffer\[84\] net94 VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload38 clknet_leaf_322_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__inv_8
XFILLER_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload49 clknet_leaf_331_clk VGND VGND VPWR VPWR clkload49/X sky130_fd_sc_hd__clkbuf_8
XFILLER_177_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15114_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[13\] _12230_ net118
+ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16094_ _13087_ _13088_ VGND VGND VPWR VPWR _13089_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_90_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19922_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[11\] _06919_ net119
+ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__mux2_1
XFILLER_138_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15045_ _12162_ _12163_ VGND VGND VPWR VPWR _12164_ sky130_fd_sc_hd__nor2_1
XFILLER_218_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19853_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[10\] VGND
+ VGND VPWR VPWR _06852_ sky130_fd_sc_hd__and2_1
XFILLER_116_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18804_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[8\]\[1\]
+ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__or2_1
X_19784_ _06784_ _06781_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__and2b_1
X_16996_ _04302_ _04303_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__a21o_1
XFILLER_7_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15947_ systolic_inst.acc_wires\[13\]\[28\] systolic_inst.acc_wires\[13\]\[29\] systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12967_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18735_ _05792_ _05797_ _05827_ _05825_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_88_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_237_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18666_ _05790_ _05791_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_237_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[19\]
+ VGND VGND VPWR VPWR _12909_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1058 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14829_ _11925_ _11952_ VGND VGND VPWR VPWR _11954_ sky130_fd_sc_hd__or2_1
XFILLER_75_1410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17617_ _04856_ _04857_ _04858_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__and3_1
XFILLER_24_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18597_ _05688_ _05689_ _05687_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__a21o_1
XFILLER_240_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17548_ _04714_ _04798_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__or2_1
XFILLER_162_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_152_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_152_clk
+ sky130_fd_sc_hd__clkbuf_8
X_17479_ _04695_ _04697_ _04732_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_17_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19218_ systolic_inst.A_outs\[7\]\[4\] systolic_inst.B_outs\[7\]\[5\] VGND VGND VPWR
+ VPWR _06282_ sky130_fd_sc_hd__nand2_1
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20490_ _07388_ _07389_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__nand2_1
XFILLER_118_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19149_ systolic_inst.A_outs\[7\]\[1\] systolic_inst.B_outs\[7\]\[6\] _06214_ VGND
+ VGND VPWR VPWR _06215_ sky130_fd_sc_hd__and3_1
XFILLER_121_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_184_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22160_ _08884_ _08907_ VGND VGND VPWR VPWR _08908_ sky130_fd_sc_hd__nand2_1
XFILLER_195_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21111_ _07980_ _07981_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__nor2_1
X_22091_ systolic_inst.B_outs\[1\]\[5\] systolic_inst.B_shift\[1\]\[5\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__mux2_1
XFILLER_161_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21042_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[6\] _07885_ _07884_
+ systolic_inst.A_outs\[4\]\[3\] VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__a32o_1
XFILLER_232_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25850_ systolic_inst.acc_wires\[10\]\[6\] C_out\[326\] net12 VGND VGND VPWR VPWR
+ _03152_ sky130_fd_sc_hd__mux2_1
XFILLER_41_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24801_ C_out\[227\] net99 net79 ser_C.shift_reg\[227\] _10870_ VGND VGND VPWR VPWR
+ _02477_ sky130_fd_sc_hd__a221o_1
XFILLER_68_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25781_ systolic_inst.acc_wires\[8\]\[1\] C_out\[257\] net21 VGND VGND VPWR VPWR
+ _03083_ sky130_fd_sc_hd__mux2_1
XFILLER_80_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22993_ _09656_ _09669_ VGND VGND VPWR VPWR _09670_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27520_ clknet_leaf_232_clk _01318_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24732_ net112 ser_C.shift_reg\[194\] VGND VGND VPWR VPWR _10836_ sky130_fd_sc_hd__and2_1
XFILLER_41_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21944_ _08721_ _08732_ VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__and2_1
XFILLER_83_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27451_ clknet_leaf_236_clk _01249_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_215_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24663_ C_out\[158\] net104 net76 ser_C.shift_reg\[158\] _10801_ VGND VGND VPWR VPWR
+ _02408_ sky130_fd_sc_hd__a221o_1
X_21875_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[3\]\[0\]
+ _08671_ _08672_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26402_ clknet_leaf_32_clk _00209_ net133 VGND VGND VPWR VPWR A_in\[70\] sky130_fd_sc_hd__dfrtp_1
X_23614_ systolic_inst.B_outs\[0\]\[6\] systolic_inst.A_outs\[0\]\[6\] _10193_ VGND
+ VGND VPWR VPWR _10235_ sky130_fd_sc_hd__a21oi_1
X_20826_ _07723_ _07722_ systolic_inst.acc_wires\[5\]\[31\] net106 VGND VGND VPWR
+ VPWR _01649_ sky130_fd_sc_hd__a2bb2o_1
X_27382_ clknet_leaf_339_clk _01180_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_5_A_in_serial_clk clknet_2_2__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_5_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_24594_ net113 ser_C.shift_reg\[125\] VGND VGND VPWR VPWR _10767_ sky130_fd_sc_hd__and2_1
XFILLER_168_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29121_ clknet_leaf_163_clk _02919_ net150 VGND VGND VPWR VPWR C_out\[93\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26333_ clknet_leaf_59_clk _00140_ net143 VGND VGND VPWR VPWR A_in\[1\] sky130_fd_sc_hd__dfrtp_1
X_23545_ _10125_ _10128_ _10166_ VGND VGND VPWR VPWR _10168_ sky130_fd_sc_hd__and3_1
X_20757_ _07663_ _07664_ _07661_ VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_143_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29052_ clknet_leaf_106_clk _02850_ net151 VGND VGND VPWR VPWR C_out\[24\] sky130_fd_sc_hd__dfrtp_1
X_26264_ clknet_leaf_4_A_in_serial_clk _00072_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23476_ _10097_ _10098_ _10054_ _10056_ VGND VGND VPWR VPWR _10101_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_33_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_33_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_20688_ net109 systolic_inst.acc_wires\[5\]\[10\] net64 _07606_ VGND VGND VPWR VPWR
+ _01628_ sky130_fd_sc_hd__a22o_1
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28003_ clknet_leaf_153_clk _01801_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25215_ C_out\[434\] net101 net73 ser_C.shift_reg\[434\] _11077_ VGND VGND VPWR VPWR
+ _02684_ sky130_fd_sc_hd__a221o_1
X_22427_ _09164_ _09165_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__xor2_1
XFILLER_137_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26195_ systolic_inst.A_shift\[30\]\[1\] net71 _11333_ A_in\[121\] VGND VGND VPWR
+ VPWR _03485_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_186_Left_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13160_ _11306_ VGND VGND VPWR VPWR _11307_ sky130_fd_sc_hd__inv_2
X_25146_ net110 ser_C.shift_reg\[401\] VGND VGND VPWR VPWR _11043_ sky130_fd_sc_hd__and2_1
XFILLER_200_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22358_ _09098_ _09099_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__or2_1
XFILLER_139_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21309_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[4\]\[9\]
+ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__nand2_1
X_22289_ _09031_ _09032_ VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_167_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25077_ C_out\[365\] net97 net77 ser_C.shift_reg\[365\] _11008_ VGND VGND VPWR VPWR
+ _02615_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_167_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24028_ _10531_ systolic_inst.B_shift\[4\]\[1\] net72 VGND VGND VPWR VPWR _02043_
+ sky130_fd_sc_hd__mux2_1
X_28905_ clknet_leaf_271_clk _02703_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16850_ _04132_ _04167_ systolic_inst.A_outs\[11\]\[7\] VGND VGND VPWR VPWR _04168_
+ sky130_fd_sc_hd__and3b_1
XFILLER_215_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28836_ clknet_leaf_327_clk _02634_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[384\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15801_ _12839_ _12840_ _12838_ VGND VGND VPWR VPWR _12843_ sky130_fd_sc_hd__a21bo_1
XFILLER_63_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28767_ clknet_leaf_224_clk _02565_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[315\]
+ sky130_fd_sc_hd__dfrtp_1
X_16781_ _04097_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__xnor2_1
X_13993_ deser_B.shift_reg\[27\] deser_B.shift_reg\[28\] net125 VGND VGND VPWR VPWR
+ _00819_ sky130_fd_sc_hd__mux2_1
X_25979_ systolic_inst.acc_wires\[14\]\[7\] ser_C.parallel_data\[455\] net25 VGND
+ VGND VPWR VPWR _03281_ sky130_fd_sc_hd__mux2_1
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_195_Left_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18520_ _05617_ _05619_ _05649_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__a211oi_1
X_27718_ clknet_leaf_188_clk _01516_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _12781_ _12782_ VGND VGND VPWR VPWR _12784_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_122_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28698_ clknet_leaf_189_clk _02496_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[246\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18451_ _05582_ _05583_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ systolic_inst.B_outs\[13\]\[6\] systolic_inst.A_outs\[13\]\[6\] _11272_ systolic_inst.A_outs\[13\]\[5\]
+ VGND VGND VPWR VPWR _12717_ sky130_fd_sc_hd__o2bb2a_1
X_27649_ clknet_leaf_325_clk _01447_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_73_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17402_ _04618_ _04620_ _04656_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__nand3_1
XFILLER_226_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14614_ net105 systolic_inst.acc_wires\[15\]\[12\] net69 _11779_ VGND VGND VPWR VPWR
+ _00990_ sky130_fd_sc_hd__a22o_1
X_18382_ _05537_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__nand2_1
XFILLER_215_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15594_ _12616_ _12649_ VGND VGND VPWR VPWR _12650_ sky130_fd_sc_hd__xor2_1
XFILLER_187_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29319_ clknet_leaf_297_clk _03117_ net138 VGND VGND VPWR VPWR C_out\[291\] sky130_fd_sc_hd__dfrtp_1
X_17333_ _04588_ _04589_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__xnor2_1
X_14545_ net69 _11718_ _11720_ systolic_inst.acc_wires\[15\]\[2\] net107 VGND VGND
+ VPWR VPWR _00980_ sky130_fd_sc_hd__a32o_1
XFILLER_230_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_134_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_230_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17264_ _04496_ _04522_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__xor2_1
XFILLER_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14476_ _11656_ _11655_ VGND VGND VPWR VPWR _11657_ sky130_fd_sc_hd__nand2b_1
XFILLER_186_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19003_ _06092_ _06093_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__nand2_1
X_16215_ systolic_inst.A_outs\[12\]\[3\] systolic_inst.A_outs\[12\]\[4\] systolic_inst.B_outs\[12\]\[6\]
+ systolic_inst.B_outs\[12\]\[7\] VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__and4b_1
XFILLER_70_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload105 clknet_leaf_279_clk VGND VGND VPWR VPWR clkload105/Y sky130_fd_sc_hd__clkinvlp_4
X_13427_ _11312_ _11313_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__nor2_1
Xclkload116 clknet_leaf_276_clk VGND VGND VPWR VPWR clkload116/Y sky130_fd_sc_hd__inv_6
X_17195_ net107 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[0\] _04459_
+ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__a21o_1
XFILLER_127_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload127 clknet_leaf_261_clk VGND VGND VPWR VPWR clkload127/Y sky130_fd_sc_hd__bufinv_16
Xclkload138 clknet_leaf_252_clk VGND VGND VPWR VPWR clkload138/Y sky130_fd_sc_hd__inv_8
X_16146_ _03527_ _03530_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__xnor2_1
Xclkload149 clknet_leaf_297_clk VGND VGND VPWR VPWR clkload149/X sky130_fd_sc_hd__clkbuf_4
X_13358_ A_in\[67\] deser_A.word_buffer\[67\] net96 VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__mux2_1
XFILLER_114_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16077_ _13067_ _13071_ VGND VGND VPWR VPWR _13073_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_226_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13289_ deser_A.word_buffer\[127\] deser_A.serial_word\[127\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19905_ _06900_ _06901_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_36_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15028_ systolic_inst.B_outs\[14\]\[5\] systolic_inst.A_outs\[14\]\[6\] VGND VGND
+ VPWR VPWR _12147_ sky130_fd_sc_hd__nand2_1
XFILLER_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19836_ _06835_ _06834_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__nand2b_1
XFILLER_9_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_239_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19767_ _06717_ _06718_ _06731_ _06730_ _06699_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__o32a_1
XFILLER_209_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 B_in_frame_sync VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
X_16979_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[11\]\[2\]
+ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__nand2_1
XFILLER_77_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18718_ _05840_ _05841_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__xnor2_1
X_19698_ _06701_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__inv_2
XFILLER_224_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18649_ _05740_ _05742_ _05741_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__o21ba_1
XFILLER_224_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21660_ _08466_ _08467_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__xor2_1
XFILLER_80_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20611_ net109 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] VGND
+ VGND VPWR VPWR _07541_ sky130_fd_sc_hd__and2_1
X_21591_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[6\] _08399_
+ _08401_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_125_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_162_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23330_ _09937_ _09957_ _09958_ VGND VGND VPWR VPWR _09959_ sky130_fd_sc_hd__and3_1
XFILLER_162_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20542_ _07435_ _07474_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_1279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23261_ _09904_ VGND VGND VPWR VPWR _09905_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_211_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20473_ _07405_ _07406_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25000_ net111 ser_C.shift_reg\[328\] VGND VGND VPWR VPWR _10970_ sky130_fd_sc_hd__and2_1
X_22212_ _08956_ _08957_ VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__or2_1
X_23192_ systolic_inst.acc_wires\[1\]\[16\] systolic_inst.acc_wires\[1\]\[17\] systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09847_ sky130_fd_sc_hd__o21a_1
X_22143_ _08880_ _08883_ VGND VGND VPWR VPWR _08891_ sky130_fd_sc_hd__and2b_1
XFILLER_195_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22074_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[31\]
+ VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__xnor2_1
X_26951_ clknet_leaf_26_A_in_serial_clk _00749_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_160_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25902_ systolic_inst.acc_wires\[11\]\[26\] C_out\[378\] net41 VGND VGND VPWR VPWR
+ _03204_ sky130_fd_sc_hd__mux2_1
X_21025_ _07896_ _07897_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_162_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29670_ clknet_leaf_29_B_in_serial_clk _03465_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_162_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26882_ clknet_leaf_9_A_in_serial_clk _00680_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28621_ clknet_leaf_141_clk _02419_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[169\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_12_B_in_serial_clk clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_12_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_25833_ systolic_inst.acc_wires\[9\]\[21\] C_out\[309\] net13 VGND VGND VPWR VPWR
+ _03135_ sky130_fd_sc_hd__mux2_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28552_ clknet_leaf_172_clk _02350_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_25764_ systolic_inst.acc_wires\[7\]\[16\] C_out\[240\] net42 VGND VGND VPWR VPWR
+ _03066_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22976_ _09516_ _09652_ VGND VGND VPWR VPWR _09653_ sky130_fd_sc_hd__or2_1
XFILLER_216_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27503_ clknet_leaf_228_clk _01301_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_24715_ C_out\[184\] net99 net79 ser_C.shift_reg\[184\] _10827_ VGND VGND VPWR VPWR
+ _02434_ sky130_fd_sc_hd__a221o_1
XFILLER_76_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28483_ clknet_leaf_108_clk _02281_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_21927_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[3\]\[10\]
+ VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__nand2_1
X_25695_ systolic_inst.acc_wires\[5\]\[11\] C_out\[171\] net31 VGND VGND VPWR VPWR
+ _02997_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27434_ clknet_leaf_235_clk _01232_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24646_ net7 ser_C.shift_reg\[151\] VGND VGND VPWR VPWR _10793_ sky130_fd_sc_hd__and2_1
X_21858_ _08657_ _08659_ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__xor2_1
XFILLER_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20809_ net106 systolic_inst.acc_wires\[5\]\[28\] net68 _07709_ VGND VGND VPWR VPWR
+ _01646_ sky130_fd_sc_hd__a22o_1
X_27365_ clknet_leaf_340_clk _01163_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24577_ C_out\[115\] net100 net80 ser_C.shift_reg\[115\] _10758_ VGND VGND VPWR VPWR
+ _02365_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_116_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_156_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21789_ _08593_ _08592_ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__nand2b_1
X_29104_ clknet_leaf_166_clk _02902_ net152 VGND VGND VPWR VPWR C_out\[76\] sky130_fd_sc_hd__dfrtp_1
XFILLER_211_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26316_ clknet_leaf_29_A_in_serial_clk _00124_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_14330_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[7\] _11485_ _11483_
+ VGND VGND VPWR VPWR _11515_ sky130_fd_sc_hd__a31o_1
XFILLER_184_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23528_ _10106_ _10149_ VGND VGND VPWR VPWR _10151_ sky130_fd_sc_hd__nand2_1
XFILLER_54_1379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27296_ clknet_leaf_292_clk _01094_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29035_ clknet_leaf_124_clk _02833_ net144 VGND VGND VPWR VPWR C_out\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14261_ systolic_inst.B_outs\[15\]\[3\] systolic_inst.A_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\]
+ systolic_inst.A_outs\[15\]\[4\] VGND VGND VPWR VPWR _11448_ sky130_fd_sc_hd__and4_1
X_26247_ clknet_leaf_18_A_in_serial_clk _00055_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_23459_ _10083_ _10082_ VGND VGND VPWR VPWR _10084_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_115_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16000_ _12992_ _12998_ VGND VGND VPWR VPWR _12999_ sky130_fd_sc_hd__or2_1
XFILLER_137_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13212_ deser_A.word_buffer\[50\] deser_A.serial_word\[50\] net128 VGND VGND VPWR
+ VPWR _00060_ sky130_fd_sc_hd__mux2_1
X_26178_ ser_C.bit_idx\[2\] _11245_ _11303_ VGND VGND VPWR VPWR _11248_ sky130_fd_sc_hd__o21ai_1
X_14192_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[3\]
+ systolic_inst.A_outs\[15\]\[4\] VGND VGND VPWR VPWR _11381_ sky130_fd_sc_hd__and4_1
XFILLER_100_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13143_ _11294_ _11295_ VGND VGND VPWR VPWR _11296_ sky130_fd_sc_hd__or2_1
X_25129_ C_out\[391\] net101 net73 ser_C.shift_reg\[391\] _11034_ VGND VGND VPWR VPWR
+ _02641_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_111_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17951_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[7\] VGND
+ VGND VPWR VPWR _05145_ sky130_fd_sc_hd__nand2_1
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_221_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_221_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16902_ _04164_ _04217_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__xor2_1
X_17882_ _05045_ _05048_ _05075_ net116 VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__o31a_1
XFILLER_215_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19621_ systolic_inst.B_outs\[5\]\[1\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__mux2_1
XFILLER_120_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16833_ _04094_ _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__nand2_1
X_28819_ clknet_leaf_237_clk _02617_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19552_ systolic_inst.acc_wires\[7\]\[20\] systolic_inst.acc_wires\[7\]\[21\] systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__o21a_1
X_16764_ _04045_ _04047_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_234_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13976_ deser_B.shift_reg\[10\] deser_B.shift_reg\[11\] net125 VGND VGND VPWR VPWR
+ _00802_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15715_ _12766_ _12767_ VGND VGND VPWR VPWR _12768_ sky130_fd_sc_hd__and2b_1
X_18503_ systolic_inst.B_outs\[8\]\[3\] systolic_inst.A_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\]
+ systolic_inst.A_outs\[8\]\[2\] VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__a22o_1
XFILLER_98_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19483_ _06516_ _06525_ _06526_ _06527_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__o211a_1
XFILLER_34_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16695_ _03987_ _04010_ _04009_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__a21boi_1
XFILLER_146_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15646_ _12684_ _12700_ VGND VGND VPWR VPWR _12701_ sky130_fd_sc_hd__xor2_1
X_18434_ systolic_inst.A_outs\[8\]\[1\] systolic_inst.B_outs\[8\]\[2\] systolic_inst.B_outs\[8\]\[3\]
+ systolic_inst.A_outs\[8\]\[0\] VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__a22oi_1
XFILLER_62_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18365_ net66 _05523_ _05524_ systolic_inst.acc_wires\[9\]\[25\] net105 VGND VGND
+ VPWR VPWR _01387_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_107_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15577_ _12581_ _12598_ _12597_ VGND VGND VPWR VPWR _12634_ sky130_fd_sc_hd__o21ba_1
XFILLER_61_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17316_ systolic_inst.A_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[4\]
+ systolic_inst.B_outs\[10\]\[3\] VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__a22oi_1
XFILLER_202_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14528_ net118 systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[15\]\[0\]
+ VGND VGND VPWR VPWR _11706_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_25_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18296_ _05457_ _05460_ _05464_ _11713_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_25_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17247_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[4\]
+ systolic_inst.A_outs\[10\]\[5\] VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_228_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14459_ _11639_ _11640_ VGND VGND VPWR VPWR _11641_ sky130_fd_sc_hd__nand2_1
XFILLER_179_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17178_ systolic_inst.A_outs\[10\]\[0\] systolic_inst.A_outs\[9\]\[0\] net120 VGND
+ VGND VPWR VPWR _01266_ sky130_fd_sc_hd__mux2_1
XFILLER_190_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16129_ systolic_inst.B_outs\[12\]\[7\] _13087_ _13088_ VGND VGND VPWR VPWR _03514_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_157_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19819_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[8\] _06817_
+ _06819_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__a22o_1
XFILLER_9_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_25__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_25__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22830_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[7\] _09511_ net122
+ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__mux2_1
XFILLER_65_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22761_ _09401_ _09419_ _09418_ VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__a21bo_1
XFILLER_198_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_346_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_346_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24500_ net113 ser_C.shift_reg\[78\] VGND VGND VPWR VPWR _10720_ sky130_fd_sc_hd__and2_1
XFILLER_225_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21712_ systolic_inst.B_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[7\]
+ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__and3_1
X_25480_ _11279_ _11214_ _11217_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__and3_1
XFILLER_240_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22692_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[1\]
+ systolic_inst.B_outs\[1\]\[0\] VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__a22o_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24431_ C_out\[42\] _11302_ net81 ser_C.shift_reg\[42\] _10685_ VGND VGND VPWR VPWR
+ _02292_ sky130_fd_sc_hd__a221o_1
XFILLER_205_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21643_ _08450_ _08451_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_213_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27150_ clknet_leaf_251_clk _00948_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_205_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24362_ net7 ser_C.shift_reg\[9\] VGND VGND VPWR VPWR _10651_ sky130_fd_sc_hd__and2_1
XANTENNA_30 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21574_ _08381_ _08384_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_41 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26101_ deser_B.serial_word\[56\] deser_B.shift_reg\[56\] net56 VGND VGND VPWR VPWR
+ _03403_ sky130_fd_sc_hd__mux2_1
XFILLER_21_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23313_ _11258_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[3\] VGND
+ VGND VPWR VPWR _09943_ sky130_fd_sc_hd__and2_1
X_20525_ _07422_ _07427_ _07458_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_151_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27081_ clknet_leaf_28_B_in_serial_clk _00879_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24293_ systolic_inst.A_shift\[12\]\[2\] A_in\[50\] net59 VGND VGND VPWR VPWR _10620_
+ sky130_fd_sc_hd__mux2_1
XFILLER_181_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26032_ systolic_inst.acc_wires\[15\]\[28\] ser_C.parallel_data\[508\] net38 VGND
+ VGND VPWR VPWR _03334_ sky130_fd_sc_hd__mux2_1
X_23244_ systolic_inst.acc_wires\[1\]\[24\] systolic_inst.acc_wires\[1\]\[25\] systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09891_ sky130_fd_sc_hd__o21a_1
XFILLER_181_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20456_ _07390_ _07391_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__nor2_1
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23175_ _09832_ _09831_ systolic_inst.acc_wires\[1\]\[15\] net109 VGND VGND VPWR
+ VPWR _01889_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_164_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20387_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] _07322_ VGND
+ VGND VPWR VPWR _07324_ sky130_fd_sc_hd__a21o_1
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22126_ _08873_ _08874_ VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__nand2_1
XFILLER_136_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27983_ clknet_leaf_151_clk _01781_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26934_ clknet_leaf_21_A_in_serial_clk _00732_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_22057_ _08828_ _08829_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__or2_1
XFILLER_212_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21008_ _07879_ _07880_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__and2_1
X_26865_ clknet_leaf_89_clk deser_B.serial_toggle net5 VGND VGND VPWR VPWR deser_B.serial_toggle_sync1
+ sky130_fd_sc_hd__dfrtp_2
X_29653_ clknet_leaf_6_B_in_serial_clk _03448_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13830_ deser_B.bit_idx\[3\] _11323_ _11321_ VGND VGND VPWR VPWR _11325_ sky130_fd_sc_hd__o21ai_1
X_28604_ clknet_leaf_135_clk _02402_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[152\]
+ sky130_fd_sc_hd__dfrtp_1
X_25816_ systolic_inst.acc_wires\[9\]\[4\] C_out\[292\] net14 VGND VGND VPWR VPWR
+ _03118_ sky130_fd_sc_hd__mux2_1
X_29584_ clknet_leaf_19_B_in_serial_clk _03379_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_26796_ clknet_leaf_85_clk _00598_ net153 VGND VGND VPWR VPWR B_in\[68\] sky130_fd_sc_hd__dfrtp_1
XFILLER_235_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap21 net22 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_8
Xmax_cap32 net33 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_8
XFILLER_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28535_ clknet_leaf_160_clk _02333_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13761_ B_in\[68\] deser_B.word_buffer\[68\] net87 VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__mux2_1
Xmax_cap43 net45 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_8
X_25747_ systolic_inst.acc_wires\[6\]\[31\] C_out\[223\] net43 VGND VGND VPWR VPWR
+ _03049_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap54 _11297_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_8
XFILLER_216_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22959_ _09627_ _09635_ VGND VGND VPWR VPWR _09637_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_337_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_337_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_56_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap65 net68 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_12
XFILLER_189_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap76 _10643_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_12
XFILLER_44_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15500_ _12551_ _12557_ VGND VGND VPWR VPWR _12559_ sky130_fd_sc_hd__xnor2_1
Xmax_cap87 net88 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_8
XFILLER_231_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28466_ clknet_leaf_99_clk _02264_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_16480_ _03837_ _03840_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13692_ deser_B.serial_toggle net123 VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__xor2_1
XFILLER_189_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap98 net99 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_12
XFILLER_182_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25678_ systolic_inst.acc_wires\[4\]\[26\] C_out\[154\] net30 VGND VGND VPWR VPWR
+ _02980_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15431_ _12489_ _12491_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[3\]
+ VGND VGND VPWR VPWR _12492_ sky130_fd_sc_hd__and4b_1
X_27417_ clknet_leaf_223_clk _01215_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_203_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24629_ C_out\[141\] net104 _10643_ ser_C.shift_reg\[141\] _10784_ VGND VGND VPWR
+ VPWR _02391_ sky130_fd_sc_hd__a221o_1
XFILLER_231_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28397_ clknet_leaf_33_clk _02195_ VGND VGND VPWR VPWR systolic_inst.A_shift\[16\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ _05335_ _05336_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__and2b_1
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27348_ clknet_leaf_233_clk _01146_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_14_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15362_ systolic_inst.A_outs\[13\]\[6\] systolic_inst.A_outs\[12\]\[6\] net115 VGND
+ VGND VPWR VPWR _01080_ sky130_fd_sc_hd__mux2_1
XFILLER_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17101_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[20\]
+ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__or2_1
XFILLER_200_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14313_ _11496_ _11497_ VGND VGND VPWR VPWR _11499_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_78_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18081_ _05262_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__nand2_1
X_15293_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[22\]
+ VGND VGND VPWR VPWR _12385_ sky130_fd_sc_hd__or2_1
X_27279_ clknet_leaf_323_clk _01077_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29018_ clknet_leaf_94_clk _02816_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17032_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[11\]\[10\]
+ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14244_ _11430_ _11431_ VGND VGND VPWR VPWR _11432_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_74_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_223_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_223_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_7_B_in_serial_clk clknet_2_2__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_7_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_14175_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[4\] VGND VGND
+ VPWR VPWR _11365_ sky130_fd_sc_hd__and2_1
XFILLER_178_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13126_ deser_A.bit_idx\[3\] deser_A.bit_idx\[5\] deser_A.bit_idx\[4\] _11280_ VGND
+ VGND VPWR VPWR _11281_ sky130_fd_sc_hd__and4_1
XFILLER_152_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18983_ _06070_ _06074_ _06071_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a21bo_1
XFILLER_26_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17934_ _05124_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17865_ systolic_inst.A_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[2\] systolic_inst.B_outs\[9\]\[3\]
+ systolic_inst.B_outs\[9\]\[4\] VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__and4_1
XFILLER_93_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19604_ _06629_ _06630_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__nand2_1
X_16816_ systolic_inst.B_outs\[11\]\[5\] systolic_inst.A_outs\[11\]\[5\] VGND VGND
+ VPWR VPWR _04135_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17796_ systolic_inst.B_outs\[8\]\[3\] systolic_inst.B_outs\[4\]\[3\] net121 VGND
+ VGND VPWR VPWR _01341_ sky130_fd_sc_hd__mux2_1
XFILLER_242_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_217_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19535_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[20\]
+ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_187_Right_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_328_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_328_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13959_ deser_A.serial_word\[120\] deser_A.shift_reg\[120\] _00002_ VGND VGND VPWR
+ VPWR _00785_ sky130_fd_sc_hd__mux2_1
X_16747_ systolic_inst.A_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[2\] systolic_inst.B_outs\[11\]\[6\]
+ systolic_inst.B_outs\[11\]\[7\] VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__and4b_1
XFILLER_59_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19466_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[7\]\[10\]
+ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16678_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.A_outs\[11\]\[1\] systolic_inst.B_outs\[11\]\[5\]
+ systolic_inst.B_outs\[11\]\[6\] VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__and4_1
XFILLER_222_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18417_ systolic_inst.B_outs\[7\]\[6\] systolic_inst.B_outs\[3\]\[6\] net119 VGND
+ VGND VPWR VPWR _01408_ sky130_fd_sc_hd__mux2_1
X_15629_ _12682_ _12683_ VGND VGND VPWR VPWR _12684_ sky130_fd_sc_hd__nand2_1
XFILLER_107_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19397_ _06373_ _06434_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18348_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__inv_2
XFILLER_72_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18279_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[9\]\[13\]
+ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__nand2_1
XFILLER_174_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20310_ _07248_ _07249_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__nor2_1
XFILLER_194_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21290_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[4\]\[6\]
+ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__and2_1
XFILLER_238_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20241_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.A_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\]
+ systolic_inst.A_outs\[5\]\[1\] VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__and4_1
XFILLER_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20172_ _07120_ _07127_ _07132_ _07137_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__nand4_1
XFILLER_153_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_206_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24980_ net111 ser_C.shift_reg\[318\] VGND VGND VPWR VPWR _10960_ sky130_fd_sc_hd__and2_1
XFILLER_233_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23931_ systolic_inst.A_shift\[3\]\[3\] net72 _11333_ A_in\[27\] VGND VGND VPWR VPWR
+ _01981_ sky130_fd_sc_hd__a22o_1
XFILLER_44_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_198_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26650_ clknet_leaf_25_B_in_serial_clk _00453_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23862_ _10451_ _10452_ VGND VGND VPWR VPWR _10453_ sky130_fd_sc_hd__nand2_1
XFILLER_45_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25601_ systolic_inst.acc_wires\[2\]\[13\] C_out\[77\] net51 VGND VGND VPWR VPWR
+ _02903_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22813_ systolic_inst.B_outs\[1\]\[5\] _11277_ _09461_ systolic_inst.A_outs\[1\]\[0\]
+ VGND VGND VPWR VPWR _09495_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_140_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26581_ clknet_leaf_28_A_in_serial_clk _00384_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23793_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[15\]
+ VGND VGND VPWR VPWR _10395_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_319_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_319_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_955 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28320_ clknet_leaf_0_clk _02118_ VGND VGND VPWR VPWR systolic_inst.A_shift\[28\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25532_ systolic_inst.acc_wires\[0\]\[8\] C_out\[8\] net33 VGND VGND VPWR VPWR _02834_
+ sky130_fd_sc_hd__mux2_1
X_22744_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[5\] VGND VGND VPWR
+ VPWR _09428_ sky130_fd_sc_hd__and2_1
XFILLER_129_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28251_ clknet_leaf_95_clk _02049_ VGND VGND VPWR VPWR systolic_inst.B_shift\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25463_ _11203_ _11204_ systolic_inst.cycle_cnt\[10\] VGND VGND VPWR VPWR _02804_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22675_ systolic_inst.A_outs\[1\]\[2\] systolic_inst.A_outs\[0\]\[2\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__mux2_1
XFILLER_241_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27202_ clknet_leaf_262_clk _01000_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_1343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24414_ net114 ser_C.shift_reg\[35\] VGND VGND VPWR VPWR _10677_ sky130_fd_sc_hd__and2_1
XFILLER_197_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21626_ _08402_ _08434_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__xnor2_1
X_28182_ clknet_leaf_66_clk _01980_ VGND VGND VPWR VPWR systolic_inst.A_shift\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25394_ _11166_ systolic_inst.A_shift\[2\]\[4\] net71 VGND VGND VPWR VPWR _02774_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27133_ clknet_leaf_71_clk _00931_ VGND VGND VPWR VPWR systolic_inst.B_shift\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24345_ net7 ser_C.shift_reg\[1\] VGND VGND VPWR VPWR _10642_ sky130_fd_sc_hd__and2_1
X_21557_ _08345_ _08367_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27064_ clknet_leaf_8_B_in_serial_clk _00862_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_20508_ _07441_ _07440_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__nand2b_1
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24276_ _10611_ systolic_inst.B_shift\[23\]\[1\] net71 VGND VGND VPWR VPWR _02211_
+ sky130_fd_sc_hd__mux2_1
X_21488_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.A_outs\[3\]\[2\] VGND VGND VPWR
+ VPWR _08303_ sky130_fd_sc_hd__nand2_1
XFILLER_181_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26015_ systolic_inst.acc_wires\[15\]\[11\] ser_C.parallel_data\[491\] net37 VGND
+ VGND VPWR VPWR _03317_ sky130_fd_sc_hd__mux2_1
XFILLER_88_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23227_ _09855_ _09862_ _09867_ _09872_ VGND VGND VPWR VPWR _09876_ sky130_fd_sc_hd__nand4_1
X_20439_ _07374_ _07373_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__nand2b_1
XFILLER_101_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23158_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[1\]\[12\]
+ _09814_ VGND VGND VPWR VPWR _09818_ sky130_fd_sc_hd__and3_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22109_ systolic_inst.A_outs\[2\]\[1\] systolic_inst.B_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[3\]
+ systolic_inst.A_outs\[2\]\[0\] VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__a22oi_1
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15980_ _12980_ _12978_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[1\]
+ net108 VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_216_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27966_ clknet_leaf_166_clk _01764_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_23089_ _09755_ _09756_ _09757_ VGND VGND VPWR VPWR _09759_ sky130_fd_sc_hd__and3_1
XFILLER_212_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14931_ _12035_ _12052_ VGND VGND VPWR VPWR _12053_ sky130_fd_sc_hd__or2_1
XFILLER_103_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26917_ clknet_leaf_10_A_in_serial_clk _00715_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27897_ clknet_leaf_46_clk _01695_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29636_ clknet_leaf_27_B_in_serial_clk _03431_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_14862_ _11983_ _11984_ _11953_ _11956_ VGND VGND VPWR VPWR _11986_ sky130_fd_sc_hd__o211a_1
X_17650_ _04876_ _04881_ _04886_ net60 VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__a31o_1
X_26848_ clknet_leaf_63_clk _00650_ net135 VGND VGND VPWR VPWR B_in\[120\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13813_ B_in\[120\] deser_B.word_buffer\[120\] net89 VGND VGND VPWR VPWR _00650_
+ sky130_fd_sc_hd__mux2_1
X_16601_ _03925_ _03926_ _03921_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__or3b_1
XFILLER_91_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17581_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[10\]\[0\]
+ _04827_ _04828_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__and4_1
XFILLER_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29567_ clknet_leaf_17_B_in_serial_clk _03362_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_26779_ clknet_leaf_54_clk _00581_ net143 VGND VGND VPWR VPWR B_in\[51\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14793_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.A_outs\[14\]\[4\] VGND VGND
+ VPWR VPWR _11919_ sky130_fd_sc_hd__nand2_1
XFILLER_63_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19320_ _06379_ _06380_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__xnor2_1
X_16532_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[24\]
+ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_63_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28518_ clknet_leaf_155_clk _02316_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_13744_ B_in\[51\] deser_B.word_buffer\[51\] net85 VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__mux2_1
XFILLER_17_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29498_ clknet_leaf_268_clk _03296_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[470\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19251_ systolic_inst.A_outs\[7\]\[3\] systolic_inst.A_outs\[7\]\[4\] systolic_inst.B_outs\[7\]\[6\]
+ systolic_inst.B_outs\[7\]\[7\] VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__and4b_1
X_16463_ _03824_ _03825_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__nand2_1
X_13675_ deser_B.word_buffer\[111\] deser_B.serial_word\[111\] net123 VGND VGND VPWR
+ VPWR _00512_ sky130_fd_sc_hd__mux2_1
X_28449_ clknet_leaf_34_clk _02247_ VGND VGND VPWR VPWR systolic_inst.A_shift\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_232_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15414_ _12473_ _12474_ _12467_ VGND VGND VPWR VPWR _12476_ sky130_fd_sc_hd__a21oi_1
X_18202_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[9\]\[2\]
+ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__nand2_1
X_19182_ _06245_ _06246_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16394_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__inv_2
X_18133_ systolic_inst.A_outs\[9\]\[6\] _11263_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__or2_1
X_15345_ _12419_ _12422_ _12425_ _12428_ VGND VGND VPWR VPWR _12429_ sky130_fd_sc_hd__o31a_1
XFILLER_223_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18064_ net116 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[10\] VGND
+ VGND VPWR VPWR _05255_ sky130_fd_sc_hd__nor2_1
X_15276_ _12366_ _12368_ _12365_ VGND VGND VPWR VPWR _12371_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17015_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[11\]\[7\]
+ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__or2_1
X_14227_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[5\] systolic_inst.B_outs\[15\]\[6\]
+ systolic_inst.A_outs\[15\]\[0\] VGND VGND VPWR VPWR _11415_ sky130_fd_sc_hd__a22oi_1
XFILLER_160_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14158_ _11340_ _11348_ VGND VGND VPWR VPWR _11349_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_242_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ systolic_inst.B_outs\[2\]\[7\] VGND VGND VPWR VPWR _11265_ sky130_fd_sc_hd__inv_2
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14089_ deser_B.shift_reg\[123\] deser_B.shift_reg\[124\] net126 VGND VGND VPWR VPWR
+ _00915_ sky130_fd_sc_hd__mux2_1
X_18966_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[24\]
+ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__and2_1
XFILLER_230_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[6\] systolic_inst.A_outs\[9\]\[7\]
+ systolic_inst.B_outs\[9\]\[0\] VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__a22o_1
XFILLER_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18897_ _05997_ _06003_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__nand2_1
XFILLER_227_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_201_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_201_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17848_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__inv_2
XFILLER_242_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17779_ _04993_ _04996_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__or2_1
XFILLER_241_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_193_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19518_ net105 systolic_inst.acc_wires\[7\]\[16\] _06556_ _06558_ VGND VGND VPWR
+ VPWR _01506_ sky130_fd_sc_hd__a22o_1
XFILLER_81_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20790_ net68 _07692_ _07693_ systolic_inst.acc_wires\[5\]\[25\] net106 VGND VGND
+ VPWR VPWR _01643_ sky130_fd_sc_hd__a32o_1
XFILLER_165_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19449_ _06497_ _06498_ _06491_ _06495_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_18_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22460_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[14\] _09198_ net122
+ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__mux2_1
XFILLER_195_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21411_ _08245_ _08249_ _08252_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__nand3_1
XFILLER_31_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22391_ _09129_ _09130_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24130_ _10566_ systolic_inst.A_shift\[29\]\[4\] net71 VGND VGND VPWR VPWR _02110_
+ sky130_fd_sc_hd__mux2_1
X_21342_ _08186_ _08189_ _08193_ _08188_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__o211a_1
XFILLER_190_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_208_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3__f_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_2_3__leaf_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
X_24061_ systolic_inst.B_shift\[19\]\[2\] B_in\[26\] net59 VGND VGND VPWR VPWR _10548_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21273_ _08125_ _08129_ _08132_ _08133_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_208_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23012_ _09686_ _09687_ VGND VGND VPWR VPWR _09688_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20224_ systolic_inst.A_outs\[5\]\[1\] systolic_inst.A_outs\[4\]\[1\] net116 VGND
+ VGND VPWR VPWR _01587_ sky130_fd_sc_hd__mux2_1
XFILLER_11_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_223_Right_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20155_ _07126_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__inv_2
X_27820_ clknet_leaf_40_clk _01618_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20086_ _07066_ _07067_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__nand2_1
X_27751_ clknet_leaf_209_clk _01549_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24963_ C_out\[308\] net103 net76 ser_C.shift_reg\[308\] _10951_ VGND VGND VPWR VPWR
+ _02558_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
X_26702_ clknet_leaf_7_B_in_serial_clk _00505_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_23914_ systolic_inst.B_shift\[22\]\[1\] B_in\[81\] _00008_ VGND VGND VPWR VPWR _10490_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27682_ clknet_leaf_200_clk _01480_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24894_ net110 ser_C.shift_reg\[275\] VGND VGND VPWR VPWR _10917_ sky130_fd_sc_hd__and2_1
XFILLER_73_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26633_ clknet_leaf_11_B_in_serial_clk _00436_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_29421_ clknet_leaf_334_clk _03219_ net131 VGND VGND VPWR VPWR C_out\[393\] sky130_fd_sc_hd__dfrtp_1
X_23845_ _10438_ _10437_ systolic_inst.acc_wires\[0\]\[23\] _11258_ VGND VGND VPWR
+ VPWR _01953_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26564_ clknet_leaf_27_A_in_serial_clk _00367_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_29352_ clknet_leaf_228_clk _03150_ net138 VGND VGND VPWR VPWR C_out\[324\] sky130_fd_sc_hd__dfrtp_1
X_23776_ _11258_ systolic_inst.acc_wires\[0\]\[12\] net63 _10380_ VGND VGND VPWR VPWR
+ _01942_ sky130_fd_sc_hd__a22o_1
XFILLER_72_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20988_ _07843_ _07861_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__xor2_1
XFILLER_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25515_ systolic_inst.cycle_cnt\[29\] _11237_ VGND VGND VPWR VPWR _11239_ sky130_fd_sc_hd__and2_1
X_28303_ clknet_leaf_67_clk _02101_ VGND VGND VPWR VPWR systolic_inst.B_shift\[27\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22727_ _09408_ _09410_ _09391_ VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__a21oi_1
X_29283_ clknet_leaf_190_clk _03081_ net146 VGND VGND VPWR VPWR C_out\[255\] sky130_fd_sc_hd__dfrtp_1
XFILLER_129_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26495_ clknet_leaf_7_A_in_serial_clk _00298_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28234_ clknet_leaf_130_clk _02032_ VGND VGND VPWR VPWR systolic_inst.B_shift\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25446_ _11193_ _11194_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__and2_1
X_13460_ deser_A.shift_reg\[24\] deser_A.shift_reg\[25\] deser_A.receiving VGND VGND
+ VPWR VPWR _00297_ sky130_fd_sc_hd__mux2_1
X_22658_ _09359_ _09362_ _09361_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__o21a_1
XFILLER_230_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28165_ clknet_leaf_91_clk _01963_ VGND VGND VPWR VPWR systolic_inst.B_shift\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21609_ systolic_inst.A_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[7\] VGND VGND VPWR
+ VPWR _08419_ sky130_fd_sc_hd__and2b_1
XFILLER_220_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25377_ systolic_inst.B_shift\[18\]\[4\] B_in\[52\] net59 VGND VGND VPWR VPWR _11158_
+ sky130_fd_sc_hd__mux2_1
X_13391_ A_in\[100\] deser_A.word_buffer\[100\] _00003_ VGND VGND VPWR VPWR _00239_
+ sky130_fd_sc_hd__mux2_1
X_22589_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[18\]
+ VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__nand2_1
XFILLER_103_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
X_27116_ clknet_leaf_31_B_in_serial_clk _00914_ net134 VGND VGND VPWR VPWR deser_B.shift_reg\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_15130_ _12175_ _12245_ VGND VGND VPWR VPWR _12246_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24328_ _10637_ systolic_inst.A_shift\[9\]\[3\] net70 VGND VGND VPWR VPWR _02237_
+ sky130_fd_sc_hd__mux2_1
X_28096_ clknet_leaf_109_clk _01894_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_194_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27047_ clknet_leaf_25_B_in_serial_clk _00845_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15061_ systolic_inst.A_outs\[14\]\[5\] systolic_inst.B_outs\[14\]\[6\] systolic_inst.A_outs\[14\]\[6\]
+ systolic_inst.B_outs\[14\]\[7\] VGND VGND VPWR VPWR _12179_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_131_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24259_ systolic_inst.A_shift\[16\]\[2\] net70 net83 systolic_inst.A_shift\[17\]\[2\]
+ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__a22o_1
XFILLER_181_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14012_ deser_B.shift_reg\[46\] deser_B.shift_reg\[47\] net125 VGND VGND VPWR VPWR
+ _00838_ sky130_fd_sc_hd__mux2_1
XFILLER_153_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18820_ _05928_ _05932_ _05935_ _05936_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__o211a_1
XFILLER_7_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28998_ clknet_leaf_104_clk _02796_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_110_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18751_ _05873_ _05874_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__nand2_1
X_27949_ clknet_leaf_178_clk _01747_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15963_ systolic_inst.A_outs\[12\]\[4\] systolic_inst.A_shift\[24\]\[4\] net115 VGND
+ VGND VPWR VPWR _01142_ sky130_fd_sc_hd__mux2_1
XFILLER_209_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_87_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_191_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17702_ _04930_ _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__xor2_1
XFILLER_208_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14914_ systolic_inst.B_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[4\]
+ systolic_inst.A_outs\[14\]\[5\] VGND VGND VPWR VPWR _12036_ sky130_fd_sc_hd__and4_1
XFILLER_62_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15894_ _12913_ _12919_ _12920_ net61 VGND VGND VPWR VPWR _12923_ sky130_fd_sc_hd__a31o_1
X_18682_ systolic_inst.A_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[5\] systolic_inst.B_outs\[8\]\[6\]
+ systolic_inst.B_outs\[8\]\[7\] VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__and4b_1
XFILLER_209_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29619_ clknet_leaf_4_B_in_serial_clk _03414_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_17633_ _04869_ _04871_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__nand2_1
XFILLER_236_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14845_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[4\] VGND VGND
+ VPWR VPWR _11969_ sky130_fd_sc_hd__nand2_1
XFILLER_223_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14776_ _11892_ _11902_ VGND VGND VPWR VPWR _11903_ sky130_fd_sc_hd__or2_1
X_17564_ _04791_ _04814_ _04793_ _04768_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_223_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19303_ _06362_ _06363_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__xnor2_1
X_13727_ B_in\[34\] deser_B.word_buffer\[34\] net86 VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__mux2_1
XFILLER_147_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16515_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[22\]
+ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__or2_1
XFILLER_32_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17495_ _04745_ _04746_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19234_ _06272_ _06297_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13658_ deser_B.word_buffer\[94\] deser_B.serial_word\[94\] net123 VGND VGND VPWR
+ VPWR _00495_ sky130_fd_sc_hd__mux2_1
X_16446_ _03807_ _03809_ _03810_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_45_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19165_ _06198_ _06229_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16377_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[12\]\[2\]
+ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__or2_1
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13589_ deser_B.word_buffer\[25\] deser_B.serial_word\[25\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__mux2_1
XFILLER_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_41_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15328_ _12408_ _12412_ _12409_ VGND VGND VPWR VPWR _12415_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_41_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18116_ _05292_ _05304_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__xnor2_1
XFILLER_219_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19096_ _06144_ _06162_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15259_ _12355_ _12356_ VGND VGND VPWR VPWR _12357_ sky130_fd_sc_hd__nand2_1
X_18047_ _05195_ _05203_ _05202_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__a21bo_1
XFILLER_201_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_182_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_203_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_203_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19998_ _06922_ _06969_ _06968_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__o21ba_1
XFILLER_101_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18949_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[22\]
+ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__nand2_1
XFILLER_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_78_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_195_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21960_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[3\]\[14\]
+ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__or2_1
XFILLER_239_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20911_ _07784_ _07785_ _07760_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__a21o_1
XFILLER_215_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21891_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[3\]\[4\]
+ VGND VGND VPWR VPWR _08688_ sky130_fd_sc_hd__and2_1
XFILLER_27_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23630_ _10248_ _10249_ VGND VGND VPWR VPWR _10251_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20842_ systolic_inst.B_outs\[3\]\[7\] systolic_inst.B_shift\[3\]\[7\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__mux2_1
XFILLER_42_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23561_ _11258_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[10\] _10181_
+ _10183_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__a22o_1
X_20773_ _07678_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__inv_2
XFILLER_126_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25300_ net111 ser_C.shift_reg\[478\] VGND VGND VPWR VPWR _11120_ sky130_fd_sc_hd__and2_1
X_22512_ net65 _09240_ _09242_ systolic_inst.acc_wires\[2\]\[6\] net109 VGND VGND
+ VPWR VPWR _01816_ sky130_fd_sc_hd__a32o_1
X_26280_ clknet_leaf_25_A_in_serial_clk _00088_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_210_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23492_ systolic_inst.B_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[6\]
+ systolic_inst.B_outs\[0\]\[3\] VGND VGND VPWR VPWR _10116_ sky130_fd_sc_hd__a22oi_1
XFILLER_161_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_99_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25231_ ser_C.parallel_data\[442\] net102 net74 ser_C.shift_reg\[442\] _11085_ VGND
+ VGND VPWR VPWR _02692_ sky130_fd_sc_hd__a221o_1
X_22443_ _09096_ _09181_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__or2_1
XFILLER_183_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25162_ net110 ser_C.shift_reg\[409\] VGND VGND VPWR VPWR _11051_ sky130_fd_sc_hd__and2_1
XFILLER_109_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22374_ _09079_ _09081_ _09115_ VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__nand3_1
XFILLER_135_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24113_ systolic_inst.B_shift\[27\]\[0\] net71 _11333_ B_in\[120\] VGND VGND VPWR
+ VPWR _02098_ sky130_fd_sc_hd__a22o_1
XFILLER_191_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21325_ _08171_ _08174_ _08177_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__a21o_1
XFILLER_136_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25093_ C_out\[373\] net98 net78 ser_C.shift_reg\[373\] _11016_ VGND VGND VPWR VPWR
+ _02623_ sky130_fd_sc_hd__a221o_1
XFILLER_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24044_ _10539_ systolic_inst.B_shift\[0\]\[1\] _11332_ VGND VGND VPWR VPWR _02051_
+ sky130_fd_sc_hd__mux2_1
X_28921_ clknet_leaf_268_clk _02719_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[469\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21256_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[4\]\[1\]
+ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__nand2_1
XFILLER_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20207_ _07170_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__inv_2
X_28852_ clknet_leaf_344_clk _02650_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[400\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_133_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21187_ _07982_ _07986_ _08022_ _08020_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__o31a_1
XFILLER_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27803_ clknet_leaf_47_clk _01601_ net137 VGND VGND VPWR VPWR systolic_inst.B_outs\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_20138_ _07103_ _07105_ _07112_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25995_ systolic_inst.acc_wires\[14\]\[23\] ser_C.parallel_data\[471\] net25 VGND
+ VGND VPWR VPWR _03297_ sky130_fd_sc_hd__mux2_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28783_ clknet_leaf_230_clk _02581_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_219_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_161_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27734_ clknet_leaf_132_clk _01532_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_20069_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[6\]\[9\]
+ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__xor2_1
XFILLER_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24946_ net111 ser_C.shift_reg\[301\] VGND VGND VPWR VPWR _10943_ sky130_fd_sc_hd__and2_1
XFILLER_180_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27665_ clknet_leaf_202_clk _01463_ net147 VGND VGND VPWR VPWR systolic_inst.A_outs\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24877_ C_out\[265\] net101 net73 ser_C.shift_reg\[265\] _10908_ VGND VGND VPWR VPWR
+ _02515_ sky130_fd_sc_hd__a221o_1
XFILLER_218_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29404_ clknet_leaf_195_clk _03202_ net146 VGND VGND VPWR VPWR C_out\[376\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14630_ net69 _11792_ _11793_ systolic_inst.acc_wires\[15\]\[14\] net105 VGND VGND
+ VPWR VPWR _00992_ sky130_fd_sc_hd__a32o_1
X_23828_ net64 _10423_ _10424_ systolic_inst.acc_wires\[0\]\[20\] _11258_ VGND VGND
+ VPWR VPWR _01950_ sky130_fd_sc_hd__a32o_1
X_26616_ clknet_leaf_21_B_in_serial_clk _00419_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27596_ clknet_leaf_33_clk _01394_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_96_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29335_ clknet_leaf_218_clk _03133_ net140 VGND VGND VPWR VPWR C_out\[307\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[15\]\[5\]
+ VGND VGND VPWR VPWR _11734_ sky130_fd_sc_hd__or2_1
X_26547_ clknet_leaf_19_A_in_serial_clk _00350_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23759_ _10363_ _10365_ VGND VGND VPWR VPWR _10366_ sky130_fd_sc_hd__xor2_1
XFILLER_18_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16300_ _03679_ _03680_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__nor2_1
XFILLER_41_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13512_ deser_A.shift_reg\[76\] deser_A.shift_reg\[77\] net129 VGND VGND VPWR VPWR
+ _00349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ systolic_inst.B_outs\[10\]\[3\] systolic_inst.A_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\]
+ systolic_inst.A_outs\[10\]\[2\] VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__a22o_1
X_29266_ clknet_leaf_191_clk _03064_ net146 VGND VGND VPWR VPWR C_out\[238\] sky130_fd_sc_hd__dfrtp_1
X_26478_ clknet_leaf_13_A_in_serial_clk _00281_ net144 VGND VGND VPWR VPWR deser_A.shift_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14492_ _11671_ _11672_ VGND VGND VPWR VPWR _11673_ sky130_fd_sc_hd__and2_1
XFILLER_202_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16231_ _03611_ _03612_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__xnor2_1
XFILLER_224_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28217_ clknet_leaf_85_clk _02015_ VGND VGND VPWR VPWR systolic_inst.B_shift\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25429_ systolic_inst.A_shift\[1\]\[6\] A_in\[6\] net59 VGND VGND VPWR VPWR _11184_
+ sky130_fd_sc_hd__mux2_1
X_13443_ deser_A.shift_reg\[7\] deser_A.shift_reg\[8\] deser_A.receiving VGND VGND
+ VPWR VPWR _00280_ sky130_fd_sc_hd__mux2_1
X_29197_ clknet_leaf_141_clk _02995_ net149 VGND VGND VPWR VPWR C_out\[169\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload309 clknet_leaf_119_clk VGND VGND VPWR VPWR clkload309/Y sky130_fd_sc_hd__inv_6
XFILLER_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16162_ _03545_ _03546_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_94_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28148_ clknet_leaf_107_clk _01946_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload17 clknet_5_19__leaf_clk VGND VGND VPWR VPWR clkload17/X sky130_fd_sc_hd__clkbuf_8
XFILLER_142_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13374_ A_in\[83\] deser_A.word_buffer\[83\] net94 VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload28 clknet_leaf_332_clk VGND VGND VPWR VPWR clkload28/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_94_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload39 clknet_leaf_338_clk VGND VGND VPWR VPWR clkload39/X sky130_fd_sc_hd__clkbuf_4
X_15113_ _12228_ _12229_ VGND VGND VPWR VPWR _12230_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28079_ clknet_leaf_108_clk _01877_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_16093_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[6\]
+ systolic_inst.A_outs\[12\]\[7\] VGND VGND VPWR VPWR _13088_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_90_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19921_ _06917_ _06918_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__and2b_1
X_15044_ _12160_ _12161_ VGND VGND VPWR VPWR _12163_ sky130_fd_sc_hd__and2b_1
XFILLER_154_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19852_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[9\] _06851_ net119
+ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18803_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[8\]\[1\]
+ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__nand2_1
XFILLER_110_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19783_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] _06783_ VGND
+ VGND VPWR VPWR _06784_ sky130_fd_sc_hd__a21o_1
XFILLER_7_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_6__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_16995_ _04297_ _04298_ _04296_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__a21bo_1
XFILLER_95_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18734_ _05858_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__inv_2
X_15946_ net107 systolic_inst.acc_wires\[13\]\[29\] net67 _12966_ VGND VGND VPWR VPWR
+ _01135_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_88_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1004 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18665_ _05790_ _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_237_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ net108 systolic_inst.acc_wires\[13\]\[18\] net67 _12908_ VGND VGND VPWR VPWR
+ _01124_ sky130_fd_sc_hd__a22o_1
XFILLER_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_237_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17616_ _04856_ _04857_ _04858_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__a21o_1
XFILLER_91_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14828_ _11925_ _11952_ VGND VGND VPWR VPWR _11953_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18596_ _05722_ _05723_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__xor2_1
XFILLER_221_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17547_ systolic_inst.B_outs\[10\]\[5\] systolic_inst.B_outs\[10\]\[6\] systolic_inst.A_outs\[10\]\[7\]
+ _04797_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__a31o_1
X_14759_ _11887_ VGND VGND VPWR VPWR _11888_ sky130_fd_sc_hd__inv_2
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17478_ _04672_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19217_ _06277_ _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__xnor2_1
X_16429_ _03794_ _03795_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__nor2_1
XFILLER_203_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19148_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[7\] VGND VGND VPWR
+ VPWR _06214_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_184_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19079_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[4\]
+ systolic_inst.A_outs\[7\]\[5\] VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__and4_1
XFILLER_173_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21110_ _07913_ _07944_ _07943_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__a21boi_1
XFILLER_191_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_B_in_serial_clk clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_20_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_195_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22090_ systolic_inst.B_outs\[1\]\[4\] systolic_inst.B_shift\[1\]\[4\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__mux2_1
XFILLER_172_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21041_ _07873_ _07880_ _07879_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24800_ net112 ser_C.shift_reg\[228\] VGND VGND VPWR VPWR _10870_ sky130_fd_sc_hd__and2_1
XFILLER_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25780_ systolic_inst.acc_wires\[8\]\[0\] C_out\[256\] net22 VGND VGND VPWR VPWR
+ _03082_ sky130_fd_sc_hd__mux2_1
X_22992_ _09667_ _09668_ VGND VGND VPWR VPWR _09669_ sky130_fd_sc_hd__nand2_1
XFILLER_41_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24731_ C_out\[192\] net100 net80 ser_C.shift_reg\[192\] _10835_ VGND VGND VPWR VPWR
+ _02442_ sky130_fd_sc_hd__a221o_1
X_21943_ _08720_ _08725_ _08726_ VGND VGND VPWR VPWR _08732_ sky130_fd_sc_hd__and3_1
XFILLER_54_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27450_ clknet_leaf_235_clk _01248_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24662_ net7 ser_C.shift_reg\[159\] VGND VGND VPWR VPWR _10801_ sky130_fd_sc_hd__and2_1
XFILLER_83_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21874_ _08673_ VGND VGND VPWR VPWR _08674_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26401_ clknet_leaf_3_clk _00208_ net133 VGND VGND VPWR VPWR A_in\[69\] sky130_fd_sc_hd__dfrtp_1
X_23613_ _10231_ _10232_ VGND VGND VPWR VPWR _10234_ sky130_fd_sc_hd__xnor2_1
XFILLER_230_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20825_ _07716_ _07720_ _07721_ net60 VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_137_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27381_ clknet_leaf_340_clk _01179_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24593_ C_out\[123\] net100 net82 ser_C.shift_reg\[123\] _10766_ VGND VGND VPWR VPWR
+ _02373_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_173_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29120_ clknet_leaf_163_clk _02918_ net151 VGND VGND VPWR VPWR C_out\[92\] sky130_fd_sc_hd__dfrtp_1
X_26332_ clknet_leaf_24_clk _00139_ net137 VGND VGND VPWR VPWR A_in\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23544_ _10125_ _10128_ _10166_ VGND VGND VPWR VPWR _10167_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_98_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20756_ _07661_ _07663_ _07664_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__or3_1
XFILLER_11_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29051_ clknet_leaf_105_clk _02849_ net151 VGND VGND VPWR VPWR C_out\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26263_ clknet_leaf_5_A_in_serial_clk _00071_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23475_ _10054_ _10056_ _10097_ _10098_ VGND VGND VPWR VPWR _10100_ sky130_fd_sc_hd__o211ai_1
XFILLER_137_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20687_ _07603_ _07605_ VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__xor2_1
X_28002_ clknet_leaf_152_clk _01800_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25214_ net110 ser_C.shift_reg\[435\] VGND VGND VPWR VPWR _11077_ sky130_fd_sc_hd__and2_1
XFILLER_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22426_ _09164_ _09165_ VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__nand2b_1
X_26194_ systolic_inst.A_shift\[30\]\[0\] net71 _11333_ A_in\[120\] VGND VGND VPWR
+ VPWR _03484_ sky130_fd_sc_hd__a22o_1
XFILLER_178_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25145_ C_out\[399\] net101 net73 ser_C.shift_reg\[399\] _11042_ VGND VGND VPWR VPWR
+ _02649_ sky130_fd_sc_hd__a221o_1
XFILLER_109_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22357_ systolic_inst.A_outs\[2\]\[5\] systolic_inst.B_outs\[2\]\[6\] _11265_ systolic_inst.A_outs\[2\]\[4\]
+ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21308_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[4\]\[9\]
+ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__nor2_1
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25076_ net112 ser_C.shift_reg\[366\] VGND VGND VPWR VPWR _11008_ sky130_fd_sc_hd__and2_1
X_22288_ systolic_inst.A_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[6\] _11265_ systolic_inst.A_outs\[2\]\[2\]
+ VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_151_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24027_ systolic_inst.B_shift\[8\]\[1\] B_in\[33\] _00008_ VGND VGND VPWR VPWR _10531_
+ sky130_fd_sc_hd__mux2_1
X_28904_ clknet_leaf_271_clk _02702_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[452\]
+ sky130_fd_sc_hd__dfrtp_1
X_21239_ _08104_ _08105_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__or2_1
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28835_ clknet_leaf_236_clk _02633_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[383\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15800_ net67 _12841_ _12842_ systolic_inst.acc_wires\[13\]\[7\] net107 VGND VGND
+ VPWR VPWR _01113_ sky130_fd_sc_hd__a32o_1
X_13992_ deser_B.shift_reg\[26\] deser_B.shift_reg\[27\] net125 VGND VGND VPWR VPWR
+ _00818_ sky130_fd_sc_hd__mux2_1
X_28766_ clknet_leaf_213_clk _02564_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[314\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16780_ _04098_ _04099_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__nor2_1
X_25978_ systolic_inst.acc_wires\[14\]\[6\] ser_C.parallel_data\[454\] net24 VGND
+ VGND VPWR VPWR _03280_ sky130_fd_sc_hd__mux2_1
XFILLER_207_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27717_ clknet_leaf_188_clk _01515_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _12782_ _12781_ VGND VGND VPWR VPWR _12783_ sky130_fd_sc_hd__and2b_1
XFILLER_150_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24929_ C_out\[291\] net102 net74 ser_C.shift_reg\[291\] _10934_ VGND VGND VPWR VPWR
+ _02541_ sky130_fd_sc_hd__a221o_1
X_28697_ clknet_leaf_193_clk _02495_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[245\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18450_ systolic_inst.A_outs\[8\]\[1\] systolic_inst.B_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\]
+ systolic_inst.A_outs\[8\]\[0\] VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__a22o_1
XFILLER_73_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15662_ _12715_ VGND VGND VPWR VPWR _12716_ sky130_fd_sc_hd__inv_2
X_27648_ clknet_leaf_313_clk _01446_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_83_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17401_ _04618_ _04620_ _04656_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__a21o_1
X_14613_ _11777_ _11778_ VGND VGND VPWR VPWR _11779_ sky130_fd_sc_hd__nor2_1
X_18381_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[28\]
+ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__nand2_1
X_15593_ systolic_inst.A_outs\[13\]\[6\] _12648_ _12647_ VGND VGND VPWR VPWR _12649_
+ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_232_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27579_ clknet_leaf_218_clk _01377_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14544_ _11719_ VGND VGND VPWR VPWR _11720_ sky130_fd_sc_hd__inv_2
X_29318_ clknet_leaf_299_clk _03116_ net138 VGND VGND VPWR VPWR C_out\[290\] sky130_fd_sc_hd__dfrtp_1
X_17332_ _04589_ _04588_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__and2b_1
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29249_ clknet_leaf_184_clk _03047_ net146 VGND VGND VPWR VPWR C_out\[221\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14475_ _11623_ _11626_ _11624_ VGND VGND VPWR VPWR _11656_ sky130_fd_sc_hd__o21ba_1
X_17263_ _04496_ _04522_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__nand2_1
XFILLER_202_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19002_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[30\]
+ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__or2_1
XFILLER_179_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16214_ systolic_inst.B_outs\[12\]\[5\] systolic_inst.A_outs\[12\]\[5\] VGND VGND
+ VPWR VPWR _03597_ sky130_fd_sc_hd__nand2_1
X_13426_ deser_A.bit_idx\[2\] _11309_ _11310_ VGND VGND VPWR VPWR _11313_ sky130_fd_sc_hd__o21ai_1
X_17194_ net120 systolic_inst.B_outs\[10\]\[0\] systolic_inst.A_outs\[10\]\[0\] VGND
+ VGND VPWR VPWR _04459_ sky130_fd_sc_hd__and3_1
Xclkload106 clknet_leaf_280_clk VGND VGND VPWR VPWR clkload106/Y sky130_fd_sc_hd__clkinv_4
Xclkload117 clknet_leaf_277_clk VGND VGND VPWR VPWR clkload117/Y sky130_fd_sc_hd__inv_6
Xclkload128 clknet_leaf_263_clk VGND VGND VPWR VPWR clkload128/Y sky130_fd_sc_hd__inv_6
XFILLER_128_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16145_ _03528_ _03529_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__nor2_1
Xclkload139 clknet_leaf_254_clk VGND VGND VPWR VPWR clkload139/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_220_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13357_ A_in\[66\] deser_A.word_buffer\[66\] net96 VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__mux2_1
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16076_ _13067_ _13068_ _13070_ VGND VGND VPWR VPWR _13072_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_226_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13288_ deser_A.word_buffer\[126\] deser_A.serial_word\[126\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_226_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19904_ _06901_ _06900_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__nand2b_1
X_15027_ _12075_ _12145_ VGND VGND VPWR VPWR _12146_ sky130_fd_sc_hd__xnor2_4
XFILLER_68_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19835_ _06793_ _06795_ _06794_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__o21ba_1
XFILLER_29_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_239_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_239_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19766_ _06751_ _06767_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16978_ net69 _04288_ _04289_ systolic_inst.acc_wires\[11\]\[1\] net105 VGND VGND
+ VPWR VPWR _01235_ sky130_fd_sc_hd__a32o_1
XFILLER_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 B_in_serial_data VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_237_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18717_ _05841_ _05840_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_177_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15929_ net107 systolic_inst.acc_wires\[13\]\[26\] net67 _12952_ VGND VGND VPWR VPWR
+ _01132_ sky130_fd_sc_hd__a22o_1
XFILLER_225_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19697_ _06692_ _06700_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__nor2_1
XFILLER_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18648_ _05771_ _05774_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18579_ _05706_ _05707_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__and2b_1
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20610_ net120 _07539_ _07540_ _07521_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__a31o_1
XFILLER_166_1380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21590_ net106 _08400_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20541_ _07471_ _07472_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23260_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[29\]
+ VGND VGND VPWR VPWR _09904_ sky130_fd_sc_hd__xor2_1
XFILLER_165_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20472_ _07406_ _07405_ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__nand2b_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22211_ systolic_inst.A_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[4\]
+ systolic_inst.B_outs\[2\]\[3\] VGND VGND VPWR VPWR _08957_ sky130_fd_sc_hd__a22oi_1
XFILLER_118_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23191_ _09844_ _09845_ VGND VGND VPWR VPWR _09846_ sky130_fd_sc_hd__nand2_1
XFILLER_134_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22142_ net109 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[4\] _08890_
+ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__a21bo_1
XFILLER_173_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22073_ net65 _08842_ _08843_ systolic_inst.acc_wires\[3\]\[30\] net106 VGND VGND
+ VPWR VPWR _01776_ sky130_fd_sc_hd__a32o_1
XFILLER_133_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26950_ clknet_leaf_26_A_in_serial_clk _00748_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_236_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25901_ systolic_inst.acc_wires\[11\]\[25\] C_out\[377\] net41 VGND VGND VPWR VPWR
+ _03203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21024_ _07848_ _07857_ _07856_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_162_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26881_ clknet_leaf_9_A_in_serial_clk _00679_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28620_ clknet_leaf_215_clk _02418_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[168\]
+ sky130_fd_sc_hd__dfrtp_1
X_25832_ systolic_inst.acc_wires\[9\]\[20\] C_out\[308\] net16 VGND VGND VPWR VPWR
+ _03134_ sky130_fd_sc_hd__mux2_1
XFILLER_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28551_ clknet_leaf_173_clk _02349_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_22975_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[7\] _09625_ _09590_
+ VGND VGND VPWR VPWR _09652_ sky130_fd_sc_hd__a31o_1
X_25763_ systolic_inst.acc_wires\[7\]\[15\] C_out\[239\] net42 VGND VGND VPWR VPWR
+ _03065_ sky130_fd_sc_hd__mux2_1
XFILLER_228_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27502_ clknet_leaf_295_clk _01300_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_21926_ net106 systolic_inst.acc_wires\[3\]\[9\] net68 _08717_ VGND VGND VPWR VPWR
+ _01755_ sky130_fd_sc_hd__a22o_1
X_24714_ net113 ser_C.shift_reg\[185\] VGND VGND VPWR VPWR _10827_ sky130_fd_sc_hd__and2_1
X_28482_ clknet_leaf_108_clk _02280_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_25694_ systolic_inst.acc_wires\[5\]\[10\] C_out\[170\] net31 VGND VGND VPWR VPWR
+ _02996_ sky130_fd_sc_hd__mux2_1
XFILLER_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24645_ C_out\[149\] net104 net76 ser_C.shift_reg\[149\] _10792_ VGND VGND VPWR VPWR
+ _02399_ sky130_fd_sc_hd__a221o_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27433_ clknet_leaf_235_clk _01231_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_21857_ _08657_ _08659_ VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__nand2_1
XFILLER_19_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20808_ _07705_ _07708_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__xor2_1
XFILLER_70_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24576_ net114 ser_C.shift_reg\[116\] VGND VGND VPWR VPWR _10758_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_156_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27364_ clknet_leaf_340_clk _01162_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_21788_ _08557_ _08559_ _08558_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__o21ba_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29103_ clknet_leaf_167_clk _02901_ net152 VGND VGND VPWR VPWR C_out\[75\] sky130_fd_sc_hd__dfrtp_1
X_23527_ _10106_ _10149_ VGND VGND VPWR VPWR _10150_ sky130_fd_sc_hd__or2_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26315_ clknet_leaf_28_A_in_serial_clk _00123_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_211_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20739_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[18\]
+ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__or2_1
X_27295_ clknet_leaf_292_clk _01093_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_184_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29034_ clknet_leaf_123_clk _02832_ net144 VGND VGND VPWR VPWR C_out\[6\] sky130_fd_sc_hd__dfrtp_1
X_14260_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[7\] VGND VGND
+ VPWR VPWR _11447_ sky130_fd_sc_hd__nand2_4
X_26246_ clknet_leaf_18_A_in_serial_clk _00054_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_23458_ _10039_ _10042_ _10040_ VGND VGND VPWR VPWR _10083_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ deser_A.word_buffer\[49\] deser_A.serial_word\[49\] net128 VGND VGND VPWR
+ VPWR _00059_ sky130_fd_sc_hd__mux2_1
X_22409_ _09148_ _09149_ VGND VGND VPWR VPWR _09150_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_169_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26177_ ser_C.bit_idx\[2\] _11245_ VGND VGND VPWR VPWR _11247_ sky130_fd_sc_hd__and2_1
X_14191_ systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[3\] systolic_inst.A_outs\[15\]\[4\]
+ systolic_inst.B_outs\[15\]\[1\] VGND VGND VPWR VPWR _11380_ sky130_fd_sc_hd__a22oi_1
XFILLER_109_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23389_ _10013_ _10014_ VGND VGND VPWR VPWR _10016_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13142_ _11291_ _11292_ _11293_ VGND VGND VPWR VPWR _11295_ sky130_fd_sc_hd__or3_1
X_25128_ net110 ser_C.shift_reg\[392\] VGND VGND VPWR VPWR _11034_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25059_ C_out\[356\] net98 net78 ser_C.shift_reg\[356\] _10999_ VGND VGND VPWR VPWR
+ _02606_ sky130_fd_sc_hd__a221o_1
X_17950_ _05103_ _05106_ _05142_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__o21a_1
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_221_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16901_ _04164_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_221_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17881_ _05076_ _05075_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__nand2b_1
XFILLER_211_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19620_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[1\]\[0\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__mux2_1
XFILLER_215_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16832_ _04148_ _04149_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__xnor2_1
X_28818_ clknet_leaf_239_clk _02616_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[366\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19551_ _06584_ _06585_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__and2_1
XFILLER_24_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16763_ _04053_ _04082_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__xor2_1
X_28749_ clknet_leaf_222_clk _02547_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[297\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_234_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13975_ deser_B.shift_reg\[9\] deser_B.shift_reg\[10\] net125 VGND VGND VPWR VPWR
+ _00801_ sky130_fd_sc_hd__mux2_1
XFILLER_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18502_ systolic_inst.A_outs\[8\]\[2\] systolic_inst.B_outs\[8\]\[3\] systolic_inst.A_outs\[8\]\[3\]
+ systolic_inst.B_outs\[8\]\[4\] VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__nand4_2
XFILLER_234_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15714_ _12732_ _12735_ _12765_ VGND VGND VPWR VPWR _12767_ sky130_fd_sc_hd__o21ai_1
XFILLER_202_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19482_ _06513_ _06519_ _06521_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__o21a_1
XFILLER_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16694_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[6\] _04016_ net119
+ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18433_ net115 _05566_ _05567_ _05560_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__a31o_1
XFILLER_94_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15645_ _12698_ _12699_ VGND VGND VPWR VPWR _12700_ sky130_fd_sc_hd__nand2_1
XFILLER_234_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18364_ _05518_ _05520_ _05522_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_29_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15576_ _12615_ _12632_ VGND VGND VPWR VPWR _12633_ sky130_fd_sc_hd__xor2_1
XFILLER_159_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17315_ systolic_inst.B_outs\[10\]\[3\] systolic_inst.A_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\]
+ systolic_inst.A_outs\[10\]\[4\] VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__and4_1
X_14527_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[15\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _11705_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_25_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18295_ _05457_ _05460_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__a21oi_1
XFILLER_222_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17246_ systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[5\]
+ systolic_inst.B_outs\[10\]\[0\] VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_228_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14458_ _11588_ _11638_ VGND VGND VPWR VPWR _11640_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_228_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_228_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13409_ A_in\[118\] deser_A.word_buffer\[118\] net92 VGND VGND VPWR VPWR _00257_
+ sky130_fd_sc_hd__mux2_1
X_17177_ _04458_ _04457_ systolic_inst.acc_wires\[11\]\[31\] net105 VGND VGND VPWR
+ VPWR _01265_ sky130_fd_sc_hd__a2bb2o_1
X_14389_ _11556_ _11572_ VGND VGND VPWR VPWR _11573_ sky130_fd_sc_hd__xor2_1
XFILLER_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16128_ _13057_ _13093_ _13091_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__a21o_1
XFILLER_227_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_291_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_291_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_103_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16059_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[3\] _13038_ _13037_
+ VGND VGND VPWR VPWR _13055_ sky130_fd_sc_hd__a31o_1
XFILLER_233_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19818_ net106 _06818_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__nor2_1
XFILLER_84_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19749_ _06714_ _06750_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22760_ _09442_ _09443_ VGND VGND VPWR VPWR _09444_ sky130_fd_sc_hd__nor2_1
XFILLER_77_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21711_ systolic_inst.B_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[6\] systolic_inst.A_outs\[3\]\[7\]
+ systolic_inst.B_outs\[3\]\[3\] VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__a22o_1
XFILLER_164_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22691_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.A_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\]
+ systolic_inst.A_outs\[1\]\[1\] VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__and4_1
XFILLER_240_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24430_ net114 ser_C.shift_reg\[43\] VGND VGND VPWR VPWR _10685_ sky130_fd_sc_hd__and2_1
X_21642_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[6\] VGND VGND VPWR
+ VPWR _08451_ sky130_fd_sc_hd__nand2_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24361_ C_out\[7\] net104 _10643_ ser_C.shift_reg\[7\] _10650_ VGND VGND VPWR VPWR
+ _02257_ sky130_fd_sc_hd__a221o_1
XFILLER_177_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_20 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21573_ _08382_ _08383_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__or2_1
XANTENNA_31 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26100_ deser_B.serial_word\[55\] deser_B.shift_reg\[55\] net56 VGND VGND VPWR VPWR
+ _03402_ sky130_fd_sc_hd__mux2_1
XANTENNA_42 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23312_ _09919_ _09927_ _09939_ _09940_ VGND VGND VPWR VPWR _09942_ sky130_fd_sc_hd__a22o_1
X_20524_ _07455_ _07457_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27080_ clknet_leaf_28_B_in_serial_clk _00878_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24292_ _10619_ systolic_inst.A_shift\[11\]\[1\] net71 VGND VGND VPWR VPWR _02219_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26031_ systolic_inst.acc_wires\[15\]\[27\] ser_C.parallel_data\[507\] net37 VGND
+ VGND VPWR VPWR _03333_ sky130_fd_sc_hd__mux2_1
X_23243_ _09888_ _09889_ VGND VGND VPWR VPWR _09890_ sky130_fd_sc_hd__nand2_1
XFILLER_181_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20455_ _07387_ _07388_ _07389_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__a21oi_1
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23174_ _09821_ _09826_ _09830_ _11713_ VGND VGND VPWR VPWR _09832_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_164_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20386_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[7\]
+ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__o21a_1
XFILLER_84_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22125_ systolic_inst.A_outs\[2\]\[1\] systolic_inst.B_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\]
+ systolic_inst.A_outs\[2\]\[0\] VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_282_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_282_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27982_ clknet_leaf_118_clk _01780_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_216_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22056_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[28\]
+ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__and2_2
XFILLER_173_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26933_ clknet_leaf_21_A_in_serial_clk _00731_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21007_ _07874_ _07878_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__or2_1
XFILLER_212_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29652_ clknet_leaf_5_B_in_serial_clk _03447_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26864_ clknet_leaf_31_B_in_serial_clk net56 net134 VGND VGND VPWR VPWR deser_B.serial_word_ready
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_60_1340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28603_ clknet_leaf_136_clk _02401_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[151\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25815_ systolic_inst.acc_wires\[9\]\[3\] C_out\[291\] net14 VGND VGND VPWR VPWR
+ _03117_ sky130_fd_sc_hd__mux2_1
X_29583_ clknet_leaf_19_B_in_serial_clk _03378_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26795_ clknet_leaf_85_clk _00597_ net153 VGND VGND VPWR VPWR B_in\[67\] sky130_fd_sc_hd__dfrtp_1
XFILLER_169_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap11 net12 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_6
Xmax_cap22 net29 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_8
XFILLER_228_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28534_ clknet_leaf_161_clk _02332_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[82\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap33 net54 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_8
X_13760_ B_in\[67\] deser_B.word_buffer\[67\] net87 VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__mux2_1
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap44 net46 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_8
X_22958_ _09627_ _09635_ VGND VGND VPWR VPWR _09636_ sky130_fd_sc_hd__nand2_1
X_25746_ systolic_inst.acc_wires\[6\]\[30\] C_out\[222\] net43 VGND VGND VPWR VPWR
+ _03048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap55 _00001_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_104_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap66 net68 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_12
XFILLER_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21909_ _08694_ _08698_ _08700_ _08702_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__o211a_1
Xmax_cap77 net80 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_12
Xmax_cap88 net90 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_6
X_28465_ clknet_leaf_100_clk _02263_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13691_ deser_B.word_buffer\[127\] deser_B.serial_word\[127\] net123 VGND VGND VPWR
+ VPWR _00528_ sky130_fd_sc_hd__mux2_1
Xmax_cap99 net100 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_12
X_22889_ _09566_ _09567_ VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__xnor2_1
X_25677_ systolic_inst.acc_wires\[4\]\[25\] C_out\[153\] net30 VGND VGND VPWR VPWR
+ _02979_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27416_ clknet_leaf_214_clk _01214_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15430_ systolic_inst.A_outs\[13\]\[2\] systolic_inst.B_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\]
+ systolic_inst.A_outs\[13\]\[1\] VGND VGND VPWR VPWR _12491_ sky130_fd_sc_hd__a22o_1
X_24628_ net7 ser_C.shift_reg\[142\] VGND VGND VPWR VPWR _10784_ sky130_fd_sc_hd__and2_1
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28396_ clknet_leaf_33_clk _02194_ VGND VGND VPWR VPWR systolic_inst.A_shift\[16\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ systolic_inst.A_outs\[13\]\[5\] systolic_inst.A_outs\[12\]\[5\] net115 VGND
+ VGND VPWR VPWR _01079_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24559_ C_out\[106\] net99 net80 ser_C.shift_reg\[106\] _10749_ VGND VGND VPWR VPWR
+ _02356_ sky130_fd_sc_hd__a221o_1
XFILLER_200_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27347_ clknet_leaf_342_clk _01145_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_196_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17100_ net105 systolic_inst.acc_wires\[11\]\[19\] net62 _04393_ VGND VGND VPWR VPWR
+ _01253_ sky130_fd_sc_hd__a22o_1
XFILLER_106_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14312_ _11496_ _11497_ VGND VGND VPWR VPWR _11498_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_78_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15292_ _12384_ _12383_ systolic_inst.acc_wires\[14\]\[21\] net107 VGND VGND VPWR
+ VPWR _01063_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18080_ _05267_ _05268_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__xnor2_1
X_27278_ clknet_leaf_326_clk _01076_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_237_Right_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29017_ clknet_leaf_94_clk _02815_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _11428_ _11429_ _11397_ _11399_ VGND VGND VPWR VPWR _11431_ sky130_fd_sc_hd__o211ai_1
X_17031_ _04330_ _04332_ _04334_ systolic_inst.acc_wires\[11\]\[9\] net105 VGND VGND
+ VPWR VPWR _01243_ sky130_fd_sc_hd__a32o_1
X_26229_ clknet_leaf_7_A_in_serial_clk _00037_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_31__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_31__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_223_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14174_ _11347_ _11362_ VGND VGND VPWR VPWR _11364_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_223_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_273_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_273_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13125_ net130 deser_A.bit_idx\[1\] deser_A.bit_idx\[0\] deser_A.bit_idx\[2\] VGND
+ VGND VPWR VPWR _11280_ sky130_fd_sc_hd__and4_1
XFILLER_98_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18982_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[27\]
+ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17933_ _05093_ _05125_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17864_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[3\] VGND VGND VPWR
+ VPWR _05060_ sky130_fd_sc_hd__nand2_1
XFILLER_121_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19603_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[30\]
+ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__or2_1
XFILLER_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16815_ _04097_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__xor2_1
XFILLER_238_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17795_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.B_outs\[4\]\[2\] net121 VGND
+ VGND VPWR VPWR _01340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19534_ net105 systolic_inst.acc_wires\[7\]\[19\] net62 _06571_ VGND VGND VPWR VPWR
+ _01509_ sky130_fd_sc_hd__a22o_1
X_16746_ systolic_inst.A_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[5\] VGND VGND
+ VPWR VPWR _04067_ sky130_fd_sc_hd__nand2_1
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13958_ deser_A.serial_word\[119\] deser_A.shift_reg\[119\] _00002_ VGND VGND VPWR
+ VPWR _00784_ sky130_fd_sc_hd__mux2_1
XFILLER_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19465_ _06508_ _06510_ _06512_ systolic_inst.acc_wires\[7\]\[9\] net105 VGND VGND
+ VPWR VPWR _01499_ sky130_fd_sc_hd__a32o_1
XFILLER_179_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16677_ systolic_inst.A_outs\[11\]\[1\] systolic_inst.B_outs\[11\]\[6\] VGND VGND
+ VPWR VPWR _04000_ sky130_fd_sc_hd__nand2_1
X_13889_ deser_A.serial_word\[50\] deser_A.shift_reg\[50\] net58 VGND VGND VPWR VPWR
+ _00715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18416_ systolic_inst.B_outs\[7\]\[5\] systolic_inst.B_outs\[3\]\[5\] net119 VGND
+ VGND VPWR VPWR _01407_ sky130_fd_sc_hd__mux2_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15628_ _12577_ _12681_ VGND VGND VPWR VPWR _12683_ sky130_fd_sc_hd__nand2_1
XFILLER_61_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19396_ _06376_ _06439_ _06437_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18347_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[23\]
+ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__xor2_1
XFILLER_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15559_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[7\] VGND VGND
+ VPWR VPWR _12616_ sky130_fd_sc_hd__nand2_4
XFILLER_188_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18278_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[9\]\[13\]
+ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__or2_1
XFILLER_175_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_204_Right_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17229_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.A_outs\[10\]\[4\] VGND VGND
+ VPWR VPWR _04490_ sky130_fd_sc_hd__nand2_1
XFILLER_162_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20240_ net109 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[0\] _07184_
+ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__a21o_1
XFILLER_157_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_264_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_264_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20171_ net62 _07139_ _07140_ systolic_inst.acc_wires\[6\]\[23\] net106 VGND VGND
+ VPWR VPWR _01577_ sky130_fd_sc_hd__a32o_1
XFILLER_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23930_ systolic_inst.A_shift\[3\]\[2\] net72 _11333_ A_in\[26\] VGND VGND VPWR VPWR
+ _01980_ sky130_fd_sc_hd__a22o_1
XFILLER_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_198_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23861_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[26\]
+ VGND VGND VPWR VPWR _10452_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_198_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25600_ systolic_inst.acc_wires\[2\]\[12\] C_out\[76\] net51 VGND VGND VPWR VPWR
+ _02902_ sky130_fd_sc_hd__mux2_1
X_22812_ _09428_ _09461_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[7\]
+ VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_140_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23792_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[15\]
+ VGND VGND VPWR VPWR _10394_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_140_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26580_ clknet_leaf_28_A_in_serial_clk _00383_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22743_ _09410_ _09426_ VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__xor2_1
X_25531_ systolic_inst.acc_wires\[0\]\[7\] C_out\[7\] net33 VGND VGND VPWR VPWR _02833_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25462_ _11204_ _11205_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__and2_1
XFILLER_213_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28250_ clknet_leaf_96_clk _02048_ VGND VGND VPWR VPWR systolic_inst.B_shift\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_22674_ systolic_inst.A_outs\[1\]\[1\] systolic_inst.A_outs\[0\]\[1\] net121 VGND
+ VGND VPWR VPWR _01843_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24413_ C_out\[33\] _11302_ net81 ser_C.shift_reg\[33\] _10676_ VGND VGND VPWR VPWR
+ _02283_ sky130_fd_sc_hd__a221o_1
XFILLER_213_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27201_ clknet_leaf_262_clk _00999_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_21625_ _08402_ _08434_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__nand2b_1
XFILLER_205_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28181_ clknet_leaf_63_clk _01979_ VGND VGND VPWR VPWR systolic_inst.A_shift\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25393_ systolic_inst.A_shift\[3\]\[4\] A_in\[20\] net59 VGND VGND VPWR VPWR _11166_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27132_ clknet_leaf_71_clk _00930_ VGND VGND VPWR VPWR systolic_inst.B_shift\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24344_ systolic_inst.A_shift\[8\]\[7\] net70 net83 systolic_inst.A_shift\[9\]\[7\]
+ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__a22o_1
XFILLER_205_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21556_ _08345_ _08367_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__nand2b_1
XFILLER_21_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27063_ clknet_leaf_6_B_in_serial_clk _00861_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[69\]
+ sky130_fd_sc_hd__dfrtp_1
X_20507_ _07401_ _07403_ _07402_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__o21ba_1
XFILLER_165_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24275_ systolic_inst.B_shift\[27\]\[1\] B_in\[89\] net59 VGND VGND VPWR VPWR _10611_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21487_ systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[1\] VGND VGND VPWR
+ VPWR _08302_ sky130_fd_sc_hd__nand2_1
XFILLER_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26014_ systolic_inst.acc_wires\[15\]\[10\] ser_C.parallel_data\[490\] net39 VGND
+ VGND VPWR VPWR _03316_ sky130_fd_sc_hd__mux2_1
X_23226_ net65 _09874_ _09875_ systolic_inst.acc_wires\[1\]\[23\] net109 VGND VGND
+ VPWR VPWR _01897_ sky130_fd_sc_hd__a32o_1
XFILLER_181_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20438_ systolic_inst.A_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[5\] _07336_ _07335_
+ VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__a31oi_1
XFILLER_49_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_255_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_255_clk
+ sky130_fd_sc_hd__clkbuf_8
X_23157_ _09808_ _09809_ _09816_ VGND VGND VPWR VPWR _09817_ sky130_fd_sc_hd__a21o_1
XFILLER_136_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20369_ _07294_ _07306_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__or2_1
XFILLER_122_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22108_ net122 _08857_ _08858_ _08851_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__a31o_1
XFILLER_175_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23088_ _09755_ _09756_ _09757_ VGND VGND VPWR VPWR _09758_ sky130_fd_sc_hd__a21o_1
X_27965_ clknet_leaf_165_clk _01763_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_62_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22039_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[26\]
+ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__or2_1
X_14930_ _12050_ _12051_ VGND VGND VPWR VPWR _12052_ sky130_fd_sc_hd__xnor2_1
X_26916_ clknet_leaf_10_A_in_serial_clk _00714_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_27896_ clknet_leaf_39_clk _01694_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29635_ clknet_leaf_26_B_in_serial_clk _03430_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26847_ clknet_leaf_68_clk _00649_ net135 VGND VGND VPWR VPWR B_in\[119\] sky130_fd_sc_hd__dfrtp_1
X_14861_ _11953_ _11956_ _11983_ _11984_ VGND VGND VPWR VPWR _11985_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_67_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _03925_ _03926_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__or2_1
X_13812_ B_in\[119\] deser_B.word_buffer\[119\] net87 VGND VGND VPWR VPWR _00649_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29566_ clknet_leaf_16_B_in_serial_clk _03361_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17580_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[10\]\[1\]
+ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__or2_1
X_26778_ clknet_leaf_52_clk _00580_ net143 VGND VGND VPWR VPWR B_in\[50\] sky130_fd_sc_hd__dfrtp_1
X_14792_ _11917_ VGND VGND VPWR VPWR _11918_ sky130_fd_sc_hd__inv_2
XFILLER_235_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28517_ clknet_leaf_155_clk _02315_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_16531_ _03863_ _03881_ _03883_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_63_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13743_ B_in\[50\] deser_B.word_buffer\[50\] net86 VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__mux2_1
X_25729_ systolic_inst.acc_wires\[6\]\[13\] C_out\[205\] net45 VGND VGND VPWR VPWR
+ _03031_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_119_Left_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29497_ clknet_5_8__leaf_clk _03295_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[469\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19250_ systolic_inst.B_outs\[7\]\[5\] systolic_inst.A_outs\[7\]\[5\] VGND VGND VPWR
+ VPWR _06313_ sky130_fd_sc_hd__nand2_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16462_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[12\]\[14\]
+ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__nand2_1
XFILLER_32_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28448_ clknet_leaf_34_clk _02246_ VGND VGND VPWR VPWR systolic_inst.A_shift\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13674_ deser_B.word_buffer\[110\] deser_B.serial_word\[110\] net123 VGND VGND VPWR
+ VPWR _00511_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18201_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[9\]\[2\]
+ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__and2_1
X_15413_ _12467_ _12473_ _12474_ VGND VGND VPWR VPWR _12475_ sky130_fd_sc_hd__and3_1
X_19181_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[6\] VGND VGND VPWR
+ VPWR _06246_ sky130_fd_sc_hd__nand2_1
XFILLER_223_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16393_ _03757_ _03760_ _03762_ _03764_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__o211a_1
X_28379_ clknet_leaf_31_clk _02177_ VGND VGND VPWR VPWR systolic_inst.A_shift\[19\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_18132_ systolic_inst.B_outs\[9\]\[6\] systolic_inst.A_outs\[9\]\[7\] VGND VGND VPWR
+ VPWR _05320_ sky130_fd_sc_hd__nand2_1
XFILLER_185_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15344_ systolic_inst.acc_wires\[14\]\[28\] systolic_inst.acc_wires\[14\]\[29\] systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12428_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_136_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18063_ _05252_ _05253_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__nand2b_1
X_15275_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[19\]
+ VGND VGND VPWR VPWR _12370_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_97_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17014_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[11\]\[7\]
+ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__nand2_1
XFILLER_176_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14226_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[6\] _11411_ _11412_
+ VGND VGND VPWR VPWR _11414_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_128_Left_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_246_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_246_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_193_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14157_ _11346_ _11347_ VGND VGND VPWR VPWR _11348_ sky130_fd_sc_hd__nand2_1
XFILLER_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_242_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_242_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13108_ systolic_inst.B_outs\[14\]\[7\] VGND VGND VPWR VPWR _11264_ sky130_fd_sc_hd__inv_2
X_14088_ deser_B.shift_reg\[122\] deser_B.shift_reg\[123\] deser_B.receiving VGND
+ VGND VPWR VPWR _00914_ sky130_fd_sc_hd__mux2_1
X_18965_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[24\]
+ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17916_ _05087_ _05089_ _05088_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__o21ba_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18896_ _05994_ _05998_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__and2_1
XFILLER_239_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_201_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17847_ _05021_ _05024_ _05043_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__a21o_1
XFILLER_54_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_137_Left_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17778_ _04993_ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_193_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19517_ net60 _06557_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__nor2_1
XFILLER_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16729_ _03983_ _03984_ _04015_ _04013_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__a31o_1
XFILLER_23_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19448_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[7\]\[7\]
+ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19379_ _06411_ _06413_ _06436_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__and3_1
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21410_ _08251_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__inv_2
XFILLER_202_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22390_ systolic_inst.B_outs\[2\]\[5\] systolic_inst.A_outs\[2\]\[7\] _09129_ VGND
+ VGND VPWR VPWR _09131_ sky130_fd_sc_hd__and3_1
XFILLER_176_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21341_ _08191_ _08192_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__nand2_1
XFILLER_11_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_187_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24060_ _10547_ systolic_inst.B_shift\[15\]\[1\] net70 VGND VGND VPWR VPWR _02059_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_208_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21272_ _08132_ _08133_ _08125_ _08129_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_208_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_208_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23011_ systolic_inst.A_outs\[1\]\[6\] _11277_ VGND VGND VPWR VPWR _09687_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_237_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_237_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20223_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.A_outs\[4\]\[0\] net116 VGND
+ VGND VPWR VPWR _01586_ sky130_fd_sc_hd__mux2_1
XFILLER_190_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_146_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20154_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[21\]
+ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_146_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27750_ clknet_leaf_209_clk _01548_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20085_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[6\]\[11\]
+ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24962_ net111 ser_C.shift_reg\[309\] VGND VGND VPWR VPWR _10951_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_5_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26701_ clknet_leaf_6_B_in_serial_clk _00504_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23913_ _10489_ systolic_inst.B_shift\[18\]\[0\] _11332_ VGND VGND VPWR VPWR _01970_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27681_ clknet_leaf_200_clk _01479_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24893_ C_out\[273\] net103 net75 ser_C.shift_reg\[273\] _10916_ VGND VGND VPWR VPWR
+ _02523_ sky130_fd_sc_hd__a221o_1
X_29420_ clknet_leaf_334_clk _03218_ net131 VGND VGND VPWR VPWR C_out\[392\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26632_ clknet_leaf_18_B_in_serial_clk _00435_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_23844_ _10429_ _10433_ _10435_ _11713_ VGND VGND VPWR VPWR _10438_ sky130_fd_sc_hd__a31o_1
XFILLER_217_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29351_ clknet_leaf_228_clk _03149_ net138 VGND VGND VPWR VPWR C_out\[323\] sky130_fd_sc_hd__dfrtp_1
X_23775_ _10378_ _10379_ VGND VGND VPWR VPWR _10380_ sky130_fd_sc_hd__nor2_1
XFILLER_26_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26563_ clknet_leaf_27_A_in_serial_clk _00366_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20987_ _07859_ _07860_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__nand2_1
XFILLER_214_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28302_ clknet_leaf_66_clk _02100_ VGND VGND VPWR VPWR systolic_inst.B_shift\[27\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25514_ _11237_ _11238_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__and2b_1
XFILLER_198_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22726_ _09391_ _09408_ _09410_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__and3_1
X_29282_ clknet_leaf_184_clk _03080_ net146 VGND VGND VPWR VPWR C_out\[254\] sky130_fd_sc_hd__dfrtp_1
X_26494_ clknet_leaf_7_A_in_serial_clk _00297_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_241_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28233_ clknet_leaf_130_clk _02031_ VGND VGND VPWR VPWR systolic_inst.B_shift\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22657_ _09364_ VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__inv_2
X_25445_ systolic_inst.cycle_cnt\[4\] _11279_ _11191_ VGND VGND VPWR VPWR _11194_
+ sky130_fd_sc_hd__a21o_1
XFILLER_199_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21608_ systolic_inst.A_outs\[3\]\[2\] systolic_inst.B_outs\[3\]\[5\] VGND VGND VPWR
+ VPWR _08418_ sky130_fd_sc_hd__nand2_1
XFILLER_138_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28164_ clknet_leaf_95_clk _01962_ VGND VGND VPWR VPWR systolic_inst.B_shift\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13390_ A_in\[99\] deser_A.word_buffer\[99\] _00003_ VGND VGND VPWR VPWR _00238_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22588_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[18\]
+ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__or2_1
XFILLER_223_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25376_ _11157_ systolic_inst.B_shift\[14\]\[3\] net71 VGND VGND VPWR VPWR _02765_
+ sky130_fd_sc_hd__mux2_1
XFILLER_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27115_ clknet_leaf_31_B_in_serial_clk _00913_ net134 VGND VGND VPWR VPWR deser_B.shift_reg\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21539_ _08346_ _08349_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24327_ systolic_inst.A_shift\[10\]\[3\] A_in\[35\] net59 VGND VGND VPWR VPWR _10637_
+ sky130_fd_sc_hd__mux2_1
X_28095_ clknet_leaf_113_clk _01893_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15060_ systolic_inst.B_outs\[14\]\[6\] systolic_inst.A_outs\[14\]\[6\] _11264_ systolic_inst.A_outs\[14\]\[5\]
+ VGND VGND VPWR VPWR _12178_ sky130_fd_sc_hd__o2bb2a_1
X_27046_ clknet_leaf_25_B_in_serial_clk _00844_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_24258_ systolic_inst.A_shift\[16\]\[1\] net70 net83 systolic_inst.A_shift\[17\]\[1\]
+ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__a22o_1
XFILLER_175_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14011_ deser_B.shift_reg\[45\] deser_B.shift_reg\[46\] net125 VGND VGND VPWR VPWR
+ _00837_ sky130_fd_sc_hd__mux2_1
XFILLER_49_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23209_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[21\]
+ VGND VGND VPWR VPWR _09861_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_228_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_228_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_175_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24189_ systolic_inst.A_shift\[24\]\[4\] net70 _10505_ systolic_inst.A_shift\[25\]\[4\]
+ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28997_ clknet_leaf_105_clk _02795_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18750_ _05806_ _05872_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__or2_1
XFILLER_237_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27948_ clknet_leaf_178_clk _01746_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15962_ systolic_inst.A_outs\[12\]\[3\] systolic_inst.A_shift\[24\]\[3\] net115 VGND
+ VGND VPWR VPWR _01141_ sky130_fd_sc_hd__mux2_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17701_ _04922_ _04924_ _04931_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__a21oi_1
XFILLER_76_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14913_ _12028_ _12034_ VGND VGND VPWR VPWR _12035_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18681_ systolic_inst.B_outs\[8\]\[5\] systolic_inst.A_outs\[8\]\[6\] VGND VGND VPWR
+ VPWR _05807_ sky130_fd_sc_hd__nand2_1
X_27879_ clknet_leaf_39_clk _01677_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15893_ _12913_ _12919_ _12920_ VGND VGND VPWR VPWR _12922_ sky130_fd_sc_hd__a21oi_1
X_29618_ clknet_leaf_4_B_in_serial_clk _03413_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17632_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[10\]\[8\]
+ _04869_ _04871_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__a211o_1
XFILLER_224_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14844_ _11966_ _11967_ VGND VGND VPWR VPWR _11968_ sky130_fd_sc_hd__or2_1
XFILLER_91_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29549_ clknet_leaf_230_clk _03344_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_17563_ _04763_ _04792_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__nor2_1
XFILLER_217_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14775_ systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[3\] VGND VGND
+ VPWR VPWR _11902_ sky130_fd_sc_hd__nand2_1
XFILLER_44_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19302_ _06363_ _06362_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__and2b_1
XFILLER_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_A_in_serial_clk clknet_2_0__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_0_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16514_ net108 systolic_inst.acc_wires\[12\]\[21\] net67 _03869_ VGND VGND VPWR VPWR
+ _01191_ sky130_fd_sc_hd__a22o_1
XFILLER_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13726_ B_in\[33\] deser_B.word_buffer\[33\] net86 VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__mux2_1
XFILLER_17_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17494_ systolic_inst.B_outs\[10\]\[5\] systolic_inst.A_outs\[10\]\[7\] _04745_ VGND
+ VGND VPWR VPWR _04747_ sky130_fd_sc_hd__and3_1
XFILLER_143_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19233_ _06294_ _06295_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__xnor2_1
X_16445_ _03794_ _03801_ _03802_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__a21bo_1
XFILLER_204_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13657_ deser_B.word_buffer\[93\] deser_B.serial_word\[93\] net123 VGND VGND VPWR
+ VPWR _00494_ sky130_fd_sc_hd__mux2_1
XFILLER_32_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19164_ _06198_ _06229_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__and2b_1
XFILLER_169_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16376_ _03750_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__inv_2
X_13588_ deser_B.word_buffer\[24\] deser_B.serial_word\[24\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18115_ _05302_ _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__nand2_1
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15327_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[27\]
+ VGND VGND VPWR VPWR _12414_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_41_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19095_ _06144_ _06162_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__nand2b_1
XFILLER_117_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18046_ _05235_ _05236_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__nand2_1
X_15258_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[16\]
+ VGND VGND VPWR VPWR _12356_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_219_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_219_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14209_ _11370_ _11396_ VGND VGND VPWR VPWR _11398_ sky130_fd_sc_hd__xor2_1
XFILLER_67_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15189_ _12296_ VGND VGND VPWR VPWR _12297_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_182_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19997_ _06922_ _06991_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__xnor2_1
XFILLER_28_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18948_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[22\]
+ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__or2_1
XFILLER_230_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_195_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18879_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[8\]\[12\]
+ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__or2_1
XFILLER_227_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20910_ _07760_ _07784_ _07785_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__nand3_1
XFILLER_67_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21890_ net65 _08685_ _08687_ systolic_inst.acc_wires\[3\]\[3\] net106 VGND VGND
+ VPWR VPWR _01749_ sky130_fd_sc_hd__a32o_1
XFILLER_94_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20841_ systolic_inst.B_outs\[3\]\[6\] systolic_inst.B_shift\[3\]\[6\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__mux2_1
XFILLER_39_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23560_ _11258_ _10182_ VGND VGND VPWR VPWR _10183_ sky130_fd_sc_hd__nor2_1
XFILLER_39_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20772_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[23\]
+ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__xor2_1
X_22511_ _09241_ VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__inv_2
XFILLER_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23491_ systolic_inst.B_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[5\]
+ systolic_inst.A_outs\[0\]\[6\] VGND VGND VPWR VPWR _10115_ sky130_fd_sc_hd__and4_1
XFILLER_210_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22442_ systolic_inst.B_outs\[2\]\[5\] systolic_inst.B_outs\[2\]\[6\] systolic_inst.A_outs\[2\]\[7\]
+ _09180_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__a31o_1
X_25230_ net111 ser_C.shift_reg\[443\] VGND VGND VPWR VPWR _11085_ sky130_fd_sc_hd__and2_1
XFILLER_195_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25161_ C_out\[407\] net101 net73 ser_C.shift_reg\[407\] _11050_ VGND VGND VPWR VPWR
+ _02657_ sky130_fd_sc_hd__a221o_1
XFILLER_202_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22373_ _09056_ _09114_ VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24112_ systolic_inst.B_shift\[1\]\[7\] _11332_ net83 systolic_inst.B_shift\[5\]\[7\]
+ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__a22o_1
X_21324_ _08171_ _08174_ _08177_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__nand3_1
XFILLER_50_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25092_ net113 ser_C.shift_reg\[374\] VGND VGND VPWR VPWR _11016_ sky130_fd_sc_hd__and2_1
XFILLER_163_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24043_ systolic_inst.B_shift\[4\]\[1\] B_in\[1\] _00008_ VGND VGND VPWR VPWR _10539_
+ sky130_fd_sc_hd__mux2_1
XFILLER_117_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28920_ clknet_leaf_282_clk _02718_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_116_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21255_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[4\]\[1\]
+ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__and2_1
XFILLER_144_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20206_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[29\]
+ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__xor2_1
XFILLER_46_1227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28851_ clknet_leaf_344_clk _02649_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[399\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21186_ _08054_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__inv_2
XFILLER_81_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27802_ clknet_leaf_47_clk _01600_ net137 VGND VGND VPWR VPWR systolic_inst.B_outs\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20137_ systolic_inst.acc_wires\[6\]\[16\] systolic_inst.acc_wires\[6\]\[17\] systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__o21a_1
X_28782_ clknet_leaf_230_clk _02580_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[330\]
+ sky130_fd_sc_hd__dfrtp_1
X_25994_ systolic_inst.acc_wires\[14\]\[22\] ser_C.parallel_data\[470\] net25 VGND
+ VGND VPWR VPWR _03296_ sky130_fd_sc_hd__mux2_1
XFILLER_58_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27733_ clknet_leaf_132_clk _01531_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_20068_ _07052_ _07051_ systolic_inst.acc_wires\[6\]\[8\] net106 VGND VGND VPWR VPWR
+ _01562_ sky130_fd_sc_hd__a2bb2o_1
X_24945_ C_out\[299\] net103 net76 ser_C.shift_reg\[299\] _10942_ VGND VGND VPWR VPWR
+ _02549_ sky130_fd_sc_hd__a221o_1
XFILLER_219_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27664_ clknet_leaf_202_clk _01462_ net147 VGND VGND VPWR VPWR systolic_inst.A_outs\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_46_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24876_ net110 ser_C.shift_reg\[266\] VGND VGND VPWR VPWR _10908_ sky130_fd_sc_hd__and2_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29403_ clknet_leaf_238_clk _03201_ net146 VGND VGND VPWR VPWR C_out\[375\] sky130_fd_sc_hd__dfrtp_1
X_26615_ clknet_leaf_17_B_in_serial_clk _00418_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_23827_ _10421_ _10422_ _10419_ VGND VGND VPWR VPWR _10424_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27595_ clknet_leaf_224_clk _01393_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29334_ clknet_leaf_218_clk _03132_ net140 VGND VGND VPWR VPWR C_out\[306\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[15\]\[5\]
+ VGND VGND VPWR VPWR _11733_ sky130_fd_sc_hd__nand2_1
XFILLER_72_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26546_ clknet_leaf_20_A_in_serial_clk _00349_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_220_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23758_ _10358_ _10364_ VGND VGND VPWR VPWR _10365_ sky130_fd_sc_hd__nand2_1
XFILLER_202_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13511_ deser_A.shift_reg\[75\] deser_A.shift_reg\[76\] net129 VGND VGND VPWR VPWR
+ _00348_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22709_ _09384_ _09393_ _09394_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__nand3_1
X_29265_ clknet_leaf_198_clk _03063_ net146 VGND VGND VPWR VPWR C_out\[237\] sky130_fd_sc_hd__dfrtp_1
XFILLER_144_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26477_ clknet_leaf_13_A_in_serial_clk _00280_ net143 VGND VGND VPWR VPWR deser_A.shift_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14491_ _11637_ _11639_ _11670_ VGND VGND VPWR VPWR _11672_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_81_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23689_ _10305_ _10306_ VGND VGND VPWR VPWR _10307_ sky130_fd_sc_hd__nand2_1
X_28216_ clknet_leaf_85_clk _02014_ VGND VGND VPWR VPWR systolic_inst.B_shift\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16230_ _03612_ _03611_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_133_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13442_ deser_A.shift_reg\[6\] deser_A.shift_reg\[7\] deser_A.receiving VGND VGND
+ VPWR VPWR _00279_ sky130_fd_sc_hd__mux2_1
X_25428_ _11183_ systolic_inst.A_shift\[0\]\[5\] net70 VGND VGND VPWR VPWR _02791_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29196_ clknet_leaf_141_clk _02994_ net149 VGND VGND VPWR VPWR C_out\[168\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28147_ clknet_leaf_100_clk _01945_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_16161_ _03504_ _03506_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__and2_1
X_13373_ A_in\[82\] deser_A.word_buffer\[82\] net95 VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25359_ ser_C.parallel_data\[506\] net98 net78 ser_C.shift_reg\[506\] _11149_ VGND
+ VGND VPWR VPWR _02756_ sky130_fd_sc_hd__a221o_1
Xclkload18 clknet_5_20__leaf_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_94_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload29 clknet_leaf_334_clk VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_94_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15112_ _12199_ _12203_ VGND VGND VPWR VPWR _12229_ sky130_fd_sc_hd__nor2_1
X_28078_ clknet_leaf_108_clk _01876_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16092_ systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[6\] systolic_inst.A_outs\[12\]\[7\]
+ systolic_inst.B_outs\[12\]\[0\] VGND VGND VPWR VPWR _13087_ sky130_fd_sc_hd__a22o_1
XFILLER_177_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27029_ clknet_leaf_11_B_in_serial_clk _00827_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_182_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19920_ _06883_ _06888_ _06914_ _06915_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__a211o_1
X_15043_ _12161_ _12160_ VGND VGND VPWR VPWR _12162_ sky130_fd_sc_hd__and2b_1
XFILLER_5_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19851_ _06849_ _06850_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_9_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18802_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[8\]\[1\]
+ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__and2_1
X_19782_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[7\]
+ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__o21ai_2
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16994_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[11\]\[4\]
+ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__or2_1
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18733_ _05855_ _05857_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__nand2_1
XFILLER_95_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15945_ _12963_ _12965_ VGND VGND VPWR VPWR _12966_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18664_ _05730_ _05755_ _05754_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__a21boi_1
XFILLER_110_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15876_ _12905_ _12907_ VGND VGND VPWR VPWR _12908_ sky130_fd_sc_hd__xor2_1
XFILLER_64_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_237_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_237_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17615_ _04851_ _04852_ _04850_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__a21bo_1
X_14827_ _11941_ _11949_ VGND VGND VPWR VPWR _11952_ sky130_fd_sc_hd__xor2_1
XFILLER_92_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18595_ _05722_ _05723_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__or2_1
XFILLER_92_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17546_ systolic_inst.A_outs\[10\]\[6\] _11275_ _04771_ _04774_ _04796_ VGND VGND
+ VPWR VPWR _04797_ sky130_fd_sc_hd__o311a_1
X_14758_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.A_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\]
+ systolic_inst.A_outs\[14\]\[1\] VGND VGND VPWR VPWR _11887_ sky130_fd_sc_hd__and4_1
XFILLER_205_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13709_ B_in\[16\] deser_B.word_buffer\[16\] net84 VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__mux2_1
XFILLER_32_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17477_ _04728_ _04729_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14689_ _11799_ _11800_ _11822_ _11842_ VGND VGND VPWR VPWR _11843_ sky130_fd_sc_hd__a211o_1
XFILLER_225_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19216_ _06278_ _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__nor2_1
X_16428_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[12\]\[10\]
+ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__nor2_1
XFILLER_177_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19147_ systolic_inst.A_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[5\] VGND VGND VPWR
+ VPWR _06213_ sky130_fd_sc_hd__nand2_1
XFILLER_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16359_ _03658_ _03659_ _03722_ _03720_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_184_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_184_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19078_ systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[5\]
+ systolic_inst.B_outs\[7\]\[0\] VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__a22oi_1
XFILLER_173_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18029_ _05150_ _05219_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__nor2_1
XFILLER_105_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21040_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[8\] _07912_ net117
+ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__mux2_1
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22991_ _09634_ _09636_ _09666_ VGND VGND VPWR VPWR _09668_ sky130_fd_sc_hd__nand3_1
XFILLER_210_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24730_ net112 ser_C.shift_reg\[193\] VGND VGND VPWR VPWR _10835_ sky130_fd_sc_hd__and2_1
X_21942_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[3\]\[10\]
+ _08725_ _08727_ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__a31o_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21873_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[3\]\[0\]
+ _08671_ _08672_ VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__and4_1
X_24661_ C_out\[157\] net104 _10643_ ser_C.shift_reg\[157\] _10800_ VGND VGND VPWR
+ VPWR _02407_ sky130_fd_sc_hd__a221o_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26400_ clknet_leaf_31_clk _00207_ net133 VGND VGND VPWR VPWR A_in\[68\] sky130_fd_sc_hd__dfrtp_1
X_20824_ _07716_ _07720_ _07721_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__a21oi_1
X_23612_ _10231_ _10232_ VGND VGND VPWR VPWR _10233_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27380_ clknet_leaf_333_clk _01178_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24592_ net114 ser_C.shift_reg\[124\] VGND VGND VPWR VPWR _10766_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_173_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26331_ clknet_leaf_30_A_in_serial_clk _00138_ net132 VGND VGND VPWR VPWR deser_A.serial_toggle
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20755_ systolic_inst.acc_wires\[5\]\[16\] systolic_inst.acc_wires\[5\]\[17\] systolic_inst.acc_wires\[5\]\[18\]
+ systolic_inst.acc_wires\[5\]\[19\] systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__o41a_1
X_23543_ _10164_ _10165_ VGND VGND VPWR VPWR _10166_ sky130_fd_sc_hd__or2_1
XFILLER_196_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29050_ clknet_leaf_103_clk _02848_ net151 VGND VGND VPWR VPWR C_out\[22\] sky130_fd_sc_hd__dfrtp_1
X_23474_ _10054_ _10056_ _10097_ _10098_ VGND VGND VPWR VPWR _10099_ sky130_fd_sc_hd__o211a_1
X_26262_ clknet_leaf_5_A_in_serial_clk _00070_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_20686_ _07598_ _07604_ VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__nand2_1
X_28001_ clknet_leaf_153_clk _01799_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22425_ _09096_ _09135_ _09134_ VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__a21bo_1
X_25213_ C_out\[433\] net101 net73 ser_C.shift_reg\[433\] _11076_ VGND VGND VPWR VPWR
+ _02683_ sky130_fd_sc_hd__a221o_1
XFILLER_210_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26193_ _11301_ _11256_ net82 ser_C.bit_idx\[8\] VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_137_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22356_ systolic_inst.A_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[5\] systolic_inst.B_outs\[2\]\[6\]
+ systolic_inst.B_outs\[2\]\[7\] VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25144_ net110 ser_C.shift_reg\[400\] VGND VGND VPWR VPWR _11042_ sky130_fd_sc_hd__and2_1
XFILLER_87_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21307_ net63 _08162_ _08163_ systolic_inst.acc_wires\[4\]\[8\] net108 VGND VGND
+ VPWR VPWR _01690_ sky130_fd_sc_hd__a32o_1
XFILLER_156_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25075_ C_out\[364\] net97 net77 ser_C.shift_reg\[364\] _11007_ VGND VGND VPWR VPWR
+ _02614_ sky130_fd_sc_hd__a221o_1
X_22287_ systolic_inst.A_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[6\]
+ systolic_inst.B_outs\[2\]\[7\] VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__and4b_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24026_ _10530_ systolic_inst.B_shift\[4\]\[0\] net72 VGND VGND VPWR VPWR _02042_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28903_ clknet_leaf_272_clk _02701_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[451\]
+ sky130_fd_sc_hd__dfrtp_1
X_21238_ _08079_ _08081_ _08103_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__and3_1
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28834_ clknet_leaf_237_clk _02632_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_238_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21169_ _08036_ _08037_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__nand2_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28765_ clknet_leaf_214_clk _02563_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13991_ deser_B.shift_reg\[25\] deser_B.shift_reg\[26\] net125 VGND VGND VPWR VPWR
+ _00817_ sky130_fd_sc_hd__mux2_1
X_25977_ systolic_inst.acc_wires\[14\]\[5\] ser_C.parallel_data\[453\] net24 VGND
+ VGND VPWR VPWR _03279_ sky130_fd_sc_hd__mux2_1
XFILLER_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27716_ clknet_leaf_189_clk _01514_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_15730_ _12715_ _12759_ _12758_ VGND VGND VPWR VPWR _12782_ sky130_fd_sc_hd__o21a_1
XFILLER_105_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24928_ net111 ser_C.shift_reg\[292\] VGND VGND VPWR VPWR _10934_ sky130_fd_sc_hd__and2_1
X_28696_ clknet_leaf_193_clk _02494_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15661_ _12713_ _12714_ VGND VGND VPWR VPWR _12715_ sky130_fd_sc_hd__nand2_1
X_27647_ clknet_leaf_314_clk _01445_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24859_ C_out\[256\] net103 net75 ser_C.shift_reg\[256\] _10899_ VGND VGND VPWR VPWR
+ _02506_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_83_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17400_ _04647_ _04655_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__xnor2_1
X_14612_ _11774_ _11775_ _11776_ VGND VGND VPWR VPWR _11778_ sky130_fd_sc_hd__a21oi_1
X_18380_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[28\]
+ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_232_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ systolic_inst.B_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[7\]
+ VGND VGND VPWR VPWR _12648_ sky130_fd_sc_hd__and3_1
X_27578_ clknet_leaf_219_clk _01376_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_232_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29317_ clknet_leaf_297_clk _03115_ net139 VGND VGND VPWR VPWR C_out\[289\] sky130_fd_sc_hd__dfrtp_1
X_17331_ _04548_ _04550_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__and2b_1
X_14543_ _11715_ _11716_ _11717_ VGND VGND VPWR VPWR _11719_ sky130_fd_sc_hd__and3_1
XFILLER_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26529_ clknet_leaf_5_A_in_serial_clk _00332_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_222_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29248_ clknet_leaf_185_clk _03046_ net146 VGND VGND VPWR VPWR C_out\[220\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17262_ _04511_ _04520_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__xor2_1
X_14474_ _11626_ _11654_ VGND VGND VPWR VPWR _11655_ sky130_fd_sc_hd__xnor2_1
X_19001_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[30\]
+ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__nand2_1
XFILLER_128_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16213_ _03560_ _03595_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__xor2_1
X_13425_ deser_A.bit_idx\[1\] deser_A.bit_idx\[2\] _11308_ VGND VGND VPWR VPWR _11312_
+ sky130_fd_sc_hd__and3_1
XFILLER_155_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29179_ clknet_leaf_136_clk _02977_ net142 VGND VGND VPWR VPWR C_out\[151\] sky130_fd_sc_hd__dfrtp_1
X_17193_ systolic_inst.B_outs\[9\]\[7\] systolic_inst.B_outs\[5\]\[7\] net116 VGND
+ VGND VPWR VPWR _01281_ sky130_fd_sc_hd__mux2_1
Xclkload107 clknet_leaf_281_clk VGND VGND VPWR VPWR clkload107/Y sky130_fd_sc_hd__bufinv_16
Xclkload118 clknet_leaf_278_clk VGND VGND VPWR VPWR clkload118/Y sky130_fd_sc_hd__bufinv_16
XFILLER_154_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload129 clknet_leaf_264_clk VGND VGND VPWR VPWR clkload129/X sky130_fd_sc_hd__clkbuf_8
X_16144_ systolic_inst.A_outs\[12\]\[2\] systolic_inst.B_outs\[12\]\[6\] _11260_ systolic_inst.A_outs\[12\]\[1\]
+ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13356_ A_in\[65\] deser_A.word_buffer\[65\] net96 VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__mux2_1
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16075_ _13068_ _13070_ VGND VGND VPWR VPWR _13071_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_226_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13287_ deser_A.word_buffer\[125\] deser_A.serial_word\[125\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_226_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19903_ _06861_ _06863_ _06862_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__o21ba_1
X_15026_ _12109_ _12144_ systolic_inst.A_outs\[14\]\[7\] VGND VGND VPWR VPWR _12145_
+ sky130_fd_sc_hd__and3b_1
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19834_ _06830_ _06833_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_239_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_239_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19765_ _06729_ _06764_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__xor2_1
X_16977_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[11\]\[0\]
+ _04285_ _04286_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__a22o_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 rst_n VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_12
XFILLER_65_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_177_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15928_ _12949_ _12951_ VGND VGND VPWR VPWR _12952_ sky130_fd_sc_hd__xnor2_1
X_18716_ _05807_ _05809_ _05808_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_177_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19696_ _06693_ _06698_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__xor2_1
XFILLER_237_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18647_ _05772_ _05773_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__nor2_1
X_15859_ _12880_ _12887_ _12888_ VGND VGND VPWR VPWR _12893_ sky130_fd_sc_hd__o21ba_1
XFILLER_40_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18578_ systolic_inst.A_outs\[8\]\[1\] _11259_ systolic_inst.B_outs\[8\]\[6\] systolic_inst.A_outs\[8\]\[2\]
+ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_224_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17529_ _04779_ _04780_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__nand2_1
XFILLER_166_1392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20540_ _07472_ _07471_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__nand2b_1
XFILLER_32_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20471_ _07369_ _07371_ _07370_ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__o21ba_1
XFILLER_192_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22210_ systolic_inst.B_outs\[2\]\[3\] systolic_inst.A_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\]
+ systolic_inst.A_outs\[2\]\[4\] VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__and4_1
X_23190_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[18\]
+ VGND VGND VPWR VPWR _09845_ sky130_fd_sc_hd__nand2_1
XFILLER_195_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_2_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_2_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22141_ net109 _08888_ _08889_ VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__or3_1
XFILLER_134_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22072_ _08829_ _08835_ _08839_ _08840_ _08841_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__o311ai_4
XFILLER_126_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25900_ systolic_inst.acc_wires\[11\]\[24\] C_out\[376\] net41 VGND VGND VPWR VPWR
+ _03202_ sky130_fd_sc_hd__mux2_1
X_21023_ _07887_ _07895_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_162_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26880_ clknet_leaf_12_A_in_serial_clk _00678_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25831_ systolic_inst.acc_wires\[9\]\[19\] C_out\[307\] net15 VGND VGND VPWR VPWR
+ _03133_ sky130_fd_sc_hd__mux2_1
XFILLER_214_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28550_ clknet_leaf_173_clk _02348_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_132_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25762_ systolic_inst.acc_wires\[7\]\[14\] C_out\[238\] net43 VGND VGND VPWR VPWR
+ _03064_ sky130_fd_sc_hd__mux2_1
X_22974_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[11\] _09651_ net122
+ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__mux2_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27501_ clknet_leaf_295_clk _01299_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_228_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24713_ C_out\[183\] net99 net79 ser_C.shift_reg\[183\] _10826_ VGND VGND VPWR VPWR
+ _02433_ sky130_fd_sc_hd__a221o_1
X_28481_ clknet_leaf_109_clk _02279_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_21925_ _08715_ _08716_ VGND VGND VPWR VPWR _08717_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25693_ systolic_inst.acc_wires\[5\]\[9\] C_out\[169\] net31 VGND VGND VPWR VPWR
+ _02995_ sky130_fd_sc_hd__mux2_1
XFILLER_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27432_ clknet_leaf_235_clk _01230_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24644_ net7 ser_C.shift_reg\[150\] VGND VGND VPWR VPWR _10792_ sky130_fd_sc_hd__and2_1
X_21856_ _08635_ _08658_ _08637_ _08612_ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_218_Right_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20807_ _07706_ _07707_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__nand2_1
XFILLER_180_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27363_ clknet_leaf_341_clk _01161_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24575_ C_out\[114\] net100 net80 ser_C.shift_reg\[114\] _10757_ VGND VGND VPWR VPWR
+ _02364_ sky130_fd_sc_hd__a221o_1
X_21787_ _08589_ _08590_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29102_ clknet_leaf_161_clk _02900_ net150 VGND VGND VPWR VPWR C_out\[74\] sky130_fd_sc_hd__dfrtp_1
X_26314_ clknet_leaf_28_A_in_serial_clk _00122_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23526_ _10144_ _10147_ VGND VGND VPWR VPWR _10149_ sky130_fd_sc_hd__xor2_1
XFILLER_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20738_ net106 systolic_inst.acc_wires\[5\]\[17\] net68 _07649_ VGND VGND VPWR VPWR
+ _01635_ sky130_fd_sc_hd__a22o_1
X_27294_ clknet_leaf_292_clk _01092_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29033_ clknet_leaf_126_clk _02831_ net144 VGND VGND VPWR VPWR C_out\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26245_ clknet_leaf_18_A_in_serial_clk _00053_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_23457_ _10078_ _10081_ VGND VGND VPWR VPWR _10082_ sky130_fd_sc_hd__xnor2_1
X_20669_ net64 _07589_ _07590_ systolic_inst.acc_wires\[5\]\[7\] net109 VGND VGND
+ VPWR VPWR _01625_ sky130_fd_sc_hd__a32o_1
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13210_ deser_A.word_buffer\[48\] deser_A.serial_word\[48\] net127 VGND VGND VPWR
+ VPWR _00058_ sky130_fd_sc_hd__mux2_1
X_22408_ _09146_ _09147_ VGND VGND VPWR VPWR _09149_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26176_ _11302_ _11245_ _11246_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__nor3_1
X_14190_ _11365_ _11367_ _11366_ VGND VGND VPWR VPWR _11379_ sky130_fd_sc_hd__a21bo_1
X_23388_ _10013_ _10014_ VGND VGND VPWR VPWR _10015_ sky130_fd_sc_hd__nand2_1
XFILLER_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13141_ systolic_inst.cycle_cnt\[11\] systolic_inst.cycle_cnt\[10\] systolic_inst.cycle_cnt\[9\]
+ systolic_inst.cycle_cnt\[8\] VGND VGND VPWR VPWR _11294_ sky130_fd_sc_hd__or4_1
XFILLER_137_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25127_ C_out\[390\] net101 net73 ser_C.shift_reg\[390\] _11033_ VGND VGND VPWR VPWR
+ _02640_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22339_ _09022_ _09080_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__or2_1
XFILLER_124_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25058_ net112 ser_C.shift_reg\[357\] VGND VGND VPWR VPWR _10999_ sky130_fd_sc_hd__and2_1
XFILLER_140_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16900_ _04215_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__nor2_1
X_24009_ systolic_inst.B_shift\[7\]\[0\] net70 net83 systolic_inst.B_shift\[11\]\[0\]
+ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__a22o_1
XFILLER_78_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_221_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17880_ _05045_ _05048_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_221_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16831_ _04149_ _04148_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__nand2b_1
XFILLER_66_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28817_ clknet_leaf_241_clk _02615_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[365\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19550_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[22\]
+ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__nand2_1
XFILLER_47_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16762_ _04082_ _04053_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__nand2b_1
X_28748_ clknet_leaf_222_clk _02546_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[296\]
+ sky130_fd_sc_hd__dfrtp_1
X_13974_ deser_B.shift_reg\[8\] deser_B.shift_reg\[9\] net125 VGND VGND VPWR VPWR
+ _00800_ sky130_fd_sc_hd__mux2_1
XFILLER_93_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_234_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18501_ _05603_ _05631_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__xor2_1
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15713_ _12732_ _12735_ _12765_ VGND VGND VPWR VPWR _12766_ sky130_fd_sc_hd__nor3_1
XFILLER_189_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19481_ _06497_ _06500_ _06509_ _06525_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__a211o_1
XFILLER_59_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_100_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28679_ clknet_leaf_196_clk _02477_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[227\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16693_ _03985_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18432_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[2\] _05565_ VGND
+ VGND VPWR VPWR _05567_ sky130_fd_sc_hd__a21o_1
X_15644_ _12657_ _12659_ _12697_ VGND VGND VPWR VPWR _12699_ sky130_fd_sc_hd__nand3_1
XFILLER_59_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18363_ _05518_ _05520_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_29_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15575_ _12629_ _12630_ VGND VGND VPWR VPWR _12632_ sky130_fd_sc_hd__xor2_1
XFILLER_226_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17314_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[5\] VGND VGND
+ VPWR VPWR _04572_ sky130_fd_sc_hd__nand2_1
XFILLER_42_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14526_ net105 systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] _11703_
+ _11704_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__a22o_1
XFILLER_186_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18294_ _05462_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__or2_1
XFILLER_226_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17245_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[2\] _04487_ _04474_
+ systolic_inst.B_outs\[10\]\[4\] VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__a32o_1
XFILLER_128_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14457_ _11588_ _11638_ VGND VGND VPWR VPWR _11639_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_228_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13408_ A_in\[117\] deser_A.word_buffer\[117\] _00003_ VGND VGND VPWR VPWR _00256_
+ sky130_fd_sc_hd__mux2_1
X_17176_ _04451_ _04455_ _04456_ net60 VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__a31o_1
X_14388_ _11569_ _11570_ VGND VGND VPWR VPWR _11572_ sky130_fd_sc_hd__xor2_1
XFILLER_196_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16127_ net108 _03510_ _03511_ _03512_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__o31ai_1
XFILLER_192_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13339_ A_in\[48\] deser_A.word_buffer\[48\] net93 VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__mux2_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16058_ net115 _13053_ _13054_ _13025_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__a31o_1
XFILLER_233_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15009_ _12126_ _12127_ VGND VGND VPWR VPWR _12129_ sky130_fd_sc_hd__xnor2_1
XFILLER_237_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19817_ _06816_ _06815_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__and2b_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19748_ _06748_ _06749_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__nor2_1
XFILLER_84_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19679_ net120 _06681_ _06682_ _06683_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__a31o_1
XFILLER_129_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21710_ _08515_ _08516_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__or2_1
XFILLER_240_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22690_ _11258_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[0\] _09378_
+ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__a21o_1
XFILLER_198_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21641_ _08448_ _08449_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__nor2_1
XFILLER_75_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24360_ net7 ser_C.shift_reg\[8\] VGND VGND VPWR VPWR _10650_ sky130_fd_sc_hd__and2_1
X_21572_ systolic_inst.B_outs\[3\]\[3\] systolic_inst.A_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\]
+ systolic_inst.A_outs\[3\]\[2\] VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__a22oi_1
XFILLER_123_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_10 systolic_inst.B_outs\[3\]\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_32 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23311_ _09924_ _09926_ _09938_ _09919_ VGND VGND VPWR VPWR _09941_ sky130_fd_sc_hd__or4b_2
X_20523_ _07417_ _07419_ _07454_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__a21o_1
X_24291_ systolic_inst.A_shift\[12\]\[1\] A_in\[49\] net59 VGND VGND VPWR VPWR _10619_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26030_ systolic_inst.acc_wires\[15\]\[26\] ser_C.parallel_data\[506\] net37 VGND
+ VGND VPWR VPWR _03332_ sky130_fd_sc_hd__mux2_1
X_23242_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[26\]
+ VGND VGND VPWR VPWR _09889_ sky130_fd_sc_hd__nand2_1
XFILLER_193_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20454_ _07387_ _07388_ _07389_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__and3_1
XFILLER_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23173_ _09821_ _09826_ _09830_ VGND VGND VPWR VPWR _09831_ sky130_fd_sc_hd__a21oi_1
XFILLER_175_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20385_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[7\]
+ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__o21ai_2
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22124_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.A_outs\[2\]\[1\] systolic_inst.B_outs\[2\]\[3\]
+ systolic_inst.B_outs\[2\]\[4\] VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_164_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27981_ clknet_leaf_118_clk _01779_ net152 VGND VGND VPWR VPWR systolic_inst.A_outs\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_82_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22055_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[28\]
+ VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26932_ clknet_leaf_16_A_in_serial_clk _00730_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21006_ _07874_ _07878_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__nand2_1
X_29651_ clknet_leaf_5_B_in_serial_clk _03446_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26863_ clknet_leaf_89_clk deser_B.serial_toggle_sync1 net5 VGND VGND VPWR VPWR deser_B.serial_toggle_sync2
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_134_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28602_ clknet_leaf_137_clk _02400_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[150\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25814_ systolic_inst.acc_wires\[9\]\[2\] C_out\[290\] net14 VGND VGND VPWR VPWR
+ _03116_ sky130_fd_sc_hd__mux2_1
XFILLER_169_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29582_ clknet_leaf_19_B_in_serial_clk _03377_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_26794_ clknet_leaf_85_clk _00596_ net153 VGND VGND VPWR VPWR B_in\[66\] sky130_fd_sc_hd__dfrtp_1
XFILLER_235_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28533_ clknet_leaf_161_clk _02331_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[81\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap23 net24 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_6
XFILLER_44_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25745_ systolic_inst.acc_wires\[6\]\[29\] C_out\[221\] net43 VGND VGND VPWR VPWR
+ _03047_ sky130_fd_sc_hd__mux2_1
Xmax_cap34 net35 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_8
X_22957_ _09632_ _09633_ VGND VGND VPWR VPWR _09635_ sky130_fd_sc_hd__xnor2_1
Xmax_cap45 net46 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_6
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap56 _00001_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_104_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap67 _11712_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_104_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28464_ clknet_leaf_121_clk _02262_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_21908_ _08700_ _08702_ _08694_ _08698_ VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__a211o_1
Xmax_cap78 net79 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_12
XFILLER_231_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13690_ deser_B.word_buffer\[126\] deser_B.serial_word\[126\] net123 VGND VGND VPWR
+ VPWR _00527_ sky130_fd_sc_hd__mux2_1
X_25676_ systolic_inst.acc_wires\[4\]\[24\] C_out\[152\] net32 VGND VGND VPWR VPWR
+ _02978_ sky130_fd_sc_hd__mux2_1
XFILLER_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap89 _00005_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_8
X_22888_ _09567_ _09566_ VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_65_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27415_ clknet_leaf_214_clk _01213_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_24627_ C_out\[140\] net103 net76 ser_C.shift_reg\[140\] _10783_ VGND VGND VPWR VPWR
+ _02390_ sky130_fd_sc_hd__a221o_1
XFILLER_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21839_ systolic_inst.B_outs\[3\]\[5\] systolic_inst.B_outs\[3\]\[6\] systolic_inst.A_outs\[3\]\[7\]
+ _08641_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__a31o_1
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28395_ clknet_leaf_33_clk _02193_ VGND VGND VPWR VPWR systolic_inst.A_shift\[17\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ systolic_inst.A_outs\[13\]\[4\] systolic_inst.A_outs\[12\]\[4\] net115 VGND
+ VGND VPWR VPWR _01078_ sky130_fd_sc_hd__mux2_1
X_27346_ clknet_leaf_342_clk _01144_ net131 VGND VGND VPWR VPWR systolic_inst.A_outs\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_24558_ net113 ser_C.shift_reg\[107\] VGND VGND VPWR VPWR _10749_ sky130_fd_sc_hd__and2_1
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14311_ _11451_ _11458_ _11457_ VGND VGND VPWR VPWR _11497_ sky130_fd_sc_hd__a21boi_1
X_23509_ _10130_ _10131_ _10113_ VGND VGND VPWR VPWR _10133_ sky130_fd_sc_hd__o21a_1
XFILLER_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15291_ _12374_ _12379_ _12381_ net61 VGND VGND VPWR VPWR _12384_ sky130_fd_sc_hd__a31o_1
X_27277_ clknet_leaf_325_clk _01075_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_78_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24489_ C_out\[71\] _11302_ net81 ser_C.shift_reg\[71\] _10714_ VGND VGND VPWR VPWR
+ _02321_ sky130_fd_sc_hd__a221o_1
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29016_ clknet_leaf_93_clk _02814_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17030_ net60 _04333_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__nor2_1
XFILLER_183_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26228_ clknet_leaf_7_A_in_serial_clk _00036_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14242_ _11397_ _11399_ _11428_ _11429_ VGND VGND VPWR VPWR _11430_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_20_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26159_ deser_B.serial_word\[114\] deser_B.shift_reg\[114\] net56 VGND VGND VPWR
+ VPWR _03461_ sky130_fd_sc_hd__mux2_1
X_14173_ _11347_ _11362_ VGND VGND VPWR VPWR _11363_ sky130_fd_sc_hd__nor2_1
XFILLER_124_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_223_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13124_ _11279_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__clkinv_16
XFILLER_125_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18981_ net108 systolic_inst.acc_wires\[8\]\[26\] net66 _06075_ VGND VGND VPWR VPWR
+ _01452_ sky130_fd_sc_hd__a22o_1
XFILLER_79_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17932_ systolic_inst.A_outs\[9\]\[1\] systolic_inst.B_outs\[9\]\[6\] _05125_ VGND
+ VGND VPWR VPWR _05126_ sky130_fd_sc_hd__and3_1
XFILLER_117_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17863_ systolic_inst.A_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[5\] VGND VGND VPWR
+ VPWR _05059_ sky130_fd_sc_hd__nand2_1
XFILLER_87_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19602_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[30\]
+ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16814_ systolic_inst.A_outs\[11\]\[6\] _04132_ _04131_ VGND VGND VPWR VPWR _04133_
+ sky130_fd_sc_hd__a21bo_1
X_17794_ systolic_inst.B_outs\[8\]\[1\] systolic_inst.B_outs\[4\]\[1\] net121 VGND
+ VGND VPWR VPWR _01339_ sky130_fd_sc_hd__mux2_1
XFILLER_238_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19533_ _06569_ _06570_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__xnor2_1
X_16745_ _04064_ _04065_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__xnor2_1
X_13957_ deser_A.serial_word\[118\] deser_A.shift_reg\[118\] _00002_ VGND VGND VPWR
+ VPWR _00783_ sky130_fd_sc_hd__mux2_1
XFILLER_62_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19464_ net60 _06511_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__nor2_1
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16676_ systolic_inst.A_outs\[11\]\[1\] systolic_inst.B_outs\[11\]\[5\] systolic_inst.B_outs\[11\]\[6\]
+ systolic_inst.A_outs\[11\]\[0\] VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__a22oi_1
XFILLER_222_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13888_ deser_A.serial_word\[49\] deser_A.shift_reg\[49\] net58 VGND VGND VPWR VPWR
+ _00714_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18415_ systolic_inst.B_outs\[7\]\[4\] systolic_inst.B_outs\[3\]\[4\] net119 VGND
+ VGND VPWR VPWR _01406_ sky130_fd_sc_hd__mux2_1
X_15627_ _12577_ _12681_ VGND VGND VPWR VPWR _12682_ sky130_fd_sc_hd__or2_1
X_19395_ _06237_ _06372_ _06444_ _06442_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__a31o_1
XFILLER_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18346_ net66 _05507_ _05508_ systolic_inst.acc_wires\[9\]\[22\] net106 VGND VGND
+ VPWR VPWR _01384_ sky130_fd_sc_hd__a32o_1
XFILLER_124_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15558_ _12613_ _12614_ VGND VGND VPWR VPWR _12615_ sky130_fd_sc_hd__or2_1
XFILLER_226_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_212_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14509_ _11686_ _11687_ VGND VGND VPWR VPWR _11689_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_13_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18277_ net107 systolic_inst.acc_wires\[9\]\[12\] net66 _05449_ VGND VGND VPWR VPWR
+ _01374_ sky130_fd_sc_hd__a22o_1
X_15489_ systolic_inst.B_outs\[13\]\[3\] systolic_inst.A_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\]
+ systolic_inst.A_outs\[13\]\[4\] VGND VGND VPWR VPWR _12548_ sky130_fd_sc_hd__and4_1
X_17228_ _04486_ _04488_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17159_ _04440_ _04443_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__xor2_1
X_20170_ _07131_ _07135_ _07138_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__a21o_1
XFILLER_104_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23860_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[26\]
+ VGND VGND VPWR VPWR _10451_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_198_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22811_ _09488_ _09492_ VGND VGND VPWR VPWR _09493_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23791_ net63 _10392_ _10393_ systolic_inst.acc_wires\[0\]\[14\] _11258_ VGND VGND
+ VPWR VPWR _01944_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_0_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25530_ systolic_inst.acc_wires\[0\]\[6\] C_out\[6\] net33 VGND VGND VPWR VPWR _02832_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22742_ _09422_ _09425_ VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_157_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25461_ systolic_inst.cycle_cnt\[8\] _11306_ _11199_ systolic_inst.cycle_cnt\[9\]
+ VGND VGND VPWR VPWR _11205_ sky130_fd_sc_hd__a31o_1
XFILLER_197_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22673_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.A_outs\[0\]\[0\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27200_ clknet_leaf_262_clk _00998_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_240_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24412_ net114 ser_C.shift_reg\[34\] VGND VGND VPWR VPWR _10676_ sky130_fd_sc_hd__and2_1
XFILLER_209_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21624_ _08403_ _08432_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__xnor2_1
X_28180_ clknet_leaf_64_clk _01978_ VGND VGND VPWR VPWR systolic_inst.A_shift\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25392_ _11165_ systolic_inst.A_shift\[2\]\[3\] net71 VGND VGND VPWR VPWR _02773_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27131_ clknet_leaf_14_clk _00929_ VGND VGND VPWR VPWR systolic_inst.A_shift\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_205_Left_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24343_ systolic_inst.A_shift\[8\]\[6\] net70 net83 systolic_inst.A_shift\[9\]\[6\]
+ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__a22o_1
X_21555_ _08365_ _08366_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__and2_1
XFILLER_178_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27062_ clknet_leaf_6_B_in_serial_clk _00860_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[68\]
+ sky130_fd_sc_hd__dfrtp_1
X_20506_ _07436_ _07439_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__xor2_1
X_21486_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[1\] _08299_
+ _08301_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__a22o_1
X_24274_ _10610_ systolic_inst.B_shift\[23\]\[0\] net71 VGND VGND VPWR VPWR _02210_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26013_ systolic_inst.acc_wires\[15\]\[9\] ser_C.parallel_data\[489\] net39 VGND
+ VGND VPWR VPWR _03315_ sky130_fd_sc_hd__mux2_1
XFILLER_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23225_ _09866_ _09870_ _09873_ VGND VGND VPWR VPWR _09875_ sky130_fd_sc_hd__a21o_1
X_20437_ _07369_ _07372_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23156_ _09810_ _09814_ VGND VGND VPWR VPWR _09816_ sky130_fd_sc_hd__nand2b_1
X_20368_ _07270_ _07305_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__xnor2_1
Xclkload290 clknet_leaf_194_clk VGND VGND VPWR VPWR clkload290/Y sky130_fd_sc_hd__clkinv_2
XFILLER_136_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22107_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[2\] _08856_ VGND
+ VGND VPWR VPWR _08858_ sky130_fd_sc_hd__a21o_1
X_23087_ _09750_ _09751_ _09749_ VGND VGND VPWR VPWR _09757_ sky130_fd_sc_hd__a21bo_1
X_27964_ clknet_leaf_168_clk _01762_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_216_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20299_ _07236_ _07237_ _07238_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__or3_1
XFILLER_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22038_ net65 _08812_ _08813_ systolic_inst.acc_wires\[3\]\[25\] net106 VGND VGND
+ VPWR VPWR _01771_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_214_Left_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26915_ clknet_leaf_10_A_in_serial_clk _00713_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27895_ clknet_leaf_39_clk _01693_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29634_ clknet_leaf_26_B_in_serial_clk _03429_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_26846_ clknet_leaf_68_clk _00648_ net135 VGND VGND VPWR VPWR B_in\[118\] sky130_fd_sc_hd__dfrtp_1
X_14860_ _11938_ _11940_ _11982_ VGND VGND VPWR VPWR _11984_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_106_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ B_in\[118\] deser_B.word_buffer\[118\] net87 VGND VGND VPWR VPWR _00648_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29565_ clknet_leaf_16_B_in_serial_clk _03360_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_26777_ clknet_leaf_78_clk _00579_ net143 VGND VGND VPWR VPWR B_in\[49\] sky130_fd_sc_hd__dfrtp_1
XFILLER_112_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14791_ _11913_ _11916_ VGND VGND VPWR VPWR _11917_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23989_ systolic_inst.B_shift\[12\]\[6\] B_in\[70\] _00008_ VGND VGND VPWR VPWR _10520_
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28516_ clknet_leaf_155_clk _02314_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16530_ _03864_ _03873_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_216_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13742_ B_in\[49\] deser_B.word_buffer\[49\] net86 VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__mux2_1
X_25728_ systolic_inst.acc_wires\[6\]\[12\] C_out\[204\] net45 VGND VGND VPWR VPWR
+ _03030_ sky130_fd_sc_hd__mux2_1
X_29496_ clknet_leaf_269_clk _03294_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16461_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[12\]\[14\]
+ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__or2_1
XFILLER_44_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28447_ clknet_leaf_35_clk _02245_ VGND VGND VPWR VPWR systolic_inst.A_shift\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_232_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13673_ deser_B.word_buffer\[109\] deser_B.serial_word\[109\] net123 VGND VGND VPWR
+ VPWR _00510_ sky130_fd_sc_hd__mux2_1
XFILLER_31_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25659_ systolic_inst.acc_wires\[4\]\[7\] C_out\[135\] net29 VGND VGND VPWR VPWR
+ _02961_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_191_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_191_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_189_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18200_ net66 _05382_ _05383_ systolic_inst.acc_wires\[9\]\[1\] net107 VGND VGND
+ VPWR VPWR _01363_ sky130_fd_sc_hd__a32o_1
XFILLER_223_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15412_ _12453_ _12471_ _12472_ VGND VGND VPWR VPWR _12474_ sky130_fd_sc_hd__or3_1
XFILLER_227_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_223_Left_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19180_ _06243_ _06244_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__nor2_1
X_16392_ _03762_ _03764_ _03757_ _03760_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__a211o_1
X_28378_ clknet_leaf_32_clk _02176_ VGND VGND VPWR VPWR systolic_inst.A_shift\[19\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18131_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[12\] _05319_ net116
+ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__mux2_1
X_15343_ net107 systolic_inst.acc_wires\[14\]\[29\] _11712_ _12427_ VGND VGND VPWR
+ VPWR _01071_ sky130_fd_sc_hd__a22o_1
X_27329_ clknet_leaf_330_clk _01127_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_12_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18062_ _05250_ _05251_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__nand2_1
XFILLER_200_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15274_ net107 systolic_inst.acc_wires\[14\]\[18\] _11712_ _12369_ VGND VGND VPWR
+ VPWR _01060_ sky130_fd_sc_hd__a22o_1
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17013_ net69 _04317_ _04319_ systolic_inst.acc_wires\[11\]\[6\] net105 VGND VGND
+ VPWR VPWR _01240_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_97_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14225_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[6\] _11411_ _11412_
+ VGND VGND VPWR VPWR _11413_ sky130_fd_sc_hd__nand4_2
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14156_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[1\] systolic_inst.A_outs\[15\]\[2\]
+ systolic_inst.B_outs\[15\]\[2\] VGND VGND VPWR VPWR _11347_ sky130_fd_sc_hd__nand4_2
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_242_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ systolic_inst.B_outs\[9\]\[7\] VGND VGND VPWR VPWR _11263_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_232_Left_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14087_ deser_B.shift_reg\[121\] deser_B.shift_reg\[122\] deser_B.receiving VGND
+ VGND VPWR VPWR _00913_ sky130_fd_sc_hd__mux2_1
X_18964_ _06040_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nor2_1
XFILLER_234_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17915_ _05079_ _05082_ _05084_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18895_ _06000_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__and2_1
XFILLER_39_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17846_ _05041_ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__or2_1
XFILLER_66_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14989_ systolic_inst.B_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[7\]
+ VGND VGND VPWR VPWR _12109_ sky130_fd_sc_hd__and3_1
X_17777_ _04994_ _04995_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_193_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19516_ _06554_ _06555_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__nor2_1
X_16728_ _04017_ _04048_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_241_Left_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19447_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[7\]\[7\]
+ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16659_ _03963_ _03981_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_182_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_182_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_18_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19378_ _06411_ _06413_ _06436_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__a21oi_1
XFILLER_194_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18329_ _05469_ _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__nor2_1
XFILLER_202_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21340_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[4\]\[13\]
+ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__nand2_1
XFILLER_198_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21271_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[4\]\[3\]
+ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__or2_1
XFILLER_190_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_208_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_208_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23010_ systolic_inst.B_outs\[1\]\[6\] systolic_inst.A_outs\[1\]\[7\] VGND VGND VPWR
+ VPWR _09686_ sky130_fd_sc_hd__nand2_1
X_20222_ _07183_ _07182_ systolic_inst.acc_wires\[6\]\[31\] net106 VGND VGND VPWR
+ VPWR _01585_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20153_ net62 _07124_ _07125_ systolic_inst.acc_wires\[6\]\[20\] net106 VGND VGND
+ VPWR VPWR _01574_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_146_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20084_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[6\]\[11\]
+ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__or2_1
X_24961_ C_out\[307\] net103 net76 ser_C.shift_reg\[307\] _10950_ VGND VGND VPWR VPWR
+ _02557_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_142_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_B_in_serial_clk clknet_0_B_in_serial_clk VGND VGND VPWR VPWR clknet_2_0__leaf_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_5_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26700_ clknet_leaf_6_B_in_serial_clk _00503_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23912_ systolic_inst.B_shift\[22\]\[0\] B_in\[80\] _00008_ VGND VGND VPWR VPWR _10489_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27680_ clknet_leaf_200_clk _01478_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24892_ net110 ser_C.shift_reg\[274\] VGND VGND VPWR VPWR _10916_ sky130_fd_sc_hd__and2_1
XFILLER_214_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26631_ clknet_leaf_19_B_in_serial_clk _00434_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23843_ _10429_ _10433_ _10435_ VGND VGND VPWR VPWR _10437_ sky130_fd_sc_hd__a21oi_1
XFILLER_85_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29350_ clknet_leaf_295_clk _03148_ net138 VGND VGND VPWR VPWR C_out\[322\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26562_ clknet_leaf_27_A_in_serial_clk _00365_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23774_ _10375_ _10376_ _10377_ VGND VGND VPWR VPWR _10379_ sky130_fd_sc_hd__a21oi_1
XFILLER_214_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20986_ _07814_ _07818_ _07858_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__a21bo_1
X_28301_ clknet_leaf_66_clk _02099_ VGND VGND VPWR VPWR systolic_inst.B_shift\[27\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25513_ systolic_inst.cycle_cnt\[27\] systolic_inst.cycle_cnt\[26\] _11233_ _11279_
+ systolic_inst.cycle_cnt\[28\] VGND VGND VPWR VPWR _11238_ sky130_fd_sc_hd__a32o_1
XFILLER_225_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22725_ systolic_inst.A_outs\[1\]\[4\] _09409_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__nand2_1
X_29281_ clknet_leaf_184_clk _03079_ net146 VGND VGND VPWR VPWR C_out\[253\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_173_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_173_clk
+ sky130_fd_sc_hd__clkbuf_8
X_26493_ clknet_leaf_8_A_in_serial_clk _00296_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28232_ clknet_leaf_129_clk _02030_ VGND VGND VPWR VPWR systolic_inst.B_shift\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_241_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25444_ systolic_inst.cycle_cnt\[4\] _11191_ VGND VGND VPWR VPWR _11193_ sky130_fd_sc_hd__nand2_1
XFILLER_90_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22656_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[29\]
+ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__xor2_1
XFILLER_198_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28163_ clknet_leaf_107_clk _01961_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_21607_ _08413_ _08416_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__xnor2_1
X_25375_ systolic_inst.B_shift\[18\]\[3\] B_in\[51\] net59 VGND VGND VPWR VPWR _11157_
+ sky130_fd_sc_hd__mux2_1
X_22587_ net109 systolic_inst.acc_wires\[2\]\[17\] net65 _09306_ VGND VGND VPWR VPWR
+ _01827_ sky130_fd_sc_hd__a22o_1
XFILLER_166_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27114_ clknet_leaf_31_B_in_serial_clk _00912_ net134 VGND VGND VPWR VPWR deser_B.shift_reg\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_24326_ _10636_ systolic_inst.A_shift\[9\]\[2\] net70 VGND VGND VPWR VPWR _02236_
+ sky130_fd_sc_hd__mux2_1
X_28094_ clknet_leaf_112_clk _01892_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_21538_ _08349_ _08346_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__nand2b_1
XFILLER_139_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27045_ clknet_leaf_25_B_in_serial_clk _00843_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_177_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24257_ systolic_inst.A_shift\[16\]\[0\] net70 net83 systolic_inst.A_shift\[17\]\[0\]
+ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__a22o_1
X_21469_ systolic_inst.A_outs\[3\]\[5\] systolic_inst.A_outs\[2\]\[5\] net122 VGND
+ VGND VPWR VPWR _01719_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14010_ deser_B.shift_reg\[44\] deser_B.shift_reg\[45\] net125 VGND VGND VPWR VPWR
+ _00836_ sky130_fd_sc_hd__mux2_1
XFILLER_88_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23208_ net65 _09859_ _09860_ systolic_inst.acc_wires\[1\]\[20\] net109 VGND VGND
+ VPWR VPWR _01894_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_92_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24188_ systolic_inst.A_shift\[24\]\[3\] net70 _10505_ systolic_inst.A_shift\[25\]\[3\]
+ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__a22o_1
XFILLER_49_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23139_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[1\]\[11\]
+ VGND VGND VPWR VPWR _09801_ sky130_fd_sc_hd__or2_1
X_28996_ clknet_leaf_92_clk _02794_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15961_ systolic_inst.A_outs\[12\]\[2\] systolic_inst.A_shift\[24\]\[2\] net115 VGND
+ VGND VPWR VPWR _01140_ sky130_fd_sc_hd__mux2_1
XFILLER_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27947_ clknet_leaf_148_clk _01745_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17700_ systolic_inst.acc_wires\[10\]\[16\] systolic_inst.acc_wires\[10\]\[17\] systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__o21a_1
XFILLER_23_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14912_ _12029_ _12032_ VGND VGND VPWR VPWR _12034_ sky130_fd_sc_hd__xnor2_1
X_27878_ clknet_leaf_37_clk _01676_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_15892_ _12920_ VGND VGND VPWR VPWR _12921_ sky130_fd_sc_hd__inv_2
X_18680_ _05735_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__xnor2_4
XFILLER_97_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29617_ clknet_leaf_4_B_in_serial_clk _03412_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_14843_ _11936_ _11965_ VGND VGND VPWR VPWR _11967_ sky130_fd_sc_hd__nor2_1
X_17631_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[10\]\[9\]
+ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__xor2_1
X_26829_ clknet_leaf_86_clk _00631_ net153 VGND VGND VPWR VPWR B_in\[101\] sky130_fd_sc_hd__dfrtp_1
XFILLER_236_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17562_ _04810_ _04811_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14774_ _11899_ _11900_ VGND VGND VPWR VPWR _11901_ sky130_fd_sc_hd__or2_1
X_29548_ clknet_leaf_229_clk _03343_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19301_ _06308_ _06326_ _06325_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__o21a_1
X_16513_ _03867_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__xor2_1
X_13725_ B_in\[32\] deser_B.word_buffer\[32\] net85 VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__mux2_1
XFILLER_147_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17493_ systolic_inst.B_outs\[10\]\[5\] systolic_inst.A_outs\[10\]\[7\] VGND VGND
+ VPWR VPWR _04746_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_164_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_164_clk
+ sky130_fd_sc_hd__clkbuf_8
X_29479_ clknet_leaf_271_clk _03277_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[451\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19232_ _06295_ _06294_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__nand2b_1
X_16444_ _03780_ _03783_ _03808_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13656_ deser_B.word_buffer\[92\] deser_B.serial_word\[92\] net123 VGND VGND VPWR
+ VPWR _00493_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19163_ _06199_ _06227_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_45_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16375_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[12\]\[2\]
+ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__nand2_1
X_13587_ deser_B.word_buffer\[23\] deser_B.serial_word\[23\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__mux2_1
XFILLER_129_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18114_ _05269_ _05271_ _05301_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__nand3_1
X_15326_ net107 systolic_inst.acc_wires\[14\]\[26\] _11712_ _12413_ VGND VGND VPWR
+ VPWR _01068_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19094_ _06137_ _06160_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_41_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18045_ _05226_ _05234_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__or2_1
X_15257_ _12353_ _12354_ VGND VGND VPWR VPWR _12355_ sky130_fd_sc_hd__and2_1
XFILLER_172_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14208_ _11370_ _11396_ VGND VGND VPWR VPWR _11397_ sky130_fd_sc_hd__nand2_1
XFILLER_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15188_ _12286_ _12290_ _12293_ _12294_ VGND VGND VPWR VPWR _12296_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_182_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14139_ systolic_inst.B_outs\[14\]\[7\] systolic_inst.B_outs\[10\]\[7\] net120 VGND
+ VGND VPWR VPWR _00961_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_203_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19996_ _06989_ _06990_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__nor2_1
XFILLER_235_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18947_ _06046_ _06045_ systolic_inst.acc_wires\[8\]\[21\] net108 VGND VGND VPWR
+ VPWR _01447_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18878_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[8\]\[11\]
+ _05982_ _05985_ _05986_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__a221oi_2
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17829_ _05025_ _05026_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__and2b_1
XFILLER_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20840_ systolic_inst.B_outs\[3\]\[5\] systolic_inst.B_shift\[3\]\[5\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__mux2_1
XFILLER_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_155_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_155_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20771_ net68 _07676_ _07677_ systolic_inst.acc_wires\[5\]\[22\] net106 VGND VGND
+ VPWR VPWR _01640_ sky130_fd_sc_hd__a32o_1
XFILLER_120_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22510_ _09237_ _09238_ _09239_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__and3_1
XFILLER_223_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23490_ systolic_inst.A_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[6\] VGND VGND VPWR
+ VPWR _10114_ sky130_fd_sc_hd__nand2_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22441_ systolic_inst.A_outs\[2\]\[6\] _11265_ _09154_ _09157_ _09179_ VGND VGND
+ VPWR VPWR _09180_ sky130_fd_sc_hd__o311a_1
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25160_ net110 ser_C.shift_reg\[408\] VGND VGND VPWR VPWR _11050_ sky130_fd_sc_hd__and2_1
X_22372_ _09112_ _09113_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__nor2_1
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24111_ systolic_inst.B_shift\[1\]\[6\] _11332_ net83 systolic_inst.B_shift\[5\]\[6\]
+ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__a22o_1
XFILLER_159_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21323_ _08175_ _08176_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__nand2_1
XFILLER_11_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25091_ C_out\[372\] net98 net78 ser_C.shift_reg\[372\] _11015_ VGND VGND VPWR VPWR
+ _02622_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_148_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24042_ _10538_ systolic_inst.B_shift\[0\]\[0\] _11332_ VGND VGND VPWR VPWR _02050_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21254_ net117 _08117_ _08118_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20205_ net106 systolic_inst.acc_wires\[6\]\[28\] net68 _07169_ VGND VGND VPWR VPWR
+ _01582_ sky130_fd_sc_hd__a22o_1
XFILLER_137_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21185_ _08052_ _08053_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__xnor2_1
X_28850_ clknet_leaf_337_clk _02648_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[398\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20136_ _07109_ _07110_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__nand2_1
X_27801_ clknet_leaf_48_clk _01599_ net137 VGND VGND VPWR VPWR systolic_inst.B_outs\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_28781_ clknet_leaf_230_clk _02579_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[329\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25993_ systolic_inst.acc_wires\[14\]\[21\] ser_C.parallel_data\[469\] net25 VGND
+ VGND VPWR VPWR _03295_ sky130_fd_sc_hd__mux2_1
XFILLER_213_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27732_ clknet_leaf_144_clk _01530_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_20067_ _07049_ _07050_ net68 VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__o21ai_1
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24944_ net111 ser_C.shift_reg\[300\] VGND VGND VPWR VPWR _10942_ sky130_fd_sc_hd__and2_1
XFILLER_219_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27663_ clknet_leaf_202_clk _01461_ net147 VGND VGND VPWR VPWR systolic_inst.A_outs\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24875_ C_out\[264\] net101 net73 ser_C.shift_reg\[264\] _10907_ VGND VGND VPWR VPWR
+ _02514_ sky130_fd_sc_hd__a221o_1
XFILLER_234_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26614_ clknet_leaf_17_B_in_serial_clk _00417_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29402_ clknet_leaf_238_clk _03200_ net146 VGND VGND VPWR VPWR C_out\[374\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23826_ _10419_ _10421_ _10422_ VGND VGND VPWR VPWR _10423_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_124_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27594_ clknet_leaf_224_clk _01392_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_205_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29333_ clknet_leaf_220_clk _03131_ net140 VGND VGND VPWR VPWR C_out\[305\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26545_ clknet_leaf_20_A_in_serial_clk _00348_ net131 VGND VGND VPWR VPWR deser_A.shift_reg\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_23757_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[0\]\[9\]
+ _10359_ VGND VGND VPWR VPWR _10364_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_146_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_120_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20969_ _07805_ _07842_ VGND VGND VPWR VPWR _07843_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13510_ deser_A.shift_reg\[74\] deser_A.shift_reg\[75\] net129 VGND VGND VPWR VPWR
+ _00347_ sky130_fd_sc_hd__mux2_1
X_22708_ systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[3\]
+ systolic_inst.B_outs\[1\]\[0\] VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__a22o_1
XFILLER_159_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29264_ clknet_leaf_191_clk _03062_ net146 VGND VGND VPWR VPWR C_out\[236\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26476_ clknet_leaf_14_A_in_serial_clk _00279_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14490_ _11637_ _11639_ _11670_ VGND VGND VPWR VPWR _11671_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_81_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23688_ _10285_ _10290_ _10297_ _10298_ net121 VGND VGND VPWR VPWR _10306_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_81_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Left_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28215_ clknet_leaf_84_clk _02013_ VGND VGND VPWR VPWR systolic_inst.B_shift\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_186_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13441_ deser_A.shift_reg\[5\] deser_A.shift_reg\[6\] deser_A.receiving VGND VGND
+ VPWR VPWR _00278_ sky130_fd_sc_hd__mux2_1
X_25427_ systolic_inst.A_shift\[1\]\[5\] A_in\[5\] net59 VGND VGND VPWR VPWR _11183_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22639_ _09348_ _09349_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__nand2_1
X_29195_ clknet_leaf_215_clk _02993_ net149 VGND VGND VPWR VPWR C_out\[167\] sky130_fd_sc_hd__dfrtp_1
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_230_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28146_ clknet_leaf_100_clk _01944_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_16160_ _03513_ _03543_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__xor2_1
X_25358_ net112 ser_C.shift_reg\[507\] VGND VGND VPWR VPWR _11149_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13372_ A_in\[81\] deser_A.word_buffer\[81\] net95 VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload19 clknet_5_21__leaf_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__clkinv_8
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15111_ _12226_ _12227_ VGND VGND VPWR VPWR _12228_ sky130_fd_sc_hd__and2b_1
XFILLER_70_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24309_ systolic_inst.A_shift\[11\]\[2\] A_in\[42\] net59 VGND VGND VPWR VPWR _10628_
+ sky130_fd_sc_hd__mux2_1
X_28077_ clknet_leaf_121_clk _01875_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_182_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16091_ _13063_ _13065_ _13064_ VGND VGND VPWR VPWR _13086_ sky130_fd_sc_hd__o21ba_1
X_25289_ ser_C.parallel_data\[471\] net102 net74 ser_C.shift_reg\[471\] _11114_ VGND
+ VGND VPWR VPWR _02721_ sky130_fd_sc_hd__a221o_1
XFILLER_182_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27028_ clknet_leaf_11_B_in_serial_clk _00826_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15042_ _12107_ _12125_ _12124_ VGND VGND VPWR VPWR _12161_ sky130_fd_sc_hd__o21a_1
XFILLER_155_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19850_ _06813_ _06818_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18801_ net115 _05920_ _05921_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19781_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[7\]
+ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__o21a_1
X_28979_ clknet_leaf_19_clk _02777_ VGND VGND VPWR VPWR systolic_inst.A_shift\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16993_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[11\]\[4\]
+ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18732_ _05853_ _05854_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__nand2_1
X_15944_ _12958_ _12961_ _12960_ VGND VGND VPWR VPWR _12965_ sky130_fd_sc_hd__o21a_1
XFILLER_95_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15875_ _12897_ _12899_ _12906_ VGND VGND VPWR VPWR _12907_ sky130_fd_sc_hd__a21oi_1
X_18663_ _05732_ _05788_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_237_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_237_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_237_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14826_ _11950_ VGND VGND VPWR VPWR _11951_ sky130_fd_sc_hd__inv_2
XFILLER_64_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17614_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[10\]\[6\]
+ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__or2_1
XFILLER_188_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18594_ _05683_ _05685_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14757_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[0\] _11886_
+ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_47_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _11275_ systolic_inst.A_outs\[10\]\[7\] _04746_ _04771_ VGND VGND VPWR VPWR
+ _04796_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_137_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_233_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13708_ B_in\[15\] deser_B.word_buffer\[15\] net84 VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17476_ _04729_ _04728_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__and2b_1
X_14688_ _11821_ _11828_ _11833_ _11838_ VGND VGND VPWR VPWR _11842_ sky130_fd_sc_hd__nand4_1
X_19215_ systolic_inst.B_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[5\]
+ systolic_inst.A_outs\[7\]\[6\] VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__and4_1
X_13639_ deser_B.word_buffer\[75\] deser_B.serial_word\[75\] net123 VGND VGND VPWR
+ VPWR _00476_ sky130_fd_sc_hd__mux2_1
X_16427_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[12\]\[10\]
+ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__and2_1
XFILLER_203_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19146_ _06208_ _06211_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__xnor2_1
X_16358_ _03516_ _03657_ _03727_ _03725_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__a31o_1
XFILLER_34_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_184_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15309_ _12378_ _12398_ VGND VGND VPWR VPWR _12399_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_184_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19077_ _06125_ _06127_ _06126_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__a21bo_1
X_16289_ _03632_ _03669_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18028_ _05191_ _05192_ _05193_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__o21ba_1
XFILLER_195_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19979_ _06944_ _06949_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__and2_1
XFILLER_140_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22990_ _09634_ _09636_ _09666_ VGND VGND VPWR VPWR _09667_ sky130_fd_sc_hd__a21o_1
XFILLER_132_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21941_ net106 systolic_inst.acc_wires\[3\]\[11\] _08729_ _08730_ VGND VGND VPWR
+ VPWR _01757_ sky130_fd_sc_hd__a22o_1
XFILLER_67_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24660_ net7 ser_C.shift_reg\[158\] VGND VGND VPWR VPWR _10800_ sky130_fd_sc_hd__and2_1
XFILLER_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21872_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[3\]\[1\]
+ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__or2_1
XFILLER_43_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23611_ _10080_ _10198_ VGND VGND VPWR VPWR _10232_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_137_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[31\]
+ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__xnor2_1
X_24591_ C_out\[122\] net100 net82 ser_C.shift_reg\[122\] _10765_ VGND VGND VPWR VPWR
+ _02372_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_128_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_137_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26330_ clknet_leaf_15_A_in_serial_clk _00004_ net143 VGND VGND VPWR VPWR deser_A.receiving
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_223_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23542_ _10158_ _10163_ VGND VGND VPWR VPWR _10165_ sky130_fd_sc_hd__and2_1
XFILLER_39_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20754_ _07641_ _07662_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26261_ clknet_leaf_5_A_in_serial_clk _00069_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_23473_ _10094_ _10095_ _10030_ _10032_ VGND VGND VPWR VPWR _10098_ sky130_fd_sc_hd__o211ai_2
X_20685_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[5\]\[9\]
+ _07599_ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__a21oi_1
X_28000_ clknet_leaf_152_clk _01798_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25212_ net110 ser_C.shift_reg\[434\] VGND VGND VPWR VPWR _11076_ sky130_fd_sc_hd__and2_1
X_22424_ _09162_ _09163_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__nand2_1
XFILLER_104_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26192_ ser_C.bit_idx\[8\] _11300_ VGND VGND VPWR VPWR _11256_ sky130_fd_sc_hd__nor2_1
XFILLER_104_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25143_ C_out\[398\] net101 net73 ser_C.shift_reg\[398\] _11041_ VGND VGND VPWR VPWR
+ _02648_ sky130_fd_sc_hd__a221o_1
X_22355_ systolic_inst.B_outs\[2\]\[5\] systolic_inst.A_outs\[2\]\[6\] VGND VGND VPWR
+ VPWR _09097_ sky130_fd_sc_hd__nand2_1
XFILLER_152_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_300_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_300_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_87_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21306_ _08155_ _08157_ _08161_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__a21o_1
X_25074_ net112 ser_C.shift_reg\[365\] VGND VGND VPWR VPWR _11007_ sky130_fd_sc_hd__and2_1
X_22286_ systolic_inst.A_outs\[2\]\[4\] systolic_inst.B_outs\[2\]\[5\] VGND VGND VPWR
+ VPWR _09030_ sky130_fd_sc_hd__nand2_1
XFILLER_152_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24025_ systolic_inst.B_shift\[8\]\[0\] B_in\[32\] _00008_ VGND VGND VPWR VPWR _10530_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28902_ clknet_leaf_273_clk _02700_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[450\]
+ sky130_fd_sc_hd__dfrtp_1
X_21237_ _08079_ _08081_ _08103_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__a21oi_1
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28833_ clknet_leaf_237_clk _02631_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21168_ _08002_ _08004_ _08035_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__or3_1
XFILLER_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20119_ _07086_ _07091_ _07095_ net60 VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__a31o_1
XFILLER_77_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13990_ deser_B.shift_reg\[24\] deser_B.shift_reg\[25\] net125 VGND VGND VPWR VPWR
+ _00816_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28764_ clknet_leaf_214_clk _02562_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[312\]
+ sky130_fd_sc_hd__dfrtp_1
X_21099_ _07967_ _07968_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__xor2_1
X_25976_ systolic_inst.acc_wires\[14\]\[4\] ser_C.parallel_data\[452\] net24 VGND
+ VGND VPWR VPWR _03278_ sky130_fd_sc_hd__mux2_1
XFILLER_120_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27715_ clknet_leaf_190_clk _01513_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24927_ C_out\[290\] net102 net74 ser_C.shift_reg\[290\] _10933_ VGND VGND VPWR VPWR
+ _02540_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_122_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28695_ clknet_leaf_193_clk _02493_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[243\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15660_ _12576_ _12712_ VGND VGND VPWR VPWR _12714_ sky130_fd_sc_hd__nand2_2
X_24858_ net110 ser_C.shift_reg\[257\] VGND VGND VPWR VPWR _10899_ sky130_fd_sc_hd__and2_1
X_27646_ clknet_leaf_314_clk _01444_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14611_ _11774_ _11775_ _11776_ VGND VGND VPWR VPWR _11777_ sky130_fd_sc_hd__and3_1
X_23809_ _10406_ _10408_ VGND VGND VPWR VPWR _10409_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_1174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_232_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15591_ systolic_inst.B_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[6\] systolic_inst.A_outs\[13\]\[7\]
+ systolic_inst.B_outs\[13\]\[3\] VGND VGND VPWR VPWR _12647_ sky130_fd_sc_hd__a22o_1
X_27577_ clknet_leaf_221_clk _01375_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_24789_ C_out\[221\] net99 net79 ser_C.shift_reg\[221\] _10864_ VGND VGND VPWR VPWR
+ _02471_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_164_Left_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_232_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_232_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17330_ _04571_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14542_ _11715_ _11716_ _11717_ VGND VGND VPWR VPWR _11718_ sky130_fd_sc_hd__a21o_1
X_29316_ clknet_leaf_300_clk _03114_ net139 VGND VGND VPWR VPWR C_out\[288\] sky130_fd_sc_hd__dfrtp_1
X_26528_ clknet_leaf_5_A_in_serial_clk _00331_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17261_ _04511_ _04520_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__nor2_1
XFILLER_109_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29247_ clknet_leaf_185_clk _03045_ net146 VGND VGND VPWR VPWR C_out\[219\] sky130_fd_sc_hd__dfrtp_1
X_14473_ _11652_ _11653_ VGND VGND VPWR VPWR _11654_ sky130_fd_sc_hd__nor2_1
X_26459_ clknet_leaf_11_clk _00266_ net132 VGND VGND VPWR VPWR A_in\[127\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16212_ systolic_inst.A_outs\[12\]\[6\] _03594_ _03593_ VGND VGND VPWR VPWR _03595_
+ sky130_fd_sc_hd__a21bo_1
X_19000_ _06081_ _06084_ _06087_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__o31a_1
X_13424_ _11309_ _11311_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__nor2_1
X_29178_ clknet_leaf_136_clk _02976_ net142 VGND VGND VPWR VPWR C_out\[150\] sky130_fd_sc_hd__dfrtp_1
X_17192_ systolic_inst.B_outs\[9\]\[6\] systolic_inst.B_outs\[5\]\[6\] net116 VGND
+ VGND VPWR VPWR _01280_ sky130_fd_sc_hd__mux2_1
XFILLER_167_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload108 clknet_leaf_282_clk VGND VGND VPWR VPWR clkload108/Y sky130_fd_sc_hd__bufinv_16
X_28129_ clknet_leaf_121_clk _01927_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16143_ systolic_inst.A_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[2\] systolic_inst.B_outs\[12\]\[6\]
+ systolic_inst.B_outs\[12\]\[7\] VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__and4b_1
Xclkload119 clknet_leaf_292_clk VGND VGND VPWR VPWR clkload119/X sky130_fd_sc_hd__clkbuf_4
X_13355_ A_in\[64\] deser_A.word_buffer\[64\] net94 VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__mux2_1
XFILLER_220_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16074_ _13035_ _13069_ VGND VGND VPWR VPWR _13070_ sky130_fd_sc_hd__nor2_1
X_13286_ deser_A.word_buffer\[124\] deser_A.serial_word\[124\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_226_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_173_Left_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_226_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_14__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_14__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_19902_ _06896_ _06899_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__xnor2_1
X_15025_ systolic_inst.B_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\] VGND VGND
+ VPWR VPWR _12144_ sky130_fd_sc_hd__or2_1
XFILLER_68_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19833_ _06831_ _06832_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__nor2_1
XFILLER_122_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_239_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_239_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19764_ _06729_ _06764_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__and2_1
XFILLER_42_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16976_ _04287_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__inv_2
XFILLER_232_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18715_ _05838_ _05839_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__xnor2_1
Xinput6 start VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_4
X_15927_ _12942_ _12944_ _12950_ VGND VGND VPWR VPWR _12951_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_177_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19695_ _06693_ _06698_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_177_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18646_ systolic_inst.A_outs\[8\]\[4\] systolic_inst.B_outs\[8\]\[6\] _11259_ systolic_inst.A_outs\[8\]\[3\]
+ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__o2bb2a_1
X_15858_ _12876_ _12883_ _12889_ _12882_ VGND VGND VPWR VPWR _12892_ sky130_fd_sc_hd__a211o_1
XFILLER_225_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_182_Left_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14809_ _11913_ _11915_ _11914_ VGND VGND VPWR VPWR _11934_ sky130_fd_sc_hd__a21bo_1
XFILLER_75_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18577_ systolic_inst.A_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[2\] systolic_inst.B_outs\[8\]\[6\]
+ systolic_inst.B_outs\[8\]\[7\] VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__and4b_1
X_15789_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[13\]\[6\]
+ VGND VGND VPWR VPWR _12833_ sky130_fd_sc_hd__or2_1
XFILLER_36_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17528_ _04714_ _04778_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__or2_1
XFILLER_177_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17459_ _04676_ _04712_ systolic_inst.A_outs\[10\]\[7\] VGND VGND VPWR VPWR _04713_
+ sky130_fd_sc_hd__and3b_1
XFILLER_127_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20470_ _07401_ _07404_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__xnor2_1
X_19129_ _06194_ _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__nor2_1
XFILLER_69_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_191_Left_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22140_ _08870_ _08886_ _08887_ VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__and3_1
XFILLER_161_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22071_ _08840_ _08841_ _08829_ _08835_ _08839_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__a2111o_1
XFILLER_195_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21022_ _07892_ _07893_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__xor2_1
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25830_ systolic_inst.acc_wires\[9\]\[18\] C_out\[306\] net15 VGND VGND VPWR VPWR
+ _03132_ sky130_fd_sc_hd__mux2_1
XFILLER_87_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25761_ systolic_inst.acc_wires\[7\]\[13\] C_out\[237\] net43 VGND VGND VPWR VPWR
+ _03063_ sky130_fd_sc_hd__mux2_1
XFILLER_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22973_ _09649_ _09650_ VGND VGND VPWR VPWR _09651_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24712_ net113 ser_C.shift_reg\[184\] VGND VGND VPWR VPWR _10826_ sky130_fd_sc_hd__and2_1
XFILLER_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27500_ clknet_leaf_296_clk _01298_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28480_ clknet_leaf_109_clk _02278_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21924_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[3\]\[8\]
+ _08711_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__a21oi_1
X_25692_ systolic_inst.acc_wires\[5\]\[8\] C_out\[168\] net31 VGND VGND VPWR VPWR
+ _02994_ sky130_fd_sc_hd__mux2_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27431_ clknet_leaf_242_clk _01229_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_182_Right_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24643_ C_out\[148\] net104 net76 ser_C.shift_reg\[148\] _10791_ VGND VGND VPWR VPWR
+ _02398_ sky130_fd_sc_hd__a221o_1
XFILLER_231_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21855_ _08607_ _08636_ VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__nor2_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20806_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[28\]
+ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__nand2_1
XFILLER_19_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27362_ clknet_leaf_341_clk _01160_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24574_ net113 ser_C.shift_reg\[115\] VGND VGND VPWR VPWR _10757_ sky130_fd_sc_hd__and2_1
X_21786_ systolic_inst.B_outs\[3\]\[5\] systolic_inst.A_outs\[3\]\[7\] _08589_ VGND
+ VGND VPWR VPWR _08591_ sky130_fd_sc_hd__and3_1
X_29101_ clknet_leaf_154_clk _02899_ net150 VGND VGND VPWR VPWR C_out\[73\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26313_ clknet_leaf_28_A_in_serial_clk _00121_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_23525_ _10144_ _10147_ VGND VGND VPWR VPWR _10148_ sky130_fd_sc_hd__or2_1
XFILLER_54_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20737_ _07646_ _07648_ VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27293_ clknet_leaf_291_clk _01091_ net141 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29032_ clknet_leaf_126_clk _02830_ net144 VGND VGND VPWR VPWR C_out\[4\] sky130_fd_sc_hd__dfrtp_1
X_26244_ clknet_leaf_11_A_in_serial_clk _00052_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_23456_ systolic_inst.A_outs\[0\]\[6\] _10080_ _10079_ VGND VGND VPWR VPWR _10081_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20668_ _07586_ _07587_ _07588_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__a21o_1
XFILLER_17_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22407_ _09146_ _09147_ VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26175_ net7 ser_C.bit_idx\[0\] ser_C.bit_idx\[1\] VGND VGND VPWR VPWR _11246_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_115_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23387_ _09968_ _09969_ _09981_ _09980_ _09979_ VGND VGND VPWR VPWR _10014_ sky130_fd_sc_hd__a32o_1
XFILLER_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20599_ _07528_ _07529_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__nor2_1
XFILLER_104_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13140_ systolic_inst.cycle_cnt\[30\] systolic_inst.cycle_cnt\[31\] systolic_inst.cycle_cnt\[29\]
+ systolic_inst.cycle_cnt\[28\] VGND VGND VPWR VPWR _11293_ sky130_fd_sc_hd__or4_1
XFILLER_152_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25126_ net110 ser_C.shift_reg\[391\] VGND VGND VPWR VPWR _11033_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22338_ _09022_ _09080_ VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25057_ C_out\[355\] net98 net78 ser_C.shift_reg\[355\] _10998_ VGND VGND VPWR VPWR
+ _02605_ sky130_fd_sc_hd__a221o_1
X_22269_ _08973_ _08975_ VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__and2_1
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24008_ _10529_ systolic_inst.B_shift\[5\]\[7\] _11332_ VGND VGND VPWR VPWR _02025_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_221_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_221_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16830_ _04096_ _04115_ _04114_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__o21ba_1
X_28816_ clknet_leaf_241_clk _02614_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[364\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13973_ deser_B.shift_reg\[7\] deser_B.shift_reg\[8\] net125 VGND VGND VPWR VPWR
+ _00799_ sky130_fd_sc_hd__mux2_1
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16761_ _04079_ _04080_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__xor2_1
X_28747_ clknet_leaf_298_clk _02545_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[295\]
+ sky130_fd_sc_hd__dfrtp_1
X_25959_ systolic_inst.acc_wires\[13\]\[19\] C_out\[435\] net20 VGND VGND VPWR VPWR
+ _03261_ sky130_fd_sc_hd__mux2_1
XFILLER_47_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18500_ _05626_ _05629_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_234_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15712_ _12714_ _12764_ VGND VGND VPWR VPWR _12765_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19480_ _06515_ _06520_ _06521_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__nand3_1
X_16692_ _04013_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__nor2_1
XFILLER_234_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28678_ clknet_leaf_197_clk _02476_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[226\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18431_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[2\] _05565_ VGND
+ VGND VPWR VPWR _05566_ sky130_fd_sc_hd__nand3_1
XFILLER_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15643_ _12657_ _12659_ _12697_ VGND VGND VPWR VPWR _12698_ sky130_fd_sc_hd__a21o_1
X_27629_ clknet_leaf_323_clk _01427_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_222_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18362_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[25\]
+ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__xor2_2
X_15574_ _12629_ _12630_ VGND VGND VPWR VPWR _12631_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_29_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14525_ _11694_ _11697_ net118 _11693_ VGND VGND VPWR VPWR _11704_ sky130_fd_sc_hd__o211a_1
X_17313_ _04533_ _04570_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18293_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[15\]
+ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__and2_1
XFILLER_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _11635_ _11636_ VGND VGND VPWR VPWR _11638_ sky130_fd_sc_hd__xnor2_1
X_17244_ _04475_ _04492_ _04494_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_228_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13407_ A_in\[116\] deser_A.word_buffer\[116\] _00003_ VGND VGND VPWR VPWR _00255_
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17175_ _04451_ _04455_ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__a21oi_1
X_14387_ _11569_ _11570_ VGND VGND VPWR VPWR _11571_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_210_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16126_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[7\] VGND
+ VGND VPWR VPWR _03512_ sky130_fd_sc_hd__nand2_1
XFILLER_196_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13338_ A_in\[47\] deser_A.word_buffer\[47\] net93 VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__mux2_1
XFILLER_170_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16057_ _13052_ _13051_ VGND VGND VPWR VPWR _13054_ sky130_fd_sc_hd__nand2b_1
X_13269_ deser_A.word_buffer\[107\] deser_A.serial_word\[107\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15008_ _12127_ _12126_ VGND VGND VPWR VPWR _12128_ sky130_fd_sc_hd__nand2b_1
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19816_ _06774_ _06777_ _06815_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__or3_1
XFILLER_233_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19747_ _06743_ _06747_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__and2_1
XFILLER_56_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16959_ _04271_ _04273_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__nand2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19678_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[4\] VGND
+ VGND VPWR VPWR _06683_ sky130_fd_sc_hd__and2_1
XFILLER_237_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18629_ _05719_ _05721_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__a21o_1
XFILLER_37_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21640_ systolic_inst.B_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[5\]
+ systolic_inst.B_outs\[3\]\[3\] VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__a22oi_1
XFILLER_80_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21571_ systolic_inst.A_outs\[3\]\[2\] systolic_inst.B_outs\[3\]\[3\] systolic_inst.A_outs\[3\]\[3\]
+ systolic_inst.B_outs\[3\]\[4\] VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_155_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_11 systolic_inst.B_outs\[3\]\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_22 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23310_ _09925_ _09938_ VGND VGND VPWR VPWR _09940_ sky130_fd_sc_hd__nand2_1
XFILLER_162_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_33 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20522_ _07455_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__inv_2
XANTENNA_44 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24290_ _10618_ systolic_inst.A_shift\[11\]\[0\] net71 VGND VGND VPWR VPWR _02218_
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23241_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[26\]
+ VGND VGND VPWR VPWR _09888_ sky130_fd_sc_hd__or2_1
XFILLER_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20453_ _07353_ _07356_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__nand2_1
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23172_ _09828_ _09829_ VGND VGND VPWR VPWR _09830_ sky130_fd_sc_hd__or2_1
XFILLER_174_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20384_ systolic_inst.B_outs\[5\]\[3\] systolic_inst.A_outs\[5\]\[4\] _07298_ _07297_
+ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__a31o_1
XFILLER_238_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22123_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[2\] VGND VGND VPWR
+ VPWR _08872_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_164_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27980_ clknet_leaf_118_clk _01778_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_122_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22054_ _08817_ _08826_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__nor2_1
X_26931_ clknet_leaf_17_A_in_serial_clk _00729_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21005_ _07837_ _07876_ _07875_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__o21a_1
XFILLER_212_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29650_ clknet_leaf_5_B_in_serial_clk _03445_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_26862_ clknet_leaf_0_B_in_serial_clk _00664_ net134 VGND VGND VPWR VPWR deser_B.bit_idx\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28601_ clknet_leaf_137_clk _02399_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[149\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25813_ systolic_inst.acc_wires\[9\]\[1\] C_out\[289\] net14 VGND VGND VPWR VPWR
+ _03115_ sky130_fd_sc_hd__mux2_1
XFILLER_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26793_ clknet_leaf_72_clk _00595_ net153 VGND VGND VPWR VPWR B_in\[65\] sky130_fd_sc_hd__dfrtp_1
X_29581_ clknet_leaf_20_B_in_serial_clk _03376_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28532_ clknet_leaf_162_clk _02330_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_25744_ systolic_inst.acc_wires\[6\]\[28\] C_out\[220\] net43 VGND VGND VPWR VPWR
+ _03046_ sky130_fd_sc_hd__mux2_1
Xmax_cap13 net16 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_4
X_22956_ _09633_ _09632_ VGND VGND VPWR VPWR _09634_ sky130_fd_sc_hd__nand2b_1
XFILLER_29_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap24 net25 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_8
Xmax_cap35 net36 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_4
XFILLER_216_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap46 net48 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_3_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21907_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[3\]\[6\]
+ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__or2_1
Xmax_cap57 _00002_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_104_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28463_ clknet_leaf_122_clk _02261_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_25675_ systolic_inst.acc_wires\[4\]\[23\] C_out\[151\] net32 VGND VGND VPWR VPWR
+ _02977_ sky130_fd_sc_hd__mux2_1
Xmax_cap68 _11712_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_104_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap79 net80 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_12
X_22887_ systolic_inst.A_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[5\] _09529_ _09528_
+ VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__a31oi_1
XFILLER_203_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27414_ clknet_leaf_214_clk _01212_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_24626_ net110 ser_C.shift_reg\[141\] VGND VGND VPWR VPWR _10783_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21838_ systolic_inst.A_outs\[3\]\[6\] _11274_ _08615_ _08618_ _08640_ VGND VGND
+ VPWR VPWR _08641_ sky130_fd_sc_hd__o311a_1
X_28394_ clknet_leaf_32_clk _02192_ VGND VGND VPWR VPWR systolic_inst.A_shift\[17\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27345_ clknet_leaf_343_clk _01143_ net131 VGND VGND VPWR VPWR systolic_inst.A_outs\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_24557_ C_out\[105\] net99 net80 ser_C.shift_reg\[105\] _10748_ VGND VGND VPWR VPWR
+ _02355_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_117_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21769_ _08538_ _08540_ _08574_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__and3_1
XFILLER_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14310_ _11486_ _11495_ VGND VGND VPWR VPWR _11496_ sky130_fd_sc_hd__xnor2_1
X_23508_ _10113_ _10130_ _10131_ VGND VGND VPWR VPWR _10132_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_78_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15290_ _12374_ _12379_ _12381_ VGND VGND VPWR VPWR _12383_ sky130_fd_sc_hd__a21oi_1
X_27276_ clknet_leaf_325_clk _01074_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_78_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24488_ net112 ser_C.shift_reg\[72\] VGND VGND VPWR VPWR _10714_ sky130_fd_sc_hd__and2_1
XFILLER_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29015_ clknet_leaf_93_clk _02813_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_200_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26227_ clknet_leaf_8_A_in_serial_clk _00035_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14241_ _11425_ _11427_ _11403_ VGND VGND VPWR VPWR _11429_ sky130_fd_sc_hd__a21oi_1
X_23439_ systolic_inst.B_outs\[0\]\[7\] _10026_ _10027_ VGND VGND VPWR VPWR _10064_
+ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_20_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26158_ deser_B.serial_word\[113\] deser_B.shift_reg\[113\] net55 VGND VGND VPWR
+ VPWR _03460_ sky130_fd_sc_hd__mux2_1
X_14172_ _11351_ _11361_ VGND VGND VPWR VPWR _11362_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_223_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13123_ B_in_valid A_in_valid net6 _11258_ VGND VGND VPWR VPWR _11279_ sky130_fd_sc_hd__nand4_4
XFILLER_124_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25109_ C_out\[381\] net99 net79 ser_C.shift_reg\[381\] _11024_ VGND VGND VPWR VPWR
+ _02631_ sky130_fd_sc_hd__a221o_1
X_26089_ deser_B.serial_word\[44\] deser_B.shift_reg\[44\] net55 VGND VGND VPWR VPWR
+ _03391_ sky130_fd_sc_hd__mux2_1
XFILLER_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18980_ _06072_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17931_ systolic_inst.A_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[7\] VGND VGND VPWR
+ VPWR _05125_ sky130_fd_sc_hd__and2b_1
XFILLER_117_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17862_ _05036_ _05056_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19601_ _06618_ _06621_ _06624_ _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__o31a_1
XFILLER_113_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16813_ systolic_inst.B_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[7\]
+ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__and3_1
XFILLER_19_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17793_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[4\]\[0\] net121 VGND
+ VGND VPWR VPWR _01338_ sky130_fd_sc_hd__mux2_1
XFILLER_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19532_ _06565_ _06567_ _06564_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_50_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16744_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[6\] VGND VGND
+ VPWR VPWR _04065_ sky130_fd_sc_hd__nand2_1
X_13956_ deser_A.serial_word\[117\] deser_A.shift_reg\[117\] _00002_ VGND VGND VPWR
+ VPWR _00782_ sky130_fd_sc_hd__mux2_1
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19463_ _06504_ _06507_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__and2_1
XFILLER_35_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16675_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[4\] _03995_ _03996_
+ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__a22o_1
X_13887_ deser_A.serial_word\[48\] deser_A.shift_reg\[48\] net58 VGND VGND VPWR VPWR
+ _00713_ sky130_fd_sc_hd__mux2_1
XFILLER_235_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18414_ systolic_inst.B_outs\[7\]\[3\] systolic_inst.B_outs\[3\]\[3\] net119 VGND
+ VGND VPWR VPWR _01405_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ systolic_inst.A_outs\[13\]\[6\] _12648_ _12649_ _12616_ VGND VGND VPWR VPWR
+ _12681_ sky130_fd_sc_hd__o2bb2a_1
X_19394_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[14\] _06452_ net119
+ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__mux2_1
XFILLER_222_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18345_ _05504_ _05505_ _05506_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__or3_1
X_15557_ _12577_ _12612_ VGND VGND VPWR VPWR _12614_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_212_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_212_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_72_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14508_ _11687_ _11686_ VGND VGND VPWR VPWR _11688_ sky130_fd_sc_hd__and2b_1
XFILLER_187_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15488_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[5\] VGND VGND
+ VPWR VPWR _12547_ sky130_fd_sc_hd__nand2_1
X_18276_ _05445_ _05448_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_13_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17227_ systolic_inst.B_outs\[10\]\[4\] _04474_ _04487_ VGND VGND VPWR VPWR _04488_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_128_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14439_ _11620_ VGND VGND VPWR VPWR _11621_ sky130_fd_sc_hd__inv_2
XFILLER_239_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17158_ _04441_ _04442_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__nand2_1
XFILLER_115_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16109_ _13100_ _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17089_ net105 systolic_inst.acc_wires\[11\]\[17\] net62 _04384_ VGND VGND VPWR VPWR
+ _01251_ sky130_fd_sc_hd__a22o_1
XFILLER_157_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_206_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_206_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_198_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22810_ _09490_ _09491_ VGND VGND VPWR VPWR _09492_ sky130_fd_sc_hd__and2b_1
XFILLER_38_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23790_ _10389_ _10391_ VGND VGND VPWR VPWR _10393_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22741_ _09423_ _09424_ VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__nor2_1
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25460_ _00008_ _11203_ VGND VGND VPWR VPWR _11204_ sky130_fd_sc_hd__nor2_1
XFILLER_80_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22672_ _09377_ _09376_ systolic_inst.acc_wires\[2\]\[31\] net109 VGND VGND VPWR
+ VPWR _01841_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_240_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24411_ C_out\[32\] _11302_ net81 ser_C.shift_reg\[32\] _10675_ VGND VGND VPWR VPWR
+ _02282_ sky130_fd_sc_hd__a221o_1
XFILLER_197_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21623_ _08403_ _08432_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__nand2b_1
XFILLER_240_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25391_ systolic_inst.A_shift\[3\]\[3\] A_in\[19\] net59 VGND VGND VPWR VPWR _11165_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
X_27130_ clknet_leaf_12_clk _00928_ VGND VGND VPWR VPWR systolic_inst.A_shift\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24342_ systolic_inst.A_shift\[8\]\[5\] net70 net83 systolic_inst.A_shift\[9\]\[5\]
+ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__a22o_1
XFILLER_240_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21554_ _08336_ _08364_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__or2_1
XFILLER_103_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27061_ clknet_leaf_6_B_in_serial_clk _00859_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_20505_ _07437_ _07438_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__or2_1
XFILLER_166_668 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24273_ systolic_inst.B_shift\[27\]\[0\] B_in\[88\] net59 VGND VGND VPWR VPWR _10610_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21485_ net122 _08300_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__and2_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26012_ systolic_inst.acc_wires\[15\]\[8\] ser_C.parallel_data\[488\] net39 VGND
+ VGND VPWR VPWR _03314_ sky130_fd_sc_hd__mux2_1
X_23224_ _09866_ _09870_ _09873_ VGND VGND VPWR VPWR _09874_ sky130_fd_sc_hd__nand3_1
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20436_ _07370_ _07371_ VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__nor2_1
XFILLER_140_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23155_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[1\]\[12\]
+ _09812_ _09814_ VGND VGND VPWR VPWR _09815_ sky130_fd_sc_hd__a211o_1
XFILLER_180_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload280 clknet_leaf_207_clk VGND VGND VPWR VPWR clkload280/X sky130_fd_sc_hd__clkbuf_4
X_20367_ _07300_ _07303_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__xor2_1
XFILLER_88_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload291 clknet_leaf_198_clk VGND VGND VPWR VPWR clkload291/Y sky130_fd_sc_hd__inv_6
X_22106_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[2\] _08856_ VGND
+ VGND VPWR VPWR _08857_ sky130_fd_sc_hd__nand3_1
XFILLER_171_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23086_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[1\]\[3\]
+ VGND VGND VPWR VPWR _09756_ sky130_fd_sc_hd__or2_1
X_27963_ clknet_leaf_149_clk _01761_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_175_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20298_ systolic_inst.A_outs\[5\]\[2\] systolic_inst.B_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\]
+ systolic_inst.A_outs\[5\]\[1\] VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__a22oi_2
Xclkbuf_leaf_99_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_216_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22037_ _08807_ _08809_ _08811_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__o21ai_1
X_26914_ clknet_leaf_11_A_in_serial_clk _00712_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27894_ clknet_leaf_39_clk _01692_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_196_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29633_ clknet_leaf_11_B_in_serial_clk _03428_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26845_ clknet_leaf_68_clk _00647_ net153 VGND VGND VPWR VPWR B_in\[117\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13810_ B_in\[117\] deser_B.word_buffer\[117\] net87 VGND VGND VPWR VPWR _00647_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29564_ clknet_leaf_15_B_in_serial_clk _03359_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14790_ _11914_ _11915_ VGND VGND VPWR VPWR _11916_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23988_ _10519_ systolic_inst.B_shift\[8\]\[5\] net72 VGND VGND VPWR VPWR _02015_
+ sky130_fd_sc_hd__mux2_1
X_26776_ clknet_leaf_79_clk _00578_ net144 VGND VGND VPWR VPWR B_in\[48\] sky130_fd_sc_hd__dfrtp_1
XFILLER_235_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28515_ clknet_leaf_156_clk _02313_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_13741_ B_in\[48\] deser_B.word_buffer\[48\] net86 VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22939_ _09580_ _09616_ _09617_ VGND VGND VPWR VPWR _09618_ sky130_fd_sc_hd__and3_1
X_25727_ systolic_inst.acc_wires\[6\]\[11\] C_out\[203\] net47 VGND VGND VPWR VPWR
+ _03029_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29495_ clknet_leaf_269_clk _03293_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[467\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13672_ deser_B.word_buffer\[108\] deser_B.serial_word\[108\] net123 VGND VGND VPWR
+ VPWR _00509_ sky130_fd_sc_hd__mux2_1
X_16460_ net108 systolic_inst.acc_wires\[12\]\[13\] _03822_ _03823_ VGND VGND VPWR
+ VPWR _01183_ sky130_fd_sc_hd__a22o_1
X_28446_ clknet_leaf_35_clk _02244_ VGND VGND VPWR VPWR systolic_inst.A_shift\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25658_ systolic_inst.acc_wires\[4\]\[6\] C_out\[134\] net29 VGND VGND VPWR VPWR
+ _02960_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15411_ _12471_ _12472_ _12453_ VGND VGND VPWR VPWR _12473_ sky130_fd_sc_hd__o21ai_1
X_16391_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[12\]\[4\]
+ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__or2_1
XFILLER_58_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24609_ C_out\[131\] net103 net75 ser_C.shift_reg\[131\] _10774_ VGND VGND VPWR VPWR
+ _02381_ sky130_fd_sc_hd__a221o_1
XFILLER_223_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25589_ systolic_inst.acc_wires\[2\]\[1\] C_out\[65\] net34 VGND VGND VPWR VPWR _02891_
+ sky130_fd_sc_hd__mux2_1
X_28377_ clknet_leaf_3_clk _02175_ VGND VGND VPWR VPWR systolic_inst.A_shift\[19\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_197_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15342_ _12424_ _12426_ VGND VGND VPWR VPWR _12427_ sky130_fd_sc_hd__xnor2_1
X_18130_ _05317_ _05318_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__nor2_1
X_27328_ clknet_leaf_330_clk _01126_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_223_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15273_ _12366_ _12368_ VGND VGND VPWR VPWR _12369_ sky130_fd_sc_hd__xor2_1
X_18061_ _05180_ _05183_ _05213_ _05214_ _05250_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__a311oi_4
X_27259_ clknet_leaf_282_clk _01057_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_185_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14224_ systolic_inst.B_outs\[15\]\[3\] systolic_inst.A_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\]
+ systolic_inst.A_outs\[15\]\[2\] VGND VGND VPWR VPWR _11412_ sky130_fd_sc_hd__a22o_1
X_17012_ _04318_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14155_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[2\]
+ systolic_inst.A_outs\[15\]\[1\] VGND VGND VPWR VPWR _11346_ sky130_fd_sc_hd__a22o_1
XFILLER_193_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13106_ systolic_inst.B_outs\[11\]\[7\] VGND VGND VPWR VPWR _11262_ sky130_fd_sc_hd__inv_2
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14086_ deser_B.shift_reg\[120\] deser_B.shift_reg\[121\] deser_B.receiving VGND
+ VGND VPWR VPWR _00912_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18963_ systolic_inst.acc_wires\[8\]\[20\] systolic_inst.acc_wires\[8\]\[21\] systolic_inst.acc_wires\[8\]\[22\]
+ systolic_inst.acc_wires\[8\]\[23\] systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__o41a_1
XFILLER_79_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17914_ _05068_ _05099_ _05101_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__o21ba_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18894_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[8\]\[14\]
+ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__nand2_1
XFILLER_239_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17845_ _05034_ _05040_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__and2_1
XFILLER_94_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_201_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17776_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[30\]
+ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__or2_1
XFILLER_240_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14988_ systolic_inst.B_outs\[14\]\[4\] systolic_inst.A_outs\[14\]\[6\] systolic_inst.A_outs\[14\]\[7\]
+ systolic_inst.B_outs\[14\]\[3\] VGND VGND VPWR VPWR _12108_ sky130_fd_sc_hd__a22o_1
XFILLER_75_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19515_ _06554_ _06555_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__nand2_1
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16727_ _04017_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_193_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13939_ deser_A.serial_word\[100\] deser_A.shift_reg\[100\] net57 VGND VGND VPWR
+ VPWR _00765_ sky130_fd_sc_hd__mux2_1
XFILLER_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19446_ net62 _06494_ _06496_ systolic_inst.acc_wires\[7\]\[6\] net105 VGND VGND
+ VPWR VPWR _01496_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_18_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16658_ _03963_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_18_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15609_ _12646_ _12664_ VGND VGND VPWR VPWR _12665_ sky130_fd_sc_hd__xor2_1
XFILLER_222_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19377_ _06434_ _06435_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__nand2_1
XFILLER_241_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16589_ systolic_inst.B_outs\[10\]\[6\] systolic_inst.B_outs\[6\]\[6\] net120 VGND
+ VGND VPWR VPWR _01216_ sky130_fd_sc_hd__mux2_1
XFILLER_72_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_18328_ _05481_ _05486_ _05492_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__or3b_1
XFILLER_33_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18259_ net66 _05432_ _05433_ systolic_inst.acc_wires\[9\]\[10\] net107 VGND VGND
+ VPWR VPWR _01372_ sky130_fd_sc_hd__a32o_1
XFILLER_200_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21270_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[4\]\[3\]
+ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__nand2_1
XFILLER_239_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_208_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20221_ _07176_ _07180_ _07181_ net60 VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__a31o_1
XFILLER_11_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20152_ _07122_ _07123_ _07120_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__o21ai_2
XFILLER_172_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24960_ net110 ser_C.shift_reg\[308\] VGND VGND VPWR VPWR _10950_ sky130_fd_sc_hd__and2_1
XFILLER_83_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20083_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[6\]\[11\]
+ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23911_ _10488_ systolic_inst.B_shift\[13\]\[7\] net72 VGND VGND VPWR VPWR _01969_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24891_ C_out\[272\] net103 net75 ser_C.shift_reg\[272\] _10915_ VGND VGND VPWR VPWR
+ _02522_ sky130_fd_sc_hd__a221o_1
XFILLER_22_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23842_ _10435_ VGND VGND VPWR VPWR _10436_ sky130_fd_sc_hd__inv_2
X_26630_ clknet_leaf_19_B_in_serial_clk _00433_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23773_ _10375_ _10376_ _10377_ VGND VGND VPWR VPWR _10378_ sky130_fd_sc_hd__and3_1
X_26561_ clknet_leaf_2_A_in_serial_clk _00364_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20985_ _07816_ _07817_ _07858_ _07814_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__or4b_1
X_28300_ clknet_leaf_63_clk _02098_ VGND VGND VPWR VPWR systolic_inst.B_shift\[27\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25512_ systolic_inst.cycle_cnt\[28\] systolic_inst.cycle_cnt\[27\] systolic_inst.cycle_cnt\[26\]
+ _11233_ VGND VGND VPWR VPWR _11237_ sky130_fd_sc_hd__and4_1
X_22724_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[3\]
+ VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29280_ clknet_leaf_187_clk _03078_ net146 VGND VGND VPWR VPWR C_out\[252\] sky130_fd_sc_hd__dfrtp_1
X_26492_ clknet_leaf_6_A_in_serial_clk _00295_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_225_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25443_ _11189_ _11192_ _11191_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__a21oi_1
X_28231_ clknet_leaf_129_clk _02029_ VGND VGND VPWR VPWR systolic_inst.B_shift\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_22655_ net109 systolic_inst.acc_wires\[2\]\[28\] net65 _09363_ VGND VGND VPWR VPWR
+ _01838_ sky130_fd_sc_hd__a22o_1
XFILLER_80_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21606_ _08414_ _08415_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__or2_1
X_28162_ clknet_leaf_107_clk _01960_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_199_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25374_ _11156_ systolic_inst.B_shift\[14\]\[2\] net71 VGND VGND VPWR VPWR _02764_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22586_ _09303_ _09305_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27113_ clknet_leaf_30_B_in_serial_clk _00911_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24325_ systolic_inst.A_shift\[10\]\[2\] A_in\[34\] net59 VGND VGND VPWR VPWR _10636_
+ sky130_fd_sc_hd__mux2_1
X_28093_ clknet_leaf_112_clk _01891_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_21537_ _08347_ _08348_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__or2_1
XFILLER_103_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27044_ clknet_leaf_19_B_in_serial_clk _00842_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24256_ systolic_inst.A_shift\[17\]\[7\] net70 net83 systolic_inst.A_shift\[18\]\[7\]
+ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__a22o_1
X_21468_ systolic_inst.A_outs\[3\]\[4\] systolic_inst.A_outs\[2\]\[4\] net122 VGND
+ VGND VPWR VPWR _01718_ sky130_fd_sc_hd__mux2_1
XFILLER_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23207_ _09857_ _09858_ _09855_ VGND VGND VPWR VPWR _09860_ sky130_fd_sc_hd__o21ai_2
X_20419_ _07355_ _07354_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__nand2b_1
XFILLER_218_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24187_ systolic_inst.A_shift\[24\]\[2\] net70 _10505_ systolic_inst.A_shift\[25\]\[2\]
+ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__a22o_1
X_21399_ _08232_ _08239_ _08240_ _11713_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23138_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[1\]\[11\]
+ VGND VGND VPWR VPWR _09800_ sky130_fd_sc_hd__nor2_1
XFILLER_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28995_ clknet_leaf_47_clk _02793_ VGND VGND VPWR VPWR systolic_inst.A_shift\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23069_ net122 systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[1\]\[0\]
+ VGND VGND VPWR VPWR _09742_ sky130_fd_sc_hd__a21oi_1
X_27946_ clknet_leaf_148_clk _01744_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_15960_ systolic_inst.A_outs\[12\]\[1\] systolic_inst.A_shift\[24\]\[1\] net115 VGND
+ VGND VPWR VPWR _01139_ sky130_fd_sc_hd__mux2_1
XFILLER_89_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14911_ _12032_ _12029_ VGND VGND VPWR VPWR _12033_ sky130_fd_sc_hd__and2b_1
XFILLER_88_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15891_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[21\]
+ VGND VGND VPWR VPWR _12920_ sky130_fd_sc_hd__xnor2_2
X_27877_ clknet_leaf_38_clk _01675_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_29616_ clknet_leaf_2_B_in_serial_clk _03411_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_17630_ _04870_ _04869_ systolic_inst.acc_wires\[10\]\[8\] net105 VGND VGND VPWR
+ VPWR _01306_ sky130_fd_sc_hd__a2bb2o_1
X_26828_ clknet_leaf_86_clk _00630_ net135 VGND VGND VPWR VPWR B_in\[100\] sky130_fd_sc_hd__dfrtp_1
X_14842_ _11936_ _11965_ VGND VGND VPWR VPWR _11966_ sky130_fd_sc_hd__and2_1
XFILLER_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29547_ clknet_leaf_229_clk _03342_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_17561_ _04811_ _04810_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__nand2b_1
X_26759_ clknet_leaf_78_clk _00561_ net143 VGND VGND VPWR VPWR B_in\[31\] sky130_fd_sc_hd__dfrtp_1
X_14773_ systolic_inst.A_outs\[14\]\[0\] systolic_inst.A_outs\[14\]\[1\] systolic_inst.B_outs\[14\]\[2\]
+ systolic_inst.B_outs\[14\]\[3\] VGND VGND VPWR VPWR _11900_ sky130_fd_sc_hd__and4_1
XFILLER_229_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19300_ _06345_ _06361_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__xor2_1
XFILLER_189_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16512_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[20\]
+ _03866_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__a21bo_1
X_13724_ B_in\[31\] deser_B.word_buffer\[31\] net86 VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__mux2_1
XFILLER_189_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29478_ clknet_leaf_274_clk _03276_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[450\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17492_ _04743_ _04744_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__nor2_1
XFILLER_147_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19231_ _06257_ _06258_ _06260_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__o21a_1
XFILLER_71_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28429_ clknet_leaf_24_clk _02227_ VGND VGND VPWR VPWR systolic_inst.A_shift\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16443_ _03785_ _03790_ _03806_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__nand3_1
XFILLER_204_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13655_ deser_B.word_buffer\[91\] deser_B.serial_word\[91\] net124 VGND VGND VPWR
+ VPWR _00492_ sky130_fd_sc_hd__mux2_1
XFILLER_232_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19162_ _06199_ _06227_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__and2b_1
XFILLER_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13586_ deser_B.word_buffer\[22\] deser_B.serial_word\[22\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__mux2_1
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16374_ net67 _03748_ _03749_ systolic_inst.acc_wires\[12\]\[1\] net108 VGND VGND
+ VPWR VPWR _01171_ sky130_fd_sc_hd__a32o_1
XFILLER_83_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18113_ _05269_ _05271_ _05301_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__a21o_1
XFILLER_200_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15325_ _12410_ _12412_ VGND VGND VPWR VPWR _12413_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_41_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19093_ _06137_ _06160_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__nand2_1
XFILLER_200_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18044_ _05226_ _05234_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__nand2_1
X_15256_ _12341_ _12347_ _12348_ VGND VGND VPWR VPWR _12354_ sky130_fd_sc_hd__o21ba_1
XFILLER_173_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14207_ _11385_ _11394_ VGND VGND VPWR VPWR _11396_ sky130_fd_sc_hd__xor2_1
X_15187_ _12293_ _12294_ _12286_ _12290_ VGND VGND VPWR VPWR _12295_ sky130_fd_sc_hd__a211o_1
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14138_ systolic_inst.B_outs\[14\]\[6\] systolic_inst.B_outs\[10\]\[6\] net120 VGND
+ VGND VPWR VPWR _00960_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19995_ _06987_ _06988_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__and2b_1
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_203_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14069_ deser_B.shift_reg\[103\] deser_B.shift_reg\[104\] net126 VGND VGND VPWR VPWR
+ _00895_ sky130_fd_sc_hd__mux2_1
X_18946_ _06036_ _06042_ _06043_ net61 VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__a31o_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_234_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18877_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[8\]\[10\]
+ _05977_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__and3_1
XFILLER_95_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17828_ _05004_ _05010_ _05013_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__o21ai_1
XFILLER_227_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17759_ net105 systolic_inst.acc_wires\[10\]\[27\] net69 _04980_ VGND VGND VPWR VPWR
+ _01325_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_59_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20770_ _07673_ _07674_ _07675_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__or3_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19429_ _06480_ _06481_ _06473_ _06477_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__a211o_1
XFILLER_74_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22440_ _11265_ systolic_inst.A_outs\[2\]\[7\] _09130_ _09154_ VGND VGND VPWR VPWR
+ _09179_ sky130_fd_sc_hd__o211ai_1
XFILLER_149_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22371_ _09110_ _09111_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__and2b_1
XFILLER_202_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24110_ systolic_inst.B_shift\[1\]\[5\] _11332_ net83 systolic_inst.B_shift\[5\]\[5\]
+ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__a22o_1
XFILLER_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21322_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[4\]\[11\]
+ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__nand2_1
XFILLER_163_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25090_ net113 ser_C.shift_reg\[373\] VGND VGND VPWR VPWR _11015_ sky130_fd_sc_hd__and2_1
XFILLER_163_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_68_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24041_ systolic_inst.B_shift\[4\]\[0\] B_in\[0\] _00008_ VGND VGND VPWR VPWR _10538_
+ sky130_fd_sc_hd__mux2_1
XFILLER_102_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21253_ net117 systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[4\]\[0\]
+ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__a21oi_1
XFILLER_190_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap150 net152 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_16
XFILLER_209_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20204_ _07165_ _07168_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__xor2_1
XFILLER_172_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21184_ _07988_ _08018_ _08017_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__a21boi_2
XFILLER_172_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27800_ clknet_leaf_45_clk _01598_ net137 VGND VGND VPWR VPWR systolic_inst.B_outs\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_20135_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[18\]
+ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__nand2_1
XFILLER_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28780_ clknet_leaf_230_clk _02578_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[328\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25992_ systolic_inst.acc_wires\[14\]\[20\] ser_C.parallel_data\[468\] net25 VGND
+ VGND VPWR VPWR _03294_ sky130_fd_sc_hd__mux2_1
XFILLER_217_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27731_ clknet_leaf_143_clk _01529_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_213_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20066_ _07049_ _07050_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__and2_1
X_24943_ C_out\[298\] net103 net76 ser_C.shift_reg\[298\] _10941_ VGND VGND VPWR VPWR
+ _02548_ sky130_fd_sc_hd__a221o_1
XFILLER_97_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27662_ clknet_leaf_202_clk _01460_ net147 VGND VGND VPWR VPWR systolic_inst.A_outs\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_24874_ net110 ser_C.shift_reg\[265\] VGND VGND VPWR VPWR _10907_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_77_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29401_ clknet_leaf_238_clk _03199_ net146 VGND VGND VPWR VPWR C_out\[373\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26613_ clknet_leaf_17_B_in_serial_clk _00416_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23825_ systolic_inst.acc_wires\[0\]\[16\] systolic_inst.acc_wires\[0\]\[17\] systolic_inst.acc_wires\[0\]\[18\]
+ systolic_inst.acc_wires\[0\]\[19\] systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _10422_ sky130_fd_sc_hd__o41a_1
XFILLER_205_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27593_ clknet_leaf_224_clk _01391_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29332_ clknet_leaf_220_clk _03130_ net140 VGND VGND VPWR VPWR C_out\[304\] sky130_fd_sc_hd__dfrtp_1
X_23756_ _10361_ _10362_ VGND VGND VPWR VPWR _10363_ sky130_fd_sc_hd__and2_1
XFILLER_54_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26544_ clknet_leaf_19_A_in_serial_clk _00347_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ _07836_ _07840_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22707_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[2\]
+ systolic_inst.A_outs\[1\]\[3\] VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__nand4_2
XFILLER_18_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29263_ clknet_leaf_192_clk _03061_ net146 VGND VGND VPWR VPWR C_out\[235\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23687_ _10284_ _10290_ _10292_ _10295_ VGND VGND VPWR VPWR _10305_ sky130_fd_sc_hd__a22o_1
X_26475_ clknet_leaf_15_A_in_serial_clk _00278_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20899_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[2\] systolic_inst.B_outs\[4\]\[3\]
+ systolic_inst.B_outs\[4\]\[4\] VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__and4_1
XFILLER_158_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28214_ clknet_leaf_72_clk _02012_ VGND VGND VPWR VPWR systolic_inst.B_shift\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13440_ deser_A.shift_reg\[4\] deser_A.shift_reg\[5\] deser_A.receiving VGND VGND
+ VPWR VPWR _00277_ sky130_fd_sc_hd__mux2_1
X_22638_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[26\]
+ VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__nand2_1
X_25426_ _11182_ systolic_inst.A_shift\[0\]\[4\] net70 VGND VGND VPWR VPWR _02790_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_230_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29194_ clknet_leaf_215_clk _02992_ net149 VGND VGND VPWR VPWR C_out\[166\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_230_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28145_ clknet_leaf_98_clk _01943_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25357_ ser_C.parallel_data\[505\] net98 net78 ser_C.shift_reg\[505\] _11148_ VGND
+ VGND VPWR VPWR _02755_ sky130_fd_sc_hd__a221o_1
X_13371_ A_in\[80\] deser_A.word_buffer\[80\] net94 VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__mux2_1
XFILLER_107_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22569_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[15\]
+ VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__nor2_1
XFILLER_210_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15110_ _12193_ _12196_ _12225_ VGND VGND VPWR VPWR _12227_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16090_ _13055_ _13058_ _13060_ VGND VGND VPWR VPWR _13085_ sky130_fd_sc_hd__a21oi_1
X_24308_ _10627_ systolic_inst.A_shift\[10\]\[1\] net71 VGND VGND VPWR VPWR _02227_
+ sky130_fd_sc_hd__mux2_1
X_28076_ clknet_leaf_101_clk _01874_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_25288_ net111 ser_C.shift_reg\[472\] VGND VGND VPWR VPWR _11114_ sky130_fd_sc_hd__and2_1
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15041_ _12143_ _12159_ VGND VGND VPWR VPWR _12160_ sky130_fd_sc_hd__xor2_1
XFILLER_68_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27027_ clknet_leaf_11_B_in_serial_clk _00825_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24239_ systolic_inst.A_shift\[19\]\[3\] A_in\[67\] net59 VGND VGND VPWR VPWR _10605_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18800_ net115 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[8\]\[0\]
+ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__a21oi_1
X_19780_ _06752_ _06754_ _06753_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__o21bai_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28978_ clknet_leaf_20_clk _02776_ VGND VGND VPWR VPWR systolic_inst.A_shift\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16992_ net69 _04299_ _04301_ systolic_inst.acc_wires\[11\]\[3\] net105 VGND VGND
+ VPWR VPWR _01237_ sky130_fd_sc_hd__a32o_1
XFILLER_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_196_Right_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18731_ _05855_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__inv_2
X_27929_ clknet_leaf_134_clk _01727_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_118_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15943_ _12963_ VGND VGND VPWR VPWR _12964_ sky130_fd_sc_hd__inv_2
XFILLER_49_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18662_ _05732_ _05788_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__nand2_1
XFILLER_236_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15874_ systolic_inst.acc_wires\[13\]\[16\] systolic_inst.acc_wires\[13\]\[17\] systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12906_ sky130_fd_sc_hd__o21a_1
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_237_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_237_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17613_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[10\]\[6\]
+ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__nand2_1
XFILLER_236_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14825_ _11941_ _11949_ VGND VGND VPWR VPWR _11950_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_237_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18593_ _05691_ _05720_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__xor2_1
XFILLER_92_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ net105 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[13\] _04794_
+ _04795_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__a22o_1
X_14756_ net118 systolic_inst.B_outs\[14\]\[0\] systolic_inst.A_outs\[14\]\[0\] VGND
+ VGND VPWR VPWR _11886_ sky130_fd_sc_hd__and3_1
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_A_in_serial_clk clknet_2_0__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_29_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_232_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13707_ B_in\[14\] deser_B.word_buffer\[14\] net84 VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__mux2_1
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17475_ _04674_ _04692_ _04691_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__o21a_1
XFILLER_189_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14687_ net69 _11840_ _11841_ systolic_inst.acc_wires\[15\]\[23\] net105 VGND VGND
+ VPWR VPWR _01001_ sky130_fd_sc_hd__a32o_1
XFILLER_149_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19214_ systolic_inst.B_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[5\] systolic_inst.A_outs\[7\]\[6\]
+ systolic_inst.B_outs\[7\]\[3\] VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__a22oi_1
XFILLER_34_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16426_ net67 _03791_ _03793_ systolic_inst.acc_wires\[12\]\[9\] net108 VGND VGND
+ VPWR VPWR _01179_ sky130_fd_sc_hd__a32o_1
X_13638_ deser_B.word_buffer\[74\] deser_B.serial_word\[74\] net123 VGND VGND VPWR
+ VPWR _00475_ sky130_fd_sc_hd__mux2_1
XFILLER_20_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19145_ _06209_ _06210_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__or2_1
X_16357_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[14\] _03733_
+ _03735_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__a22o_1
XFILLER_9_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13569_ deser_B.word_buffer\[5\] deser_B.serial_word\[5\] net124 VGND VGND VPWR VPWR
+ _00406_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15308_ systolic_inst.acc_wires\[14\]\[20\] systolic_inst.acc_wires\[14\]\[21\] systolic_inst.acc_wires\[14\]\[22\]
+ systolic_inst.acc_wires\[14\]\[23\] systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12398_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_184_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19076_ _06133_ _06136_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_184_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16288_ _03666_ _03667_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18027_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[9\] _05218_ net116
+ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__mux2_1
X_15239_ net67 _12336_ _12339_ systolic_inst.acc_wires\[14\]\[13\] net107 VGND VGND
+ VPWR VPWR _01055_ sky130_fd_sc_hd__a32o_1
XFILLER_172_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19978_ _06972_ _06973_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__and2b_1
XFILLER_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18929_ net66 _06030_ _06031_ systolic_inst.acc_wires\[8\]\[18\] net108 VGND VGND
+ VPWR VPWR _01444_ sky130_fd_sc_hd__a32o_1
XFILLER_101_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21940_ _08718_ _08724_ _08728_ net60 VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__a31oi_1
XFILLER_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21871_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[3\]\[1\]
+ VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__nand2_1
XFILLER_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23610_ _10229_ _10230_ VGND VGND VPWR VPWR _10231_ sky130_fd_sc_hd__nor2_1
X_20822_ net68 _07719_ _07720_ systolic_inst.acc_wires\[5\]\[30\] net106 VGND VGND
+ VPWR VPWR _01648_ sky130_fd_sc_hd__a32o_1
XFILLER_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_951 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24590_ net114 ser_C.shift_reg\[123\] VGND VGND VPWR VPWR _10765_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23541_ _10158_ _10163_ VGND VGND VPWR VPWR _10164_ sky130_fd_sc_hd__nor2_1
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20753_ _07642_ _07647_ _07652_ _07656_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__or4_1
XFILLER_168_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26260_ clknet_leaf_5_A_in_serial_clk _00068_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_196_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23472_ _10030_ _10032_ _10094_ _10095_ VGND VGND VPWR VPWR _10097_ sky130_fd_sc_hd__a211o_1
X_20684_ _07601_ _07602_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__and2_1
XFILLER_51_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25211_ C_out\[432\] net101 net73 ser_C.shift_reg\[432\] _11075_ VGND VGND VPWR VPWR
+ _02682_ sky130_fd_sc_hd__a221o_1
X_22423_ _09096_ _09161_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__or2_1
X_26191_ _11254_ _11255_ ser_C.bit_idx\[7\] VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__mux2_1
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25142_ net110 ser_C.shift_reg\[399\] VGND VGND VPWR VPWR _11041_ sky130_fd_sc_hd__and2_1
XFILLER_104_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22354_ _09025_ _09095_ VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__xnor2_4
X_21305_ _08155_ _08157_ _08161_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__nand3_1
XFILLER_237_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25073_ C_out\[363\] net97 net77 ser_C.shift_reg\[363\] _11006_ VGND VGND VPWR VPWR
+ _02613_ sky130_fd_sc_hd__a221o_1
X_22285_ _09025_ _09028_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24024_ systolic_inst.B_shift\[6\]\[7\] net70 net83 systolic_inst.B_shift\[10\]\[7\]
+ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__a22o_1
X_28901_ clknet_leaf_273_clk _02699_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_113_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21236_ _08073_ _08102_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28832_ clknet_leaf_195_clk _02630_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21167_ _08002_ _08004_ _08035_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__o21ai_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20118_ _07086_ _07091_ _07095_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28763_ clknet_leaf_214_clk _02561_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[311\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21098_ _07967_ _07968_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__and2_1
X_25975_ systolic_inst.acc_wires\[14\]\[3\] ser_C.parallel_data\[451\] net24 VGND
+ VGND VPWR VPWR _03277_ sky130_fd_sc_hd__mux2_1
XFILLER_213_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27714_ clknet_leaf_189_clk _01512_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_218_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20049_ _07036_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__inv_2
XFILLER_4_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24926_ net111 ser_C.shift_reg\[291\] VGND VGND VPWR VPWR _10933_ sky130_fd_sc_hd__and2_1
XFILLER_111_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28694_ clknet_leaf_193_clk _02492_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[242\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27645_ clknet_leaf_313_clk _01443_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_24857_ C_out\[255\] net99 net79 ser_C.shift_reg\[255\] _10898_ VGND VGND VPWR VPWR
+ _02505_ sky130_fd_sc_hd__a221o_1
XFILLER_74_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14610_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[15\]\[12\]
+ VGND VGND VPWR VPWR _11776_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23808_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[16\]
+ _10404_ VGND VGND VPWR VPWR _10408_ sky130_fd_sc_hd__a21oi_1
XFILLER_215_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15590_ _12644_ _12645_ VGND VGND VPWR VPWR _12646_ sky130_fd_sc_hd__or2_1
XFILLER_92_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27576_ clknet_leaf_221_clk _01374_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_232_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24788_ net113 ser_C.shift_reg\[222\] VGND VGND VPWR VPWR _10864_ sky130_fd_sc_hd__and2_1
XFILLER_2_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_232_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29315_ clknet_leaf_301_clk _03113_ net141 VGND VGND VPWR VPWR C_out\[287\] sky130_fd_sc_hd__dfrtp_1
XFILLER_199_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14541_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[15\]\[0\]
+ _11709_ _11707_ VGND VGND VPWR VPWR _11717_ sky130_fd_sc_hd__a31o_1
X_26527_ clknet_leaf_5_A_in_serial_clk _00330_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23739_ _10346_ _10347_ _10348_ VGND VGND VPWR VPWR _10349_ sky130_fd_sc_hd__a21o_1
XFILLER_144_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29246_ clknet_leaf_187_clk _03044_ net146 VGND VGND VPWR VPWR C_out\[218\] sky130_fd_sc_hd__dfrtp_1
XFILLER_144_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17260_ _04512_ _04518_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__xor2_1
XFILLER_92_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14472_ _11650_ _11651_ VGND VGND VPWR VPWR _11653_ sky130_fd_sc_hd__nor2_1
X_26458_ clknet_leaf_11_clk _00265_ net132 VGND VGND VPWR VPWR A_in\[126\] sky130_fd_sc_hd__dfrtp_1
XFILLER_202_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16211_ systolic_inst.B_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[7\]
+ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__and3_1
X_25409_ systolic_inst.A_shift\[2\]\[4\] A_in\[12\] net59 VGND VGND VPWR VPWR _11174_
+ sky130_fd_sc_hd__mux2_1
X_13423_ deser_A.bit_idx\[1\] _11308_ _11310_ VGND VGND VPWR VPWR _11311_ sky130_fd_sc_hd__o21ai_1
X_29177_ clknet_leaf_137_clk _02975_ net142 VGND VGND VPWR VPWR C_out\[149\] sky130_fd_sc_hd__dfrtp_1
X_17191_ systolic_inst.B_outs\[9\]\[5\] systolic_inst.B_outs\[5\]\[5\] net116 VGND
+ VGND VPWR VPWR _01279_ sky130_fd_sc_hd__mux2_1
XFILLER_220_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26389_ clknet_leaf_17_clk _00196_ net134 VGND VGND VPWR VPWR A_in\[57\] sky130_fd_sc_hd__dfrtp_1
XFILLER_220_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload109 clknet_leaf_284_clk VGND VGND VPWR VPWR clkload109/Y sky130_fd_sc_hd__inv_6
X_28128_ clknet_leaf_124_clk _01926_ net153 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_16142_ systolic_inst.A_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[5\] VGND VGND
+ VPWR VPWR _03527_ sky130_fd_sc_hd__nand2_1
X_13354_ A_in\[63\] deser_A.word_buffer\[63\] net95 VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__mux2_1
XFILLER_155_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28059_ clknet_leaf_98_clk _01857_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_16073_ systolic_inst.A_outs\[12\]\[1\] systolic_inst.B_outs\[12\]\[6\] VGND VGND
+ VPWR VPWR _13069_ sky130_fd_sc_hd__nand2_1
X_13285_ deser_A.word_buffer\[123\] deser_A.serial_word\[123\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_226_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19901_ _06897_ _06898_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__nor2_1
X_15024_ _12141_ _12142_ VGND VGND VPWR VPWR _12143_ sky130_fd_sc_hd__nand2_1
XFILLER_69_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19832_ systolic_inst.A_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[6\] _11278_ systolic_inst.A_outs\[6\]\[2\]
+ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_36_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_239_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19763_ _06729_ _06764_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_239_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16975_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[11\]\[0\]
+ _04285_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__and4_1
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18714_ systolic_inst.B_outs\[8\]\[5\] systolic_inst.A_outs\[8\]\[7\] VGND VGND VPWR
+ VPWR _05839_ sky130_fd_sc_hd__nand2_1
XFILLER_232_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15926_ systolic_inst.acc_wires\[13\]\[24\] systolic_inst.acc_wires\[13\]\[25\] systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12950_ sky130_fd_sc_hd__o21a_1
XFILLER_77_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19694_ _06694_ _06697_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_177_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18645_ systolic_inst.A_outs\[8\]\[3\] systolic_inst.A_outs\[8\]\[4\] systolic_inst.B_outs\[8\]\[6\]
+ systolic_inst.B_outs\[8\]\[7\] VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__and4b_1
X_15857_ _12891_ _12890_ systolic_inst.acc_wires\[13\]\[15\] net108 VGND VGND VPWR
+ VPWR _01121_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_237_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14808_ _11900_ _11921_ _11923_ VGND VGND VPWR VPWR _11933_ sky130_fd_sc_hd__a21oi_1
X_18576_ systolic_inst.A_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[5\] VGND VGND VPWR
+ VPWR _05705_ sky130_fd_sc_hd__nand2_1
XFILLER_91_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15788_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[13\]\[6\]
+ VGND VGND VPWR VPWR _12832_ sky130_fd_sc_hd__nand2_1
X_17527_ _04714_ _04778_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__nand2_1
X_14739_ _11885_ _11884_ systolic_inst.acc_wires\[15\]\[31\] net105 VGND VGND VPWR
+ VPWR _01009_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17458_ systolic_inst.B_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\] VGND VGND
+ VPWR VPWR _04712_ sky130_fd_sc_hd__or2_1
XFILLER_178_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16409_ net67 _03777_ _03779_ systolic_inst.acc_wires\[12\]\[6\] net108 VGND VGND
+ VPWR VPWR _01176_ sky130_fd_sc_hd__a32o_1
XFILLER_203_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17389_ systolic_inst.B_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[5\]
+ systolic_inst.A_outs\[10\]\[6\] VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__and4_1
X_19128_ _06192_ _06193_ _06161_ _06163_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__o211a_1
XFILLER_199_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_232_Right_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_294_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_294_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_238_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19059_ _06126_ _06127_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__nand2_1
XFILLER_12_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22070_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[30\]
+ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__or2_1
XFILLER_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21021_ _07892_ _07893_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__and2_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22972_ _09614_ _09619_ VGND VGND VPWR VPWR _09650_ sky130_fd_sc_hd__nand2_1
X_25760_ systolic_inst.acc_wires\[7\]\[12\] C_out\[236\] net42 VGND VGND VPWR VPWR
+ _03062_ sky130_fd_sc_hd__mux2_1
XFILLER_142_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24711_ C_out\[182\] net99 net79 ser_C.shift_reg\[182\] _10825_ VGND VGND VPWR VPWR
+ _02432_ sky130_fd_sc_hd__a221o_1
X_21923_ _08713_ _08714_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__nor2_1
XFILLER_83_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25691_ systolic_inst.acc_wires\[5\]\[7\] C_out\[167\] net16 VGND VGND VPWR VPWR
+ _02993_ sky130_fd_sc_hd__mux2_1
XFILLER_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27430_ clknet_leaf_242_clk _01228_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_21854_ _08654_ _08655_ VGND VGND VPWR VPWR _08657_ sky130_fd_sc_hd__xnor2_1
X_24642_ net7 ser_C.shift_reg\[149\] VGND VGND VPWR VPWR _10791_ sky130_fd_sc_hd__and2_1
XFILLER_83_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20805_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[28\]
+ VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__or2_1
XFILLER_145_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27361_ clknet_leaf_322_clk _01159_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24573_ C_out\[113\] net100 net80 ser_C.shift_reg\[113\] _10756_ VGND VGND VPWR VPWR
+ _02363_ sky130_fd_sc_hd__a221o_1
X_21785_ systolic_inst.B_outs\[3\]\[5\] systolic_inst.A_outs\[3\]\[7\] VGND VGND VPWR
+ VPWR _08590_ sky130_fd_sc_hd__nand2_1
XFILLER_51_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29100_ clknet_leaf_154_clk _02898_ net150 VGND VGND VPWR VPWR C_out\[72\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_20__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_20__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_169_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26312_ clknet_leaf_27_A_in_serial_clk _00120_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_20736_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[16\]
+ _07644_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__a21oi_1
X_23524_ _10145_ _10146_ VGND VGND VPWR VPWR _10147_ sky130_fd_sc_hd__or2_1
X_27292_ clknet_leaf_291_clk _01090_ net141 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29031_ clknet_leaf_126_clk _02829_ net144 VGND VGND VPWR VPWR C_out\[3\] sky130_fd_sc_hd__dfrtp_1
X_23455_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[7\]
+ VGND VGND VPWR VPWR _10080_ sky130_fd_sc_hd__and3_2
XFILLER_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26243_ clknet_leaf_17_A_in_serial_clk _00051_ net143 VGND VGND VPWR VPWR deser_A.word_buffer\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_20667_ _07586_ _07587_ _07588_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__nand3_1
XFILLER_137_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22406_ _09056_ _09114_ _09112_ VGND VGND VPWR VPWR _09147_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_115_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26174_ net7 ser_C.bit_idx\[0\] ser_C.bit_idx\[1\] VGND VGND VPWR VPWR _11245_ sky130_fd_sc_hd__and3_1
X_23386_ _09997_ _10011_ VGND VGND VPWR VPWR _10013_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_115_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20598_ _07499_ _07502_ _07527_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_115_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_285_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_285_clk
+ sky130_fd_sc_hd__clkbuf_8
X_22337_ _09077_ _09078_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__xnor2_1
X_25125_ C_out\[389\] net101 net73 ser_C.shift_reg\[389\] _11032_ VGND VGND VPWR VPWR
+ _02639_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25056_ net112 ser_C.shift_reg\[356\] VGND VGND VPWR VPWR _10998_ sky130_fd_sc_hd__and2_1
X_22268_ _08981_ _09011_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__xor2_1
XFILLER_140_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24007_ systolic_inst.B_shift\[9\]\[7\] B_in\[15\] _00008_ VGND VGND VPWR VPWR _10529_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21219_ _08085_ _08086_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22199_ _08915_ _08938_ _08937_ VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_221_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_221_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28815_ clknet_leaf_240_clk _02613_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[363\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28746_ clknet_leaf_298_clk _02544_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[294\]
+ sky130_fd_sc_hd__dfrtp_1
X_16760_ _04080_ _04079_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__nand2b_1
X_13972_ deser_B.shift_reg\[6\] deser_B.shift_reg\[7\] net125 VGND VGND VPWR VPWR
+ _00798_ sky130_fd_sc_hd__mux2_1
X_25958_ systolic_inst.acc_wires\[13\]\[18\] C_out\[434\] net20 VGND VGND VPWR VPWR
+ _03260_ sky130_fd_sc_hd__mux2_1
XFILLER_4_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15711_ _12762_ _12763_ VGND VGND VPWR VPWR _12764_ sky130_fd_sc_hd__nor2_1
XFILLER_58_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24909_ C_out\[281\] net103 net75 ser_C.shift_reg\[281\] _10924_ VGND VGND VPWR VPWR
+ _02531_ sky130_fd_sc_hd__a221o_1
X_28677_ clknet_leaf_197_clk _02475_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[225\]
+ sky130_fd_sc_hd__dfrtp_1
X_16691_ _04011_ _04012_ _03980_ _03982_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__o211a_1
XFILLER_46_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25889_ systolic_inst.acc_wires\[11\]\[13\] C_out\[365\] net40 VGND VGND VPWR VPWR
+ _03191_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18430_ _05557_ _05563_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15642_ _12687_ _12695_ VGND VGND VPWR VPWR _12697_ sky130_fd_sc_hd__xnor2_1
X_27628_ clknet_leaf_323_clk _01426_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_234_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18361_ _05521_ _05520_ systolic_inst.acc_wires\[9\]\[24\] net106 VGND VGND VPWR
+ VPWR _01386_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_29_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15573_ _12586_ _12594_ _12593_ VGND VGND VPWR VPWR _12630_ sky130_fd_sc_hd__a21o_1
X_27559_ clknet_leaf_305_clk _01357_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17312_ _04568_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__and2_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14524_ _11699_ _11702_ VGND VGND VPWR VPWR _11703_ sky130_fd_sc_hd__xnor2_1
X_18292_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[15\]
+ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__nor2_1
XFILLER_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29229_ clknet_leaf_203_clk _03027_ net147 VGND VGND VPWR VPWR C_out\[201\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17243_ net107 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[4\] _04501_
+ _04503_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__a22o_1
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14455_ _11636_ _11635_ VGND VGND VPWR VPWR _11637_ sky130_fd_sc_hd__nand2b_1
XFILLER_70_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13406_ A_in\[115\] deser_A.word_buffer\[115\] _00003_ VGND VGND VPWR VPWR _00254_
+ sky130_fd_sc_hd__mux2_1
X_17174_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[31\]
+ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14386_ _11527_ _11536_ _11535_ VGND VGND VPWR VPWR _11570_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_210_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_210_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16125_ _13079_ _13082_ _03509_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_276_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_276_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_227_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13337_ A_in\[46\] deser_A.word_buffer\[46\] net93 VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16056_ _13020_ _13023_ _13051_ VGND VGND VPWR VPWR _13053_ sky130_fd_sc_hd__or3_1
XFILLER_142_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13268_ deser_A.word_buffer\[106\] deser_A.serial_word\[106\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__mux2_1
XFILLER_124_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_23_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15007_ _12074_ _12091_ _12089_ VGND VGND VPWR VPWR _12127_ sky130_fd_sc_hd__o21a_1
X_13199_ deser_A.word_buffer\[37\] deser_A.serial_word\[37\] net127 VGND VGND VPWR
+ VPWR _00047_ sky130_fd_sc_hd__mux2_1
XFILLER_111_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19815_ _06774_ _06777_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__nor2_1
XFILLER_116_1057 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19746_ _06743_ _06747_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__nor2_1
X_16958_ _04224_ _04225_ _04250_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__a31o_1
XFILLER_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15909_ _12914_ _12921_ _12926_ _12931_ VGND VGND VPWR VPWR _12935_ sky130_fd_sc_hd__nand4_1
X_19677_ _06661_ _06680_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__nand2_1
X_16889_ _04170_ _04172_ _04171_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_200_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_200_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18628_ _05730_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18559_ _05621_ _05622_ _05653_ _05651_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__a31o_1
XFILLER_162_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21570_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[4\] VGND VGND VPWR
+ VPWR _08381_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_155_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_12 systolic_inst.B_shift\[3\]\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1058 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_23 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20521_ _07417_ _07419_ _07454_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__nand3_1
XFILLER_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_34 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_45 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23240_ net65 _09886_ _09887_ systolic_inst.acc_wires\[1\]\[25\] net109 VGND VGND
+ VPWR VPWR _01899_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_151_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20452_ _07348_ _07350_ _07386_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__nand3_1
XFILLER_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_267_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_267_clk
+ sky130_fd_sc_hd__clkbuf_8
X_23171_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[15\]
+ VGND VGND VPWR VPWR _09829_ sky130_fd_sc_hd__and2_1
X_20383_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.A_outs\[5\]\[7\] _07289_ _07288_
+ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_41_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22122_ net109 _08869_ _08870_ _08871_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_164_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22053_ systolic_inst.acc_wires\[3\]\[26\] systolic_inst.acc_wires\[3\]\[27\] systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__o21a_1
XFILLER_121_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26930_ clknet_leaf_3_A_in_serial_clk _00728_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21004_ _07837_ _07876_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__nor2_1
X_26861_ clknet_leaf_1_B_in_serial_clk _00663_ net135 VGND VGND VPWR VPWR deser_B.bit_idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28600_ clknet_leaf_138_clk _02398_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[148\]
+ sky130_fd_sc_hd__dfrtp_1
X_25812_ systolic_inst.acc_wires\[9\]\[0\] C_out\[288\] net14 VGND VGND VPWR VPWR
+ _03114_ sky130_fd_sc_hd__mux2_1
X_29580_ clknet_leaf_25_B_in_serial_clk _03375_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_214_1181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26792_ clknet_leaf_72_clk _00594_ net153 VGND VGND VPWR VPWR B_in\[64\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28531_ clknet_leaf_162_clk _02329_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25743_ systolic_inst.acc_wires\[6\]\[27\] C_out\[219\] net43 VGND VGND VPWR VPWR
+ _03045_ sky130_fd_sc_hd__mux2_1
Xmax_cap14 net15 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_8
X_22955_ _09593_ _09595_ _09594_ VGND VGND VPWR VPWR _09633_ sky130_fd_sc_hd__o21ba_1
XFILLER_90_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap25 net26 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_50_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap36 net54 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_8
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21906_ _08700_ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__inv_2
X_28462_ clknet_leaf_122_clk _02260_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25674_ systolic_inst.acc_wires\[4\]\[22\] C_out\[150\] net32 VGND VGND VPWR VPWR
+ _02976_ sky130_fd_sc_hd__mux2_1
Xmax_cap69 _11712_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_12
XFILLER_83_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22886_ _09562_ _09565_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27413_ clknet_leaf_213_clk _01211_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_65_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24625_ C_out\[139\] net103 net75 ser_C.shift_reg\[139\] _10782_ VGND VGND VPWR VPWR
+ _02389_ sky130_fd_sc_hd__a221o_1
XFILLER_19_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21837_ _11274_ systolic_inst.A_outs\[3\]\[7\] _08590_ _08615_ VGND VGND VPWR VPWR
+ _08640_ sky130_fd_sc_hd__o211ai_1
X_28393_ clknet_leaf_32_clk _02191_ VGND VGND VPWR VPWR systolic_inst.A_shift\[17\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27344_ clknet_leaf_343_clk _01142_ net131 VGND VGND VPWR VPWR systolic_inst.A_outs\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_62_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24556_ net113 ser_C.shift_reg\[106\] VGND VGND VPWR VPWR _10748_ sky130_fd_sc_hd__and2_1
XFILLER_200_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21768_ _08515_ _08573_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20719_ net64 _07632_ _07633_ systolic_inst.acc_wires\[5\]\[14\] net109 VGND VGND
+ VPWR VPWR _01632_ sky130_fd_sc_hd__a32o_1
X_23507_ _10084_ _10086_ _10129_ VGND VGND VPWR VPWR _10131_ sky130_fd_sc_hd__and3_1
XFILLER_141_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27275_ clknet_leaf_271_clk _01073_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24487_ C_out\[70\] _11302_ net81 ser_C.shift_reg\[70\] _10713_ VGND VGND VPWR VPWR
+ _02320_ sky130_fd_sc_hd__a221o_1
X_21699_ _08468_ _08470_ _08506_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29014_ clknet_leaf_93_clk _02812_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26226_ clknet_leaf_8_A_in_serial_clk _00034_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14240_ _11403_ _11425_ _11427_ VGND VGND VPWR VPWR _11428_ sky130_fd_sc_hd__and3_1
X_23438_ _10063_ _10061_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[7\]
+ _11258_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_172_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_258_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_258_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14171_ _11359_ _11360_ VGND VGND VPWR VPWR _11361_ sky130_fd_sc_hd__nor2_1
X_26157_ deser_B.serial_word\[112\] deser_B.shift_reg\[112\] _00001_ VGND VGND VPWR
+ VPWR _03459_ sky130_fd_sc_hd__mux2_1
X_23369_ _09966_ _09994_ VGND VGND VPWR VPWR _09996_ sky130_fd_sc_hd__or2_1
XFILLER_125_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_223_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13122_ systolic_inst.B_outs\[6\]\[7\] VGND VGND VPWR VPWR _11278_ sky130_fd_sc_hd__inv_2
X_25108_ net112 ser_C.shift_reg\[382\] VGND VGND VPWR VPWR _11024_ sky130_fd_sc_hd__and2_1
X_26088_ deser_B.serial_word\[43\] deser_B.shift_reg\[43\] net55 VGND VGND VPWR VPWR
+ _03390_ sky130_fd_sc_hd__mux2_1
XFILLER_113_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17930_ systolic_inst.A_outs\[9\]\[2\] systolic_inst.B_outs\[9\]\[5\] VGND VGND VPWR
+ VPWR _05124_ sky130_fd_sc_hd__nand2_1
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25039_ C_out\[346\] net97 net77 ser_C.shift_reg\[346\] _10989_ VGND VGND VPWR VPWR
+ _02596_ sky130_fd_sc_hd__a221o_1
XFILLER_26_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17861_ _05036_ _05056_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__nand2_1
XFILLER_61_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19600_ systolic_inst.acc_wires\[7\]\[28\] systolic_inst.acc_wires\[7\]\[29\] systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_1388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16812_ systolic_inst.B_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[6\] systolic_inst.A_outs\[11\]\[7\]
+ systolic_inst.B_outs\[11\]\[3\] VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__a22o_1
XFILLER_66_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17792_ systolic_inst.A_outs\[9\]\[7\] systolic_inst.A_outs\[8\]\[7\] net117 VGND
+ VGND VPWR VPWR _01337_ sky130_fd_sc_hd__mux2_1
XFILLER_94_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19531_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[19\]
+ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_50_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28729_ clknet_leaf_326_clk _02527_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[277\]
+ sky130_fd_sc_hd__dfrtp_1
X_16743_ _04062_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__nor2_1
XFILLER_98_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13955_ deser_A.serial_word\[116\] deser_A.shift_reg\[116\] _00002_ VGND VGND VPWR
+ VPWR _00781_ sky130_fd_sc_hd__mux2_1
XFILLER_98_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19462_ _06501_ _06509_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__or2_1
XFILLER_228_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16674_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[4\] _03995_ _03996_
+ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__nand4_2
XFILLER_98_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13886_ deser_A.serial_word\[47\] deser_A.shift_reg\[47\] net58 VGND VGND VPWR VPWR
+ _00712_ sky130_fd_sc_hd__mux2_1
XFILLER_234_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18413_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.B_outs\[3\]\[2\] net119 VGND
+ VGND VPWR VPWR _01404_ sky130_fd_sc_hd__mux2_1
X_15625_ net115 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[11\] VGND
+ VGND VPWR VPWR _12680_ sky130_fd_sc_hd__or2_1
X_19393_ _06448_ _06450_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_191_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _05505_ _05506_ _05504_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15556_ _12577_ _12612_ VGND VGND VPWR VPWR _12613_ sky130_fd_sc_hd__nor2_1
XFILLER_43_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_212_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _11622_ _11664_ _11663_ VGND VGND VPWR VPWR _11687_ sky130_fd_sc_hd__o21ba_1
XFILLER_30_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18275_ _05446_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15487_ _12510_ _12545_ VGND VGND VPWR VPWR _12546_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17226_ systolic_inst.A_outs\[10\]\[1\] systolic_inst.B_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\]
+ systolic_inst.A_outs\[10\]\[0\] VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__a22o_1
X_14438_ _11517_ _11618_ VGND VGND VPWR VPWR _11620_ sky130_fd_sc_hd__and2_2
XFILLER_128_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_249_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_249_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_190_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17157_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[28\]
+ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__nand2_1
X_14369_ _11447_ _11524_ _11525_ VGND VGND VPWR VPWR _11553_ sky130_fd_sc_hd__o21ba_1
XFILLER_183_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16108_ _13069_ _03492_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17088_ _04381_ _04383_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16039_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[3\] VGND VGND
+ VPWR VPWR _13036_ sky130_fd_sc_hd__nand2_1
XFILLER_233_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19729_ _06719_ _06731_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22740_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[4\]
+ systolic_inst.A_outs\[1\]\[5\] VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_0_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22671_ _09370_ _09374_ _09375_ net60 VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__a31o_1
XFILLER_53_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24410_ net114 ser_C.shift_reg\[33\] VGND VGND VPWR VPWR _10675_ sky130_fd_sc_hd__and2_1
X_21622_ _08429_ _08430_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_153_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25390_ _11164_ systolic_inst.A_shift\[2\]\[2\] net71 VGND VGND VPWR VPWR _02772_
+ sky130_fd_sc_hd__mux2_1
XFILLER_200_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21553_ _08336_ _08364_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__nand2_1
XFILLER_21_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24341_ systolic_inst.A_shift\[8\]\[4\] net70 net83 systolic_inst.A_shift\[9\]\[4\]
+ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__a22o_1
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20504_ systolic_inst.A_outs\[5\]\[5\] systolic_inst.B_outs\[5\]\[6\] _11276_ systolic_inst.A_outs\[5\]\[4\]
+ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__o2bb2a_1
X_24272_ systolic_inst.B_shift\[17\]\[7\] net72 _11333_ B_in\[111\] VGND VGND VPWR
+ VPWR _02209_ sky130_fd_sc_hd__a22o_1
X_27060_ clknet_leaf_4_B_in_serial_clk _00858_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21484_ systolic_inst.A_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[1\]
+ systolic_inst.B_outs\[3\]\[0\] VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__a22o_1
XFILLER_165_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23223_ _09872_ VGND VGND VPWR VPWR _09873_ sky130_fd_sc_hd__inv_2
XFILLER_181_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26011_ systolic_inst.acc_wires\[15\]\[7\] ser_C.parallel_data\[487\] net37 VGND
+ VGND VPWR VPWR _03313_ sky130_fd_sc_hd__mux2_1
X_20435_ systolic_inst.A_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[6\] _11276_ systolic_inst.A_outs\[5\]\[2\]
+ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23154_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[1\]\[13\]
+ VGND VGND VPWR VPWR _09814_ sky130_fd_sc_hd__xor2_1
XFILLER_180_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload270 clknet_leaf_141_clk VGND VGND VPWR VPWR clkload270/X sky130_fd_sc_hd__clkbuf_8
X_20366_ _07300_ _07303_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__nand2_1
Xclkload281 clknet_leaf_183_clk VGND VGND VPWR VPWR clkload281/Y sky130_fd_sc_hd__clkinv_8
XFILLER_161_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload292 clknet_leaf_199_clk VGND VGND VPWR VPWR clkload292/Y sky130_fd_sc_hd__clkinv_8
X_22105_ _08848_ _08854_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23085_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[1\]\[3\]
+ VGND VGND VPWR VPWR _09755_ sky130_fd_sc_hd__nand2_1
X_27962_ clknet_leaf_149_clk _01760_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_20297_ systolic_inst.A_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[2\] systolic_inst.B_outs\[5\]\[3\]
+ systolic_inst.B_outs\[5\]\[4\] VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__and4_1
X_22036_ _08807_ _08809_ _08811_ VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__or3_1
X_26913_ clknet_leaf_11_A_in_serial_clk _00711_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27893_ clknet_leaf_39_clk _01691_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_212_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29632_ clknet_leaf_11_B_in_serial_clk _03427_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_26844_ clknet_leaf_74_clk _00646_ net153 VGND VGND VPWR VPWR B_in\[116\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29563_ clknet_leaf_15_B_in_serial_clk _03358_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26775_ clknet_leaf_80_clk _00577_ net153 VGND VGND VPWR VPWR B_in\[47\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23987_ systolic_inst.B_shift\[12\]\[5\] B_in\[69\] _00008_ VGND VGND VPWR VPWR _10519_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28514_ clknet_leaf_158_clk _02312_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_216_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13740_ B_in\[47\] deser_B.word_buffer\[47\] net84 VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__mux2_1
X_25726_ systolic_inst.acc_wires\[6\]\[10\] C_out\[202\] net47 VGND VGND VPWR VPWR
+ _03028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22938_ _09581_ _09583_ VGND VGND VPWR VPWR _09617_ sky130_fd_sc_hd__nand2_1
X_29494_ clknet_leaf_282_clk _03292_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28445_ clknet_leaf_36_clk _02243_ VGND VGND VPWR VPWR systolic_inst.A_shift\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_232_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13671_ deser_B.word_buffer\[107\] deser_B.serial_word\[107\] net123 VGND VGND VPWR
+ VPWR _00508_ sky130_fd_sc_hd__mux2_1
X_25657_ systolic_inst.acc_wires\[4\]\[5\] C_out\[133\] net29 VGND VGND VPWR VPWR
+ _02959_ sky130_fd_sc_hd__mux2_1
X_22869_ _09547_ _09548_ VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__nand2b_1
XFILLER_186_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15410_ _12468_ _12470_ _12451_ VGND VGND VPWR VPWR _12472_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24608_ net110 ser_C.shift_reg\[132\] VGND VGND VPWR VPWR _10774_ sky130_fd_sc_hd__and2_1
X_16390_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__inv_2
X_28376_ clknet_leaf_32_clk _02174_ VGND VGND VPWR VPWR systolic_inst.A_shift\[19\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_25588_ systolic_inst.acc_wires\[2\]\[0\] C_out\[64\] net34 VGND VGND VPWR VPWR _02890_
+ sky130_fd_sc_hd__mux2_1
XFILLER_197_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15341_ _12419_ _12422_ _12421_ VGND VGND VPWR VPWR _12426_ sky130_fd_sc_hd__o21a_1
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27327_ clknet_leaf_331_clk _01125_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_24539_ C_out\[96\] net99 net79 ser_C.shift_reg\[96\] _10739_ VGND VGND VPWR VPWR
+ _02346_ sky130_fd_sc_hd__a221o_1
XFILLER_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18060_ _05180_ _05183_ _05213_ _05214_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__a31o_1
X_15272_ _12358_ _12360_ _12367_ VGND VGND VPWR VPWR _12368_ sky130_fd_sc_hd__a21oi_1
X_27258_ clknet_leaf_280_clk _01056_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17011_ _04314_ _04315_ _04316_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__and3_1
X_26209_ clknet_leaf_14_A_in_serial_clk _00017_ net143 VGND VGND VPWR VPWR deser_A.word_buffer\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14223_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[3\] systolic_inst.A_outs\[15\]\[3\]
+ systolic_inst.B_outs\[15\]\[4\] VGND VGND VPWR VPWR _11411_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_97_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27189_ clknet_leaf_255_clk _00987_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_208_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14154_ net118 _11344_ _11345_ _11338_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__a31o_1
XFILLER_193_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13105_ systolic_inst.B_outs\[7\]\[7\] VGND VGND VPWR VPWR _11261_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14085_ deser_B.shift_reg\[119\] deser_B.shift_reg\[120\] deser_B.receiving VGND
+ VGND VPWR VPWR _00911_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18962_ _06012_ _06013_ _06038_ _06058_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__a211o_1
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17913_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[6\] _05105_
+ _05107_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18893_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[8\]\[14\]
+ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__or2_1
XFILLER_234_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17844_ _05034_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17775_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[30\]
+ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__nand2_1
XFILLER_226_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14987_ _12105_ _12106_ VGND VGND VPWR VPWR _12107_ sky130_fd_sc_hd__or2_1
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19514_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[16\]
+ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__xnor2_1
X_16726_ _04018_ _04046_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_193_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13938_ deser_A.serial_word\[99\] deser_A.shift_reg\[99\] net57 VGND VGND VPWR VPWR
+ _00764_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19445_ _06495_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__inv_2
XFILLER_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16657_ _03956_ _03979_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__xor2_1
X_13869_ deser_A.serial_word\[30\] deser_A.shift_reg\[30\] _00002_ VGND VGND VPWR
+ VPWR _00695_ sky130_fd_sc_hd__mux2_1
XFILLER_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15608_ _12661_ _12662_ VGND VGND VPWR VPWR _12664_ sky130_fd_sc_hd__xor2_1
X_19376_ _06348_ _06433_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__nand2_1
XFILLER_50_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16588_ systolic_inst.B_outs\[10\]\[5\] systolic_inst.B_outs\[6\]\[5\] net120 VGND
+ VGND VPWR VPWR _01215_ sky130_fd_sc_hd__mux2_1
XFILLER_241_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18327_ _05470_ _05471_ _05476_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__and3_1
XFILLER_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15539_ _12596_ _12595_ VGND VGND VPWR VPWR _12597_ sky130_fd_sc_hd__and2b_1
XFILLER_202_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18258_ _05424_ _05428_ _05431_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__nand3_1
XFILLER_147_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17209_ _04469_ _04470_ net120 VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__o21a_1
X_18189_ net116 _05364_ _05374_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__and3_1
XFILLER_11_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_208_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20220_ _07176_ _07180_ _07181_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__a21oi_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20151_ _07120_ _07122_ _07123_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__or3_1
XFILLER_131_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20082_ net106 systolic_inst.acc_wires\[6\]\[10\] net68 _07064_ VGND VGND VPWR VPWR
+ _01564_ sky130_fd_sc_hd__a22o_1
XFILLER_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23910_ systolic_inst.B_shift\[17\]\[7\] B_in\[79\] _00008_ VGND VGND VPWR VPWR _10488_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24890_ net110 ser_C.shift_reg\[273\] VGND VGND VPWR VPWR _10915_ sky130_fd_sc_hd__and2_1
XFILLER_97_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23841_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[23\]
+ VGND VGND VPWR VPWR _10435_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26560_ clknet_leaf_1_A_in_serial_clk _00363_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23772_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[0\]\[12\]
+ VGND VGND VPWR VPWR _10377_ sky130_fd_sc_hd__xnor2_1
X_20984_ _07848_ _07857_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__xnor2_1
XFILLER_232_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25511_ systolic_inst.cycle_cnt\[27\] systolic_inst.cycle_cnt\[26\] _11233_ _11236_
+ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__a31oi_1
XFILLER_225_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22723_ systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[3\] systolic_inst.A_outs\[1\]\[4\]
+ systolic_inst.B_outs\[1\]\[0\] VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26491_ clknet_leaf_8_A_in_serial_clk _00294_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28230_ clknet_leaf_48_clk _02028_ VGND VGND VPWR VPWR systolic_inst.B_shift\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25442_ systolic_inst.cycle_cnt\[3\] _11279_ VGND VGND VPWR VPWR _11192_ sky130_fd_sc_hd__nand2_1
XFILLER_240_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22654_ _09359_ _09362_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__xor2_1
XFILLER_94_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28161_ clknet_leaf_108_clk _01959_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_21605_ systolic_inst.A_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[4\]
+ systolic_inst.B_outs\[3\]\[3\] VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__a22oi_1
XFILLER_240_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22585_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[16\]
+ _09301_ VGND VGND VPWR VPWR _09305_ sky130_fd_sc_hd__a21oi_1
X_25373_ systolic_inst.B_shift\[18\]\[2\] B_in\[50\] net59 VGND VGND VPWR VPWR _11156_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_1223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27112_ clknet_leaf_30_B_in_serial_clk _00910_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24324_ _10635_ systolic_inst.A_shift\[9\]\[1\] net70 VGND VGND VPWR VPWR _02235_
+ sky130_fd_sc_hd__mux2_1
X_28092_ clknet_leaf_111_clk _01890_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_21536_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[4\]
+ systolic_inst.A_outs\[3\]\[5\] VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__and4_1
XFILLER_142_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27043_ clknet_leaf_20_B_in_serial_clk _00841_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_21467_ systolic_inst.A_outs\[3\]\[3\] systolic_inst.A_outs\[2\]\[3\] net122 VGND
+ VGND VPWR VPWR _01717_ sky130_fd_sc_hd__mux2_1
XFILLER_154_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24255_ systolic_inst.A_shift\[17\]\[6\] net70 net83 systolic_inst.A_shift\[18\]\[6\]
+ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__a22o_1
XFILLER_193_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_177_Right_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23206_ _09855_ _09857_ _09858_ VGND VGND VPWR VPWR _09859_ sky130_fd_sc_hd__or3_1
X_20418_ _07315_ _07317_ _07314_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__a21oi_1
XFILLER_175_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21398_ _08232_ _08239_ _08240_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__a21oi_1
X_24186_ systolic_inst.A_shift\[24\]\[1\] net70 _10505_ systolic_inst.A_shift\[25\]\[1\]
+ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__a22o_1
XFILLER_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23137_ net109 systolic_inst.acc_wires\[1\]\[10\] net64 _09799_ VGND VGND VPWR VPWR
+ _01884_ sky130_fd_sc_hd__a22o_1
XFILLER_175_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20349_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[6\] VGND VGND VPWR
+ VPWR _07287_ sky130_fd_sc_hd__nand2_1
XFILLER_134_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28994_ clknet_leaf_47_clk _02792_ VGND VGND VPWR VPWR systolic_inst.A_shift\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_241_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23068_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[1\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _09741_ sky130_fd_sc_hd__a21o_1
X_27945_ clknet_leaf_148_clk _01743_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22019_ _08789_ _08790_ _08797_ VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14910_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] _12031_ VGND
+ VGND VPWR VPWR _12032_ sky130_fd_sc_hd__a21o_1
XFILLER_62_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15890_ net67 _12918_ _12919_ systolic_inst.acc_wires\[13\]\[20\] net108 VGND VGND
+ VPWR VPWR _01126_ sky130_fd_sc_hd__a32o_1
X_27876_ clknet_leaf_38_clk _01674_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26827_ clknet_leaf_86_clk _00629_ net135 VGND VGND VPWR VPWR B_in\[99\] sky130_fd_sc_hd__dfrtp_1
X_29615_ clknet_leaf_1_B_in_serial_clk _03410_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_14841_ _11961_ _11964_ VGND VGND VPWR VPWR _11965_ sky130_fd_sc_hd__xor2_1
XFILLER_124_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29546_ clknet_leaf_250_clk _03341_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_95_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17560_ _04740_ _04788_ _04787_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__o21ba_1
X_26758_ clknet_leaf_75_clk _00560_ net143 VGND VGND VPWR VPWR B_in\[30\] sky130_fd_sc_hd__dfrtp_1
X_14772_ systolic_inst.A_outs\[14\]\[1\] systolic_inst.B_outs\[14\]\[2\] systolic_inst.B_outs\[14\]\[3\]
+ systolic_inst.A_outs\[14\]\[0\] VGND VGND VPWR VPWR _11899_ sky130_fd_sc_hd__a22oi_1
XFILLER_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16511_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[21\]
+ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__xor2_1
XFILLER_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25709_ systolic_inst.acc_wires\[5\]\[25\] C_out\[185\] net45 VGND VGND VPWR VPWR
+ _03011_ sky130_fd_sc_hd__mux2_1
X_13723_ B_in\[30\] deser_B.word_buffer\[30\] net85 VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__mux2_1
X_29477_ clknet_leaf_273_clk _03275_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[449\]
+ sky130_fd_sc_hd__dfrtp_1
X_17491_ systolic_inst.A_outs\[10\]\[5\] systolic_inst.B_outs\[10\]\[6\] systolic_inst.A_outs\[10\]\[6\]
+ systolic_inst.B_outs\[10\]\[7\] VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__and4b_1
X_26689_ clknet_leaf_30_B_in_serial_clk _00492_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19230_ _06276_ _06293_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__xor2_1
XFILLER_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28428_ clknet_leaf_24_clk _02226_ VGND VGND VPWR VPWR systolic_inst.A_shift\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16442_ _03797_ _03806_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__and2_1
X_13654_ deser_B.word_buffer\[90\] deser_B.serial_word\[90\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__mux2_1
XFILLER_143_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19161_ _06224_ _06225_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28359_ clknet_leaf_74_clk _02157_ VGND VGND VPWR VPWR systolic_inst.B_shift\[22\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16373_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[12\]\[0\]
+ _03744_ _03746_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13585_ deser_B.word_buffer\[21\] deser_B.serial_word\[21\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__mux2_1
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18112_ _05262_ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__xnor2_1
X_15324_ _12403_ _12405_ _12411_ VGND VGND VPWR VPWR _12412_ sky130_fd_sc_hd__a21o_1
X_19092_ _06150_ _06158_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__xor2_1
XFILLER_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18043_ _05231_ _05232_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__xnor2_1
X_15255_ _12329_ _12337_ _12351_ _12352_ VGND VGND VPWR VPWR _12353_ sky130_fd_sc_hd__o31a_1
XFILLER_173_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14206_ _11385_ _11394_ VGND VGND VPWR VPWR _11395_ sky130_fd_sc_hd__nor2_1
XFILLER_193_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15186_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[14\]\[6\]
+ VGND VGND VPWR VPWR _12294_ sky130_fd_sc_hd__or2_1
XFILLER_158_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14137_ systolic_inst.B_outs\[14\]\[5\] systolic_inst.B_outs\[10\]\[5\] net120 VGND
+ VGND VPWR VPWR _00959_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19994_ _06988_ _06987_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__and2b_1
XFILLER_140_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_203_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14068_ deser_B.shift_reg\[102\] deser_B.shift_reg\[103\] net126 VGND VGND VPWR VPWR
+ _00894_ sky130_fd_sc_hd__mux2_1
X_18945_ _06036_ _06042_ _06043_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__a21oi_1
XFILLER_234_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18876_ _05962_ _05966_ _05967_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17827_ _05017_ _05023_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17758_ _04978_ _04979_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16709_ _04027_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__xnor2_1
X_17689_ _04919_ _04920_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__nor2_1
XFILLER_39_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_1__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_139_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19428_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[7\]\[4\]
+ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__or2_1
XFILLER_62_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19359_ _06376_ _06418_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22370_ _09111_ _09110_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_171_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21321_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[4\]\[11\]
+ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__or2_1
XFILLER_198_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24040_ _10537_ systolic_inst.B_shift\[4\]\[7\] net72 VGND VGND VPWR VPWR _02049_
+ sky130_fd_sc_hd__mux2_1
X_21252_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[4\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap140 net141 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_16
Xmax_cap151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_16
X_20203_ _07166_ _07167_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__nand2_1
XFILLER_172_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21183_ _08026_ _08050_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__xor2_1
XFILLER_176_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20134_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[18\]
+ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__or2_1
XFILLER_137_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25991_ systolic_inst.acc_wires\[14\]\[19\] ser_C.parallel_data\[467\] net25 VGND
+ VGND VPWR VPWR _03293_ sky130_fd_sc_hd__mux2_1
XFILLER_48_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27730_ clknet_leaf_142_clk _01528_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_20065_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[6\]\[8\]
+ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__xor2_1
X_24942_ net111 ser_C.shift_reg\[299\] VGND VGND VPWR VPWR _10941_ sky130_fd_sc_hd__and2_1
XFILLER_225_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27661_ clknet_leaf_202_clk _01459_ net147 VGND VGND VPWR VPWR systolic_inst.A_outs\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_24873_ C_out\[263\] net101 net73 ser_C.shift_reg\[263\] _10906_ VGND VGND VPWR VPWR
+ _02513_ sky130_fd_sc_hd__a221o_1
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29400_ clknet_leaf_239_clk _03198_ net145 VGND VGND VPWR VPWR C_out\[372\] sky130_fd_sc_hd__dfrtp_1
X_26612_ clknet_leaf_16_B_in_serial_clk _00415_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_23824_ _10401_ _10420_ VGND VGND VPWR VPWR _10421_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27592_ clknet_leaf_224_clk _01390_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29331_ clknet_leaf_219_clk _03129_ net140 VGND VGND VPWR VPWR C_out\[303\] sky130_fd_sc_hd__dfrtp_1
X_26543_ clknet_leaf_20_A_in_serial_clk _00346_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_23755_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[0\]\[10\]
+ VGND VGND VPWR VPWR _10362_ sky130_fd_sc_hd__or2_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20967_ _07840_ _07836_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__nand2b_1
XFILLER_214_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22706_ _09390_ _09391_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__nor2_1
X_29262_ clknet_leaf_192_clk _03060_ net146 VGND VGND VPWR VPWR C_out\[234\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26474_ clknet_leaf_15_A_in_serial_clk _00277_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23686_ systolic_inst.ce_local _10303_ _10304_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_81_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ systolic_inst.A_outs\[4\]\[2\] systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\]
+ systolic_inst.A_outs\[4\]\[1\] VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__a22oi_1
XFILLER_198_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28213_ clknet_leaf_72_clk _02011_ VGND VGND VPWR VPWR systolic_inst.B_shift\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25425_ systolic_inst.A_shift\[1\]\[4\] A_in\[4\] net59 VGND VGND VPWR VPWR _11182_
+ sky130_fd_sc_hd__mux2_1
X_22637_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[26\]
+ VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__or2_1
X_29193_ clknet_leaf_217_clk _02991_ net149 VGND VGND VPWR VPWR C_out\[165\] sky130_fd_sc_hd__dfrtp_1
XFILLER_224_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_230_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_230_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_A_in_serial_clk clknet_2_3__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_16_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_28144_ clknet_leaf_122_clk _01942_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25356_ net112 ser_C.shift_reg\[506\] VGND VGND VPWR VPWR _11148_ sky130_fd_sc_hd__and2_1
X_13370_ A_in\[79\] deser_A.word_buffer\[79\] net94 VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__mux2_1
XFILLER_224_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22568_ net65 _09289_ _09290_ systolic_inst.acc_wires\[2\]\[14\] net109 VGND VGND
+ VPWR VPWR _01824_ sky130_fd_sc_hd__a32o_1
XFILLER_221_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24307_ systolic_inst.A_shift\[11\]\[1\] A_in\[41\] net59 VGND VGND VPWR VPWR _10627_
+ sky130_fd_sc_hd__mux2_1
X_28075_ clknet_leaf_151_clk _01873_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_186_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21519_ _08313_ _08330_ _08331_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__a21oi_1
XFILLER_166_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25287_ ser_C.parallel_data\[470\] net102 net74 ser_C.shift_reg\[470\] _11113_ VGND
+ VGND VPWR VPWR _02720_ sky130_fd_sc_hd__a221o_1
X_22499_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[2\]\[5\]
+ VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__nand2_1
X_27026_ clknet_leaf_19_B_in_serial_clk _00824_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_15040_ _12157_ _12158_ VGND VGND VPWR VPWR _12159_ sky130_fd_sc_hd__nand2_1
XFILLER_170_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24238_ _10604_ systolic_inst.A_shift\[18\]\[2\] net70 VGND VGND VPWR VPWR _02180_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24169_ systolic_inst.A_shift\[26\]\[0\] net70 net83 systolic_inst.A_shift\[27\]\[0\]
+ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__a22o_1
XFILLER_150_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16991_ _04300_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__inv_2
XFILLER_150_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28977_ clknet_leaf_19_clk _02775_ VGND VGND VPWR VPWR systolic_inst.A_shift\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15942_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[29\]
+ VGND VGND VPWR VPWR _12963_ sky130_fd_sc_hd__xor2_1
XFILLER_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18730_ _05853_ _05854_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__or2_1
X_27928_ clknet_leaf_134_clk _01726_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_62_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _05785_ _05786_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__xnor2_1
X_15873_ _12903_ _12904_ VGND VGND VPWR VPWR _12905_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27859_ clknet_leaf_36_clk _01657_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_97_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_237_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14824_ _11942_ _11947_ VGND VGND VPWR VPWR _11949_ sky130_fd_sc_hd__xor2_1
X_17612_ _11712_ _04853_ _04855_ systolic_inst.acc_wires\[10\]\[5\] net105 VGND VGND
+ VPWR VPWR _01303_ sky130_fd_sc_hd__a32o_1
XFILLER_76_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_237_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18592_ _05720_ _05691_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_237_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17543_ _04763_ _04768_ _04793_ net118 VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__o31a_1
X_29529_ clknet_leaf_262_clk _03327_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[501\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ systolic_inst.B_outs\[13\]\[7\] systolic_inst.B_outs\[9\]\[7\] net115 VGND
+ VGND VPWR VPWR _01025_ sky130_fd_sc_hd__mux2_1
XFILLER_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13706_ B_in\[13\] deser_B.word_buffer\[13\] net84 VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__mux2_1
XFILLER_72_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17474_ _04711_ _04727_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__xor2_1
XFILLER_220_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_213_Right_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14686_ _11832_ _11836_ _11839_ VGND VGND VPWR VPWR _11841_ sky130_fd_sc_hd__a21o_1
XFILLER_232_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19213_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[7\] VGND VGND VPWR
+ VPWR _06277_ sky130_fd_sc_hd__nand2_4
X_16425_ _03786_ _03790_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__a21oi_1
X_13637_ deser_B.word_buffer\[73\] deser_B.serial_word\[73\] net123 VGND VGND VPWR
+ VPWR _00474_ sky130_fd_sc_hd__mux2_1
XFILLER_220_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19144_ systolic_inst.A_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[4\]
+ systolic_inst.B_outs\[7\]\[3\] VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__a22oi_1
XFILLER_125_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16356_ net108 _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__nor2_1
X_13568_ deser_B.word_buffer\[4\] deser_B.serial_word\[4\] net124 VGND VGND VPWR VPWR
+ _00405_ sky130_fd_sc_hd__mux2_1
XFILLER_34_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15307_ _12353_ _12354_ _12376_ _12396_ VGND VGND VPWR VPWR _12397_ sky130_fd_sc_hd__a211o_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_229_Left_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19075_ net105 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[4\] _06143_
+ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__a21bo_1
XFILLER_12_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16287_ _03667_ _03666_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_184_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13499_ deser_A.shift_reg\[63\] deser_A.shift_reg\[64\] net129 VGND VGND VPWR VPWR
+ _00336_ sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18026_ _05216_ _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__xnor2_1
X_15238_ _12333_ _12335_ _12338_ VGND VGND VPWR VPWR _12339_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15169_ _11712_ _12277_ _12279_ systolic_inst.acc_wires\[14\]\[3\] net107 VGND VGND
+ VPWR VPWR _01045_ sky130_fd_sc_hd__a32o_1
XFILLER_99_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19977_ _06939_ _06941_ _06971_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__o21ai_1
XFILLER_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18928_ _06027_ _06028_ _06029_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__nand3_1
XFILLER_80_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_238_Left_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18859_ _05962_ _05964_ _05968_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__a21bo_1
XFILLER_28_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21870_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[3\]\[1\]
+ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__and2_1
XFILLER_242_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20821_ _07715_ _07718_ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__or2_1
XFILLER_82_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23540_ _10161_ _10162_ VGND VGND VPWR VPWR _10163_ sky130_fd_sc_hd__or2_1
X_20752_ _07659_ _07660_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__and2_1
XFILLER_165_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23471_ _10030_ _10032_ _10094_ _10095_ VGND VGND VPWR VPWR _10096_ sky130_fd_sc_hd__a211oi_1
X_20683_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[5\]\[10\]
+ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__or2_1
XFILLER_11_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25210_ net110 ser_C.shift_reg\[433\] VGND VGND VPWR VPWR _11075_ sky130_fd_sc_hd__and2_1
X_22422_ _09096_ _09161_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__nand2_1
XFILLER_149_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26190_ _11252_ _11255_ ser_C.bit_idx\[6\] VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__mux2_1
XFILLER_164_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25141_ C_out\[397\] net101 net73 ser_C.shift_reg\[397\] _11040_ VGND VGND VPWR VPWR
+ _02647_ sky130_fd_sc_hd__a221o_1
X_22353_ _09060_ _09094_ systolic_inst.A_outs\[2\]\[7\] VGND VGND VPWR VPWR _09095_
+ sky130_fd_sc_hd__and3b_1
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21304_ _08159_ _08160_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__nand2_1
X_22284_ _09026_ _09027_ VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__nor2_1
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25072_ net112 ser_C.shift_reg\[364\] VGND VGND VPWR VPWR _11006_ sky130_fd_sc_hd__and2_1
XFILLER_117_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24023_ systolic_inst.B_shift\[6\]\[6\] _11332_ net83 systolic_inst.B_shift\[10\]\[6\]
+ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__a22o_1
X_21235_ _08100_ _08101_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_113_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28900_ clknet_leaf_272_clk _02698_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[448\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28831_ clknet_leaf_194_clk _02629_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[379\]
+ sky130_fd_sc_hd__dfrtp_1
X_21166_ _08033_ _08034_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20117_ _07093_ _07094_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__or2_1
X_28762_ clknet_leaf_214_clk _02560_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21097_ systolic_inst.A_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[6\] _07928_ _07929_
+ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__a31o_1
X_25974_ systolic_inst.acc_wires\[14\]\[2\] ser_C.parallel_data\[450\] net24 VGND
+ VGND VPWR VPWR _03276_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27713_ clknet_leaf_189_clk _01511_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_20048_ _07032_ _07033_ _07034_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__and3_1
X_24925_ C_out\[289\] net102 net74 ser_C.shift_reg\[289\] _10932_ VGND VGND VPWR VPWR
+ _02539_ sky130_fd_sc_hd__a221o_1
XFILLER_213_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28693_ clknet_leaf_194_clk _02491_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[241\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_207_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27644_ clknet_leaf_314_clk _01442_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24856_ net110 ser_C.shift_reg\[256\] VGND VGND VPWR VPWR _10898_ sky130_fd_sc_hd__and2_4
XFILLER_171_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23807_ _10406_ VGND VGND VPWR VPWR _10407_ sky130_fd_sc_hd__inv_2
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27575_ clknet_leaf_305_clk _01373_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_24787_ C_out\[220\] net99 net79 ser_C.shift_reg\[220\] _10863_ VGND VGND VPWR VPWR
+ _02470_ sky130_fd_sc_hd__a221o_1
X_21999_ _08773_ _08777_ _08779_ net60 VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__a31o_1
XFILLER_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_232_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29314_ clknet_leaf_301_clk _03112_ net141 VGND VGND VPWR VPWR C_out\[286\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_232_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14540_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[15\]\[2\]
+ VGND VGND VPWR VPWR _11716_ sky130_fd_sc_hd__or2_1
X_26526_ clknet_leaf_6_A_in_serial_clk _00329_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_215_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23738_ _10341_ _10342_ _10340_ VGND VGND VPWR VPWR _10348_ sky130_fd_sc_hd__a21bo_1
XFILLER_109_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29245_ clknet_leaf_187_clk _03043_ net148 VGND VGND VPWR VPWR C_out\[217\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _11650_ _11651_ VGND VGND VPWR VPWR _11652_ sky130_fd_sc_hd__and2_1
X_26457_ clknet_leaf_10_clk _00264_ net132 VGND VGND VPWR VPWR A_in\[125\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23669_ _10258_ _10287_ _10080_ VGND VGND VPWR VPWR _10288_ sky130_fd_sc_hd__o21ba_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16210_ systolic_inst.B_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[6\] systolic_inst.A_outs\[12\]\[7\]
+ systolic_inst.B_outs\[12\]\[3\] VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__a22o_1
XFILLER_224_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25408_ _11173_ systolic_inst.A_shift\[1\]\[3\] net70 VGND VGND VPWR VPWR _02781_
+ sky130_fd_sc_hd__mux2_1
X_13422_ net130 net1 VGND VGND VPWR VPWR _11310_ sky130_fd_sc_hd__nand2b_1
X_29176_ clknet_leaf_138_clk _02974_ net142 VGND VGND VPWR VPWR C_out\[148\] sky130_fd_sc_hd__dfrtp_1
X_17190_ systolic_inst.B_outs\[9\]\[4\] systolic_inst.B_outs\[5\]\[4\] net116 VGND
+ VGND VPWR VPWR _01278_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26388_ clknet_leaf_17_clk _00195_ net133 VGND VGND VPWR VPWR A_in\[56\] sky130_fd_sc_hd__dfrtp_1
XFILLER_155_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28127_ clknet_leaf_123_clk _01925_ net144 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16141_ _03524_ _03525_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__xnor2_1
X_25339_ ser_C.parallel_data\[496\] net97 net77 ser_C.shift_reg\[496\] _11139_ VGND
+ VGND VPWR VPWR _02746_ sky130_fd_sc_hd__a221o_1
X_13353_ A_in\[62\] deser_A.word_buffer\[62\] net92 VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__mux2_1
XFILLER_194_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28058_ clknet_leaf_98_clk _01856_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16072_ systolic_inst.A_outs\[12\]\[1\] systolic_inst.B_outs\[12\]\[5\] systolic_inst.B_outs\[12\]\[6\]
+ systolic_inst.A_outs\[12\]\[0\] VGND VGND VPWR VPWR _13068_ sky130_fd_sc_hd__a22oi_1
X_13284_ deser_A.word_buffer\[122\] deser_A.serial_word\[122\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__mux2_1
XFILLER_142_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27009_ clknet_leaf_17_B_in_serial_clk _00807_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_19900_ systolic_inst.A_outs\[6\]\[5\] systolic_inst.B_outs\[6\]\[6\] _11278_ systolic_inst.A_outs\[6\]\[4\]
+ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__o2bb2a_1
X_15023_ _12031_ _12140_ VGND VGND VPWR VPWR _12142_ sky130_fd_sc_hd__nand2_1
XFILLER_68_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19831_ systolic_inst.A_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[6\]
+ systolic_inst.B_outs\[6\]\[7\] VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_36_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_239_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19762_ _06756_ _06762_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16974_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[11\]\[1\]
+ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__or2_1
XFILLER_49_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18713_ _05836_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__nor2_1
X_15925_ _12947_ _12948_ VGND VGND VPWR VPWR _12949_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19693_ _06695_ _06696_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_177_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15856_ _12880_ _12885_ _12889_ net61 VGND VGND VPWR VPWR _12891_ sky130_fd_sc_hd__a31o_1
X_18644_ systolic_inst.B_outs\[8\]\[5\] systolic_inst.A_outs\[8\]\[5\] VGND VGND VPWR
+ VPWR _05771_ sky130_fd_sc_hd__nand2_1
XFILLER_225_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14807_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[4\] _11932_
+ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__a21bo_1
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15787_ net67 _12829_ _12831_ systolic_inst.acc_wires\[13\]\[5\] net107 VGND VGND
+ VPWR VPWR _01111_ sky130_fd_sc_hd__a32o_1
X_18575_ _05702_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14738_ _11878_ _11882_ _11883_ net61 VGND VGND VPWR VPWR _11885_ sky130_fd_sc_hd__a31o_1
X_17526_ _04776_ _04777_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__and2_1
XFILLER_166_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17457_ _04709_ _04710_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__nand2_1
XFILLER_221_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14669_ net69 _11825_ _11826_ systolic_inst.acc_wires\[15\]\[20\] net107 VGND VGND
+ VPWR VPWR _00998_ sky130_fd_sc_hd__a32o_1
XFILLER_20_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16408_ _03778_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__inv_2
XFILLER_242_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17388_ systolic_inst.B_outs\[10\]\[4\] systolic_inst.A_outs\[10\]\[5\] systolic_inst.A_outs\[10\]\[6\]
+ systolic_inst.B_outs\[10\]\[3\] VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__a22oi_1
XFILLER_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19127_ _06161_ _06163_ _06192_ _06193_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__a211oi_1
X_16339_ _03632_ _03716_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__nand2_1
XFILLER_203_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19058_ systolic_inst.A_outs\[7\]\[1\] systolic_inst.B_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\]
+ systolic_inst.A_outs\[7\]\[0\] VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__a22o_1
XFILLER_146_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18009_ _05160_ _05162_ _05161_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__o21ba_1
XFILLER_82_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21020_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[6\] _07854_ _07853_
+ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__a31o_1
XFILLER_0_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_162_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_162_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22971_ _09647_ _09648_ VGND VGND VPWR VPWR _09649_ sky130_fd_sc_hd__nand2b_1
X_24710_ net113 ser_C.shift_reg\[183\] VGND VGND VPWR VPWR _10825_ sky130_fd_sc_hd__and2_1
XFILLER_110_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21922_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[3\]\[9\]
+ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__and2_1
XFILLER_132_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25690_ systolic_inst.acc_wires\[5\]\[6\] C_out\[166\] net16 VGND VGND VPWR VPWR
+ _02992_ sky130_fd_sc_hd__mux2_1
XFILLER_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24641_ C_out\[147\] net104 net76 ser_C.shift_reg\[147\] _10790_ VGND VGND VPWR VPWR
+ _02397_ sky130_fd_sc_hd__a221o_1
XFILLER_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21853_ _08655_ _08654_ VGND VGND VPWR VPWR _08656_ sky130_fd_sc_hd__nand2b_1
XFILLER_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20804_ _07689_ _07691_ _07703_ _07704_ _07697_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__a311oi_4
X_27360_ clknet_leaf_327_clk _01158_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24572_ net113 ser_C.shift_reg\[114\] VGND VGND VPWR VPWR _10756_ sky130_fd_sc_hd__and2_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21784_ _08587_ _08588_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__nor2_1
X_26311_ clknet_leaf_28_A_in_serial_clk _00119_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_223_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23523_ systolic_inst.B_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[5\] _10025_ VGND
+ VGND VPWR VPWR _10146_ sky130_fd_sc_hd__a21oi_1
X_20735_ _07646_ VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__inv_2
X_27291_ clknet_leaf_319_clk _01089_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_208_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29030_ clknet_leaf_127_clk _02828_ net144 VGND VGND VPWR VPWR C_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26242_ clknet_leaf_12_A_in_serial_clk _00050_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_23454_ systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[6\] systolic_inst.A_outs\[0\]\[7\]
+ systolic_inst.B_outs\[0\]\[1\] VGND VGND VPWR VPWR _10079_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_119_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20666_ _07581_ _07582_ _07580_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__a21bo_1
XFILLER_91_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22405_ _09091_ _09144_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__xor2_1
X_26173_ net7 _10643_ ser_C.bit_idx\[0\] VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20597_ _07499_ _07502_ _07527_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__a21oi_1
X_23385_ _09997_ _10011_ VGND VGND VPWR VPWR _10012_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25124_ net110 ser_C.shift_reg\[390\] VGND VGND VPWR VPWR _11032_ sky130_fd_sc_hd__and2_1
X_22336_ _09078_ _09077_ VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_76_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25055_ C_out\[354\] net98 net78 ser_C.shift_reg\[354\] _10997_ VGND VGND VPWR VPWR
+ _02604_ sky130_fd_sc_hd__a221o_1
X_22267_ _09011_ _08981_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_72_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24006_ _10528_ systolic_inst.B_shift\[5\]\[6\] _11332_ VGND VGND VPWR VPWR _02024_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21218_ _08052_ _08053_ _08057_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__o21ba_1
X_22198_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[6\] _08944_ net122
+ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__mux2_1
XFILLER_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_221_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_221_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28814_ clknet_leaf_243_clk _02612_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[362\]
+ sky130_fd_sc_hd__dfrtp_1
X_21149_ _07988_ _08018_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13971_ deser_B.shift_reg\[5\] deser_B.shift_reg\[6\] net125 VGND VGND VPWR VPWR
+ _00797_ sky130_fd_sc_hd__mux2_1
X_25957_ systolic_inst.acc_wires\[13\]\[17\] C_out\[433\] net20 VGND VGND VPWR VPWR
+ _03259_ sky130_fd_sc_hd__mux2_1
X_28745_ clknet_leaf_297_clk _02543_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[293\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15710_ _12760_ _12761_ VGND VGND VPWR VPWR _12763_ sky130_fd_sc_hd__and2b_1
XFILLER_46_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24908_ net110 ser_C.shift_reg\[282\] VGND VGND VPWR VPWR _10924_ sky130_fd_sc_hd__and2_1
X_28676_ clknet_leaf_197_clk _02474_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[224\]
+ sky130_fd_sc_hd__dfrtp_1
X_16690_ _03980_ _03982_ _04011_ _04012_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__a211oi_1
X_25888_ systolic_inst.acc_wires\[11\]\[12\] C_out\[364\] net39 VGND VGND VPWR VPWR
+ _03190_ sky130_fd_sc_hd__mux2_1
X_15641_ _12687_ _12695_ VGND VGND VPWR VPWR _12696_ sky130_fd_sc_hd__nand2_1
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24839_ C_out\[246\] net98 net78 ser_C.shift_reg\[246\] _10889_ VGND VGND VPWR VPWR
+ _02496_ sky130_fd_sc_hd__a221o_1
X_27627_ clknet_leaf_317_clk _01425_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18360_ _05514_ _05516_ _05519_ net60 VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__a31o_1
X_15572_ _12620_ _12628_ VGND VGND VPWR VPWR _12629_ sky130_fd_sc_hd__xnor2_1
X_27558_ clknet_leaf_305_clk _01356_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _04566_ _04567_ _04538_ _04540_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__o211ai_1
XFILLER_202_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _11700_ _11701_ VGND VGND VPWR VPWR _11702_ sky130_fd_sc_hd__xnor2_1
X_26509_ clknet_leaf_17_A_in_serial_clk _00312_ net143 VGND VGND VPWR VPWR deser_A.shift_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18291_ net66 _05460_ _05461_ systolic_inst.acc_wires\[9\]\[14\] net107 VGND VGND
+ VPWR VPWR _01376_ sky130_fd_sc_hd__a32o_1
XFILLER_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27489_ clknet_leaf_228_clk _01287_ net140 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ net107 _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__nor2_1
XFILLER_175_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29228_ clknet_leaf_210_clk _03026_ net147 VGND VGND VPWR VPWR C_out\[200\] sky130_fd_sc_hd__dfrtp_1
X_14454_ _11590_ _11607_ _11606_ VGND VGND VPWR VPWR _11636_ sky130_fd_sc_hd__o21a_1
XFILLER_109_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13405_ A_in\[114\] deser_A.word_buffer\[114\] _00003_ VGND VGND VPWR VPWR _00253_
+ sky130_fd_sc_hd__mux2_1
X_17173_ net62 _04454_ _04455_ systolic_inst.acc_wires\[11\]\[30\] net105 VGND VGND
+ VPWR VPWR _01264_ sky130_fd_sc_hd__a32o_1
X_29159_ clknet_leaf_309_clk _02957_ net142 VGND VGND VPWR VPWR C_out\[131\] sky130_fd_sc_hd__dfrtp_1
X_14385_ _11560_ _11568_ VGND VGND VPWR VPWR _11569_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_210_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16124_ _13079_ _13082_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__nor3_1
X_13336_ A_in\[45\] deser_A.word_buffer\[45\] net95 VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__mux2_1
XFILLER_227_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16055_ _13020_ _13023_ VGND VGND VPWR VPWR _13052_ sky130_fd_sc_hd__nor2_1
X_13267_ deser_A.word_buffer\[105\] deser_A.serial_word\[105\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__mux2_1
XFILLER_108_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15006_ _12107_ _12125_ VGND VGND VPWR VPWR _12126_ sky130_fd_sc_hd__xor2_1
XFILLER_68_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13198_ deser_A.word_buffer\[36\] deser_A.serial_word\[36\] net127 VGND VGND VPWR
+ VPWR _00046_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_18_B_in_serial_clk clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_18_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_19814_ _06813_ _06814_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__nor2_1
XFILLER_97_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19745_ _11278_ _06746_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16957_ _04221_ _04248_ _04249_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__o21ai_1
XFILLER_238_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15908_ net67 _12933_ _12934_ systolic_inst.acc_wires\[13\]\[23\] net108 VGND VGND
+ VPWR VPWR _01129_ sky130_fd_sc_hd__a32o_1
X_19676_ _06661_ _06680_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__or2_1
X_16888_ _04203_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18627_ _05752_ _05753_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__xnor2_1
X_15839_ _12867_ _12868_ _12875_ VGND VGND VPWR VPWR _12876_ sky130_fd_sc_hd__a21o_1
XFILLER_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18558_ _05655_ _05686_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17509_ _04672_ _04731_ _04730_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18489_ _05619_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__and2_1
XFILLER_162_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_13 systolic_inst.load_acc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20520_ _07394_ _07453_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__xnor2_1
XANTENNA_24 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_35 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_46 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20451_ _07348_ _07350_ _07386_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__a21o_1
XFILLER_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23170_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[15\]
+ VGND VGND VPWR VPWR _09828_ sky130_fd_sc_hd__nor2_1
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20382_ _07285_ _07291_ _07293_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__a21oi_1
X_22121_ net109 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[3\] VGND
+ VGND VPWR VPWR _08871_ sky130_fd_sc_hd__nand2_1
XFILLER_161_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22052_ _08805_ _08808_ _08821_ _08824_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__or4_1
XFILLER_161_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21003_ systolic_inst.B_outs\[4\]\[4\] systolic_inst.A_outs\[4\]\[5\] VGND VGND VPWR
+ VPWR _07876_ sky130_fd_sc_hd__nand2_1
X_26860_ clknet_leaf_1_B_in_serial_clk _00662_ net135 VGND VGND VPWR VPWR deser_B.bit_idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25811_ systolic_inst.acc_wires\[8\]\[31\] C_out\[287\] net27 VGND VGND VPWR VPWR
+ _03113_ sky130_fd_sc_hd__mux2_1
XFILLER_101_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26791_ clknet_leaf_72_clk _00593_ net153 VGND VGND VPWR VPWR B_in\[63\] sky130_fd_sc_hd__dfrtp_1
X_28530_ clknet_leaf_166_clk _02328_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_214_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25742_ systolic_inst.acc_wires\[6\]\[26\] C_out\[218\] net44 VGND VGND VPWR VPWR
+ _03044_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22954_ _09628_ _09631_ VGND VGND VPWR VPWR _09632_ sky130_fd_sc_hd__xor2_1
XFILLER_233_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap15 net16 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_6
XFILLER_210_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap26 net27 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_8
XFILLER_228_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21905_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[3\]\[6\]
+ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__nand2_1
X_28461_ clknet_leaf_124_clk _02259_ net153 VGND VGND VPWR VPWR ser_C.shift_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap48 net49 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_8
X_25673_ systolic_inst.acc_wires\[4\]\[21\] C_out\[149\] net32 VGND VGND VPWR VPWR
+ _02975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22885_ _09563_ _09564_ VGND VGND VPWR VPWR _09565_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_104_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27412_ clknet_leaf_223_clk _01210_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_24624_ net110 ser_C.shift_reg\[140\] VGND VGND VPWR VPWR _10782_ sky130_fd_sc_hd__and2_1
X_21836_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[13\] _08638_
+ _08639_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28392_ clknet_leaf_32_clk _02190_ VGND VGND VPWR VPWR systolic_inst.A_shift\[17\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27343_ clknet_leaf_342_clk _01141_ net131 VGND VGND VPWR VPWR systolic_inst.A_outs\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24555_ C_out\[104\] net99 net79 ser_C.shift_reg\[104\] _10747_ VGND VGND VPWR VPWR
+ _02354_ sky130_fd_sc_hd__a221o_1
XFILLER_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21767_ _08570_ _08571_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23506_ _10084_ _10086_ _10129_ VGND VGND VPWR VPWR _10130_ sky130_fd_sc_hd__a21oi_2
XFILLER_145_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20718_ _07629_ _07631_ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__or2_1
X_27274_ clknet_leaf_272_clk _01072_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_24486_ net112 ser_C.shift_reg\[71\] VGND VGND VPWR VPWR _10713_ sky130_fd_sc_hd__and2_1
XFILLER_141_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21698_ _08480_ _08505_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29013_ clknet_leaf_93_clk _02811_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26225_ clknet_leaf_8_A_in_serial_clk _00033_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23437_ net121 _10062_ VGND VGND VPWR VPWR _10063_ sky130_fd_sc_hd__nand2_1
X_20649_ net64 _07571_ _07573_ systolic_inst.acc_wires\[5\]\[4\] net109 VGND VGND
+ VPWR VPWR _01622_ sky130_fd_sc_hd__a32o_1
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_227_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26156_ deser_B.serial_word\[111\] deser_B.shift_reg\[111\] _00001_ VGND VGND VPWR
+ VPWR _03458_ sky130_fd_sc_hd__mux2_1
XFILLER_194_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14170_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[2\]
+ systolic_inst.A_outs\[15\]\[3\] VGND VGND VPWR VPWR _11360_ sky130_fd_sc_hd__and4_1
X_23368_ _09966_ _09994_ VGND VGND VPWR VPWR _09995_ sky130_fd_sc_hd__nand2_1
XFILLER_180_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13121_ systolic_inst.B_outs\[1\]\[7\] VGND VGND VPWR VPWR _11277_ sky130_fd_sc_hd__inv_2
X_25107_ C_out\[380\] net99 net79 ser_C.shift_reg\[380\] _11023_ VGND VGND VPWR VPWR
+ _02630_ sky130_fd_sc_hd__a221o_1
XFILLER_30_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_223_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22319_ _09025_ _09061_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__xor2_1
X_26087_ deser_B.serial_word\[42\] deser_B.shift_reg\[42\] net55 VGND VGND VPWR VPWR
+ _03389_ sky130_fd_sc_hd__mux2_1
X_23299_ systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[3\] VGND VGND VPWR
+ VPWR _09929_ sky130_fd_sc_hd__nand2_1
XFILLER_124_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25038_ net112 ser_C.shift_reg\[347\] VGND VGND VPWR VPWR _10989_ sky130_fd_sc_hd__and2_1
XFILLER_152_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17860_ _05051_ _05054_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16811_ _04128_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__or2_1
XFILLER_8_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17791_ systolic_inst.A_outs\[9\]\[6\] systolic_inst.A_outs\[8\]\[6\] net117 VGND
+ VGND VPWR VPWR _01336_ sky130_fd_sc_hd__mux2_1
X_26989_ clknet_leaf_30_A_in_serial_clk _00787_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19530_ net105 systolic_inst.acc_wires\[7\]\[18\] net62 _06568_ VGND VGND VPWR VPWR
+ _01508_ sky130_fd_sc_hd__a22o_1
XFILLER_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13954_ deser_A.serial_word\[115\] deser_A.shift_reg\[115\] _00002_ VGND VGND VPWR
+ VPWR _00780_ sky130_fd_sc_hd__mux2_1
X_28728_ clknet_leaf_325_clk _02526_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[276\]
+ sky130_fd_sc_hd__dfrtp_1
X_16742_ systolic_inst.B_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[5\]
+ systolic_inst.B_outs\[11\]\[3\] VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_50_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19461_ _06505_ _06507_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__nand2_1
X_16673_ systolic_inst.B_outs\[11\]\[3\] systolic_inst.A_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\]
+ systolic_inst.A_outs\[11\]\[2\] VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__a22o_1
XFILLER_185_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28659_ clknet_leaf_182_clk _02457_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[207\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_194_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_194_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13885_ deser_A.serial_word\[46\] deser_A.shift_reg\[46\] net58 VGND VGND VPWR VPWR
+ _00711_ sky130_fd_sc_hd__mux2_1
XFILLER_234_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18412_ systolic_inst.B_outs\[7\]\[1\] systolic_inst.B_outs\[3\]\[1\] net119 VGND
+ VGND VPWR VPWR _01403_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15624_ net115 _12677_ _12678_ _12679_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__a31o_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19392_ _06448_ _06450_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__nand2_1
XFILLER_185_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_191_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18343_ _05497_ _05498_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15555_ _12583_ _12585_ _12582_ VGND VGND VPWR VPWR _12612_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_191_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_212_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14506_ _11622_ _11685_ VGND VGND VPWR VPWR _11686_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18274_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[9\]\[12\]
+ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__nand2_1
XFILLER_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15486_ _12539_ _12543_ VGND VGND VPWR VPWR _12545_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14437_ _11517_ _11618_ VGND VGND VPWR VPWR _11619_ sky130_fd_sc_hd__or2_1
X_17225_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[2\] VGND VGND
+ VPWR VPWR _04486_ sky130_fd_sc_hd__nand2_1
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17156_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[28\]
+ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__or2_1
X_14368_ _11515_ _11516_ _11517_ _11521_ VGND VGND VPWR VPWR _11552_ sky130_fd_sc_hd__a31o_1
XFILLER_239_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16107_ systolic_inst.A_outs\[12\]\[1\] systolic_inst.B_outs\[12\]\[6\] _03492_ VGND
+ VGND VPWR VPWR _03493_ sky130_fd_sc_hd__and3_1
X_13319_ A_in\[28\] deser_A.word_buffer\[28\] net91 VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17087_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[16\]
+ _04379_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__a21oi_1
X_14299_ _11483_ _11484_ VGND VGND VPWR VPWR _11485_ sky130_fd_sc_hd__nor2_1
XFILLER_100_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16038_ systolic_inst.A_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[5\] VGND VGND
+ VPWR VPWR _13035_ sky130_fd_sc_hd__nand2_1
XFILLER_135_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_206_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_179_Left_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17989_ _05180_ _05181_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__and2_1
XFILLER_38_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19728_ _06699_ _06730_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19659_ systolic_inst.A_outs\[6\]\[0\] systolic_inst.A_outs\[6\]\[1\] systolic_inst.B_outs\[6\]\[3\]
+ systolic_inst.B_outs\[6\]\[4\] VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_0_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_185_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_185_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_157_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22670_ _09370_ _09374_ _09375_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21621_ _08430_ _08429_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_153_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_188_Left_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24340_ systolic_inst.A_shift\[8\]\[3\] net70 net83 systolic_inst.A_shift\[9\]\[3\]
+ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__a22o_1
X_21552_ _08353_ _08361_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_60_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20503_ systolic_inst.A_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[5\] systolic_inst.B_outs\[5\]\[6\]
+ systolic_inst.B_outs\[5\]\[7\] VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__and4b_1
XFILLER_138_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24271_ systolic_inst.B_shift\[17\]\[6\] net72 _11333_ B_in\[110\] VGND VGND VPWR
+ VPWR _02208_ sky130_fd_sc_hd__a22o_1
X_21483_ _08298_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__inv_2
XFILLER_148_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26010_ systolic_inst.acc_wires\[15\]\[6\] ser_C.parallel_data\[486\] net37 VGND
+ VGND VPWR VPWR _03312_ sky130_fd_sc_hd__mux2_1
XFILLER_88_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23222_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[23\]
+ VGND VGND VPWR VPWR _09872_ sky130_fd_sc_hd__xor2_1
XFILLER_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20434_ systolic_inst.A_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[6\]
+ systolic_inst.B_outs\[5\]\[7\] VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__and4b_1
XFILLER_193_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload260 clknet_leaf_103_clk VGND VGND VPWR VPWR clkload260/Y sky130_fd_sc_hd__bufinv_16
X_23153_ net109 systolic_inst.acc_wires\[1\]\[12\] net64 _09813_ VGND VGND VPWR VPWR
+ _01886_ sky130_fd_sc_hd__a22o_1
XFILLER_146_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20365_ _07301_ _07302_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__nand2_1
XFILLER_88_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload271 clknet_leaf_208_clk VGND VGND VPWR VPWR clkload271/Y sky130_fd_sc_hd__clkinv_2
Xclkload282 clknet_leaf_184_clk VGND VGND VPWR VPWR clkload282/Y sky130_fd_sc_hd__clkinv_2
XFILLER_122_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22104_ _08852_ _08853_ _08848_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__or3b_1
Xclkload293 clknet_leaf_203_clk VGND VGND VPWR VPWR clkload293/Y sky130_fd_sc_hd__inv_6
X_23084_ net64 _09752_ _09754_ systolic_inst.acc_wires\[1\]\[2\] _11258_ VGND VGND
+ VPWR VPWR _01876_ sky130_fd_sc_hd__a32o_1
X_27961_ clknet_leaf_148_clk _01759_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_161_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20296_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[3\] VGND VGND VPWR
+ VPWR _07236_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_197_Left_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22035_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[25\]
+ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__xor2_1
X_26912_ clknet_leaf_18_A_in_serial_clk _00710_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_27892_ clknet_leaf_38_clk _01690_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29631_ clknet_leaf_10_B_in_serial_clk _03426_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26843_ clknet_leaf_74_clk _00645_ net153 VGND VGND VPWR VPWR B_in\[115\] sky130_fd_sc_hd__dfrtp_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29562_ clknet_leaf_15_B_in_serial_clk _03357_ net152 VGND VGND VPWR VPWR deser_B.serial_word\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_26774_ clknet_leaf_96_clk _00576_ net153 VGND VGND VPWR VPWR B_in\[46\] sky130_fd_sc_hd__dfrtp_1
X_23986_ _10518_ systolic_inst.B_shift\[8\]\[4\] net72 VGND VGND VPWR VPWR _02014_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28513_ clknet_leaf_157_clk _02311_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_25725_ systolic_inst.acc_wires\[6\]\[9\] C_out\[201\] net47 VGND VGND VPWR VPWR
+ _03027_ sky130_fd_sc_hd__mux2_1
XFILLER_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22937_ _09614_ _09615_ VGND VGND VPWR VPWR _09616_ sky130_fd_sc_hd__nand2_1
XFILLER_5_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_216_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_176_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_176_clk
+ sky130_fd_sc_hd__clkbuf_8
X_29493_ clknet_leaf_281_clk _03291_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_216_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13670_ deser_B.word_buffer\[106\] deser_B.serial_word\[106\] net123 VGND VGND VPWR
+ VPWR _00507_ sky130_fd_sc_hd__mux2_1
X_28444_ clknet_leaf_25_clk _02242_ VGND VGND VPWR VPWR systolic_inst.A_shift\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25656_ systolic_inst.acc_wires\[4\]\[4\] C_out\[132\] net29 VGND VGND VPWR VPWR
+ _02958_ sky130_fd_sc_hd__mux2_1
XFILLER_231_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22868_ _09548_ _09547_ VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__nand2b_1
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24607_ C_out\[130\] net103 net75 ser_C.shift_reg\[130\] _10773_ VGND VGND VPWR VPWR
+ _02380_ sky130_fd_sc_hd__a221o_1
X_21819_ _08556_ _08622_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__nand2_1
XFILLER_169_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28375_ clknet_leaf_31_clk _02173_ VGND VGND VPWR VPWR systolic_inst.A_shift\[19\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25587_ systolic_inst.acc_wires\[1\]\[31\] C_out\[63\] net34 VGND VGND VPWR VPWR
+ _02889_ sky130_fd_sc_hd__mux2_1
XFILLER_71_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22799_ systolic_inst.B_outs\[1\]\[1\] systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[5\]
+ systolic_inst.A_outs\[1\]\[6\] VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__and4_1
XFILLER_19_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15340_ _12424_ VGND VGND VPWR VPWR _12425_ sky130_fd_sc_hd__inv_2
X_27326_ clknet_leaf_330_clk _01124_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_212_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24538_ net113 ser_C.shift_reg\[97\] VGND VGND VPWR VPWR _10739_ sky130_fd_sc_hd__and2_1
XFILLER_19_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27257_ clknet_leaf_280_clk _01055_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_15271_ systolic_inst.acc_wires\[14\]\[16\] systolic_inst.acc_wires\[14\]\[17\] systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12367_ sky130_fd_sc_hd__o21a_1
XFILLER_40_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24469_ C_out\[61\] net100 net82 ser_C.shift_reg\[61\] _10704_ VGND VGND VPWR VPWR
+ _02311_ sky130_fd_sc_hd__a221o_1
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17010_ _04314_ _04315_ _04316_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__a21o_1
X_26208_ clknet_leaf_15_A_in_serial_clk _00016_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14222_ _11381_ _11409_ VGND VGND VPWR VPWR _11410_ sky130_fd_sc_hd__xor2_1
XFILLER_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27188_ clknet_leaf_254_clk _00986_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26139_ deser_B.serial_word\[94\] deser_B.shift_reg\[94\] net56 VGND VGND VPWR VPWR
+ _03441_ sky130_fd_sc_hd__mux2_1
X_14153_ _11336_ _11343_ VGND VGND VPWR VPWR _11345_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_100_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_193_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13104_ systolic_inst.B_outs\[12\]\[7\] VGND VGND VPWR VPWR _11260_ sky130_fd_sc_hd__inv_2
XFILLER_98_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14084_ deser_B.shift_reg\[118\] deser_B.shift_reg\[119\] deser_B.receiving VGND
+ VGND VPWR VPWR _00910_ sky130_fd_sc_hd__mux2_1
XFILLER_113_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18961_ _06037_ _06044_ _06049_ _06054_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_56_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17912_ net107 _05106_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__nor2_1
XFILLER_191_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18892_ net108 systolic_inst.acc_wires\[8\]\[13\] net63 _05999_ VGND VGND VPWR VPWR
+ _01439_ sky130_fd_sc_hd__a22o_1
XFILLER_224_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17843_ _05019_ _05038_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_7_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_201_Left_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17774_ _04983_ _04986_ _04989_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__o31a_1
X_14986_ _12031_ _12104_ VGND VGND VPWR VPWR _12106_ sky130_fd_sc_hd__and2_1
XFILLER_78_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19513_ _06552_ _06553_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__and2_1
XFILLER_235_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16725_ _04018_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_167_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_167_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13937_ deser_A.serial_word\[98\] deser_A.shift_reg\[98\] net57 VGND VGND VPWR VPWR
+ _00763_ sky130_fd_sc_hd__mux2_1
XFILLER_208_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_193_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19444_ _06485_ _06489_ _06492_ _06493_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__o211a_1
X_13868_ deser_A.serial_word\[29\] deser_A.shift_reg\[29\] _00002_ VGND VGND VPWR
+ VPWR _00694_ sky130_fd_sc_hd__mux2_1
XFILLER_35_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16656_ _03956_ _03979_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__nand2_1
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15607_ _12661_ _12662_ VGND VGND VPWR VPWR _12663_ sky130_fd_sc_hd__nand2b_1
X_19375_ _06348_ _06433_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__or2_1
XFILLER_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13799_ B_in\[106\] deser_B.word_buffer\[106\] net90 VGND VGND VPWR VPWR _00636_
+ sky130_fd_sc_hd__mux2_1
X_16587_ systolic_inst.B_outs\[10\]\[4\] systolic_inst.B_outs\[6\]\[4\] net120 VGND
+ VGND VPWR VPWR _01214_ sky130_fd_sc_hd__mux2_1
XFILLER_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18326_ _05489_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__and2_1
XFILLER_241_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15538_ _12521_ _12556_ _12558_ VGND VGND VPWR VPWR _12596_ sky130_fd_sc_hd__a21oi_1
XFILLER_230_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_210_Left_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15469_ _12497_ _12527_ _12528_ VGND VGND VPWR VPWR _12529_ sky130_fd_sc_hd__and3_1
X_18257_ _05424_ _05428_ _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__a21o_1
XFILLER_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17208_ _04469_ _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__nand2_1
XFILLER_163_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18188_ _05370_ _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__xnor2_1
XFILLER_239_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17139_ _04422_ _04424_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__or3_1
XFILLER_144_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20150_ systolic_inst.acc_wires\[6\]\[16\] systolic_inst.acc_wires\[6\]\[17\] systolic_inst.acc_wires\[6\]\[18\]
+ systolic_inst.acc_wires\[6\]\[19\] systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__o41a_1
XFILLER_235_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20081_ _07061_ _07063_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__xor2_1
XFILLER_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_227_Right_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23840_ net64 _10433_ _10434_ systolic_inst.acc_wires\[0\]\[22\] _11258_ VGND VGND
+ VPWR VPWR _01952_ sky130_fd_sc_hd__a32o_1
XFILLER_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23771_ _10361_ _10367_ _10369_ VGND VGND VPWR VPWR _10376_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_158_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_158_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_101_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20983_ _07817_ _07855_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__xor2_1
X_25510_ systolic_inst.cycle_cnt\[27\] _11279_ _11233_ systolic_inst.cycle_cnt\[26\]
+ VGND VGND VPWR VPWR _11236_ sky130_fd_sc_hd__a22oi_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_A_in_serial_clk clknet_2_1__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_24_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_226_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22722_ _09403_ _09406_ VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__xnor2_1
X_26490_ clknet_leaf_8_A_in_serial_clk _00293_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25441_ systolic_inst.ce_local _11190_ VGND VGND VPWR VPWR _11191_ sky130_fd_sc_hd__and2_1
XFILLER_214_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22653_ _09360_ _09361_ VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__nand2_1
XFILLER_230_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28160_ clknet_leaf_109_clk _01958_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_21604_ systolic_inst.B_outs\[3\]\[3\] systolic_inst.A_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\]
+ systolic_inst.A_outs\[3\]\[4\] VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__and4_1
XFILLER_16_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25372_ _11155_ systolic_inst.B_shift\[14\]\[1\] _11332_ VGND VGND VPWR VPWR _02763_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22584_ _09303_ VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__inv_2
XFILLER_222_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27111_ clknet_leaf_29_B_in_serial_clk _00909_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24323_ systolic_inst.A_shift\[10\]\[1\] A_in\[33\] net59 VGND VGND VPWR VPWR _10635_
+ sky130_fd_sc_hd__mux2_1
X_28091_ clknet_leaf_113_clk _01889_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_193_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21535_ systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[5\]
+ systolic_inst.B_outs\[3\]\[0\] VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__a22oi_1
XFILLER_193_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_330_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_330_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_135_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27042_ clknet_leaf_18_B_in_serial_clk _00840_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_239_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24254_ systolic_inst.A_shift\[17\]\[5\] net70 net83 systolic_inst.A_shift\[18\]\[5\]
+ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__a22o_1
X_21466_ systolic_inst.A_outs\[3\]\[2\] systolic_inst.A_outs\[2\]\[2\] net122 VGND
+ VGND VPWR VPWR _01716_ sky130_fd_sc_hd__mux2_1
XFILLER_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23205_ systolic_inst.acc_wires\[1\]\[16\] systolic_inst.acc_wires\[1\]\[17\] systolic_inst.acc_wires\[1\]\[18\]
+ systolic_inst.acc_wires\[1\]\[19\] systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09858_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_131_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20417_ _07351_ _07352_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_131_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24185_ systolic_inst.A_shift\[24\]\[0\] net70 _10505_ systolic_inst.A_shift\[25\]\[0\]
+ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__a22o_1
X_21397_ _08240_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__inv_2
XFILLER_218_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23136_ _09796_ _09798_ VGND VGND VPWR VPWR _09799_ sky130_fd_sc_hd__xor2_1
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20348_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.A_outs\[5\]\[7\] VGND VGND VPWR
+ VPWR _07286_ sky130_fd_sc_hd__nand2_1
X_28993_ clknet_leaf_36_clk _02791_ VGND VGND VPWR VPWR systolic_inst.A_shift\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_241_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_241_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27944_ clknet_leaf_148_clk _01742_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_23067_ net109 systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] _09734_
+ _09740_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__a22o_1
X_20279_ _07199_ _07217_ _07218_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__nor3_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22018_ systolic_inst.acc_wires\[3\]\[20\] systolic_inst.acc_wires\[3\]\[21\] systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__o21a_1
XFILLER_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27875_ clknet_leaf_38_clk _01673_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29614_ clknet_leaf_1_B_in_serial_clk _03409_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26826_ clknet_leaf_86_clk _00628_ net135 VGND VGND VPWR VPWR B_in\[98\] sky130_fd_sc_hd__dfrtp_1
X_14840_ _11962_ _11963_ VGND VGND VPWR VPWR _11964_ sky130_fd_sc_hd__nor2_1
XFILLER_64_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14771_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[2\] _11897_
+ _11898_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__a22o_1
X_29545_ clknet_leaf_250_clk _03340_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_217_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23969_ systolic_inst.B_shift\[13\]\[4\] B_in\[44\] _00008_ VGND VGND VPWR VPWR _10510_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_149_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_149_clk
+ sky130_fd_sc_hd__clkbuf_8
X_26757_ clknet_leaf_52_clk _00559_ net143 VGND VGND VPWR VPWR B_in\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_229_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13722_ B_in\[29\] deser_B.word_buffer\[29\] net85 VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__mux2_1
X_16510_ net67 _03865_ _03866_ systolic_inst.acc_wires\[12\]\[20\] net108 VGND VGND
+ VPWR VPWR _01190_ sky130_fd_sc_hd__a32o_1
XFILLER_217_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25708_ systolic_inst.acc_wires\[5\]\[24\] C_out\[184\] net45 VGND VGND VPWR VPWR
+ _03010_ sky130_fd_sc_hd__mux2_1
XFILLER_17_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26688_ clknet_leaf_31_B_in_serial_clk _00491_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29476_ clknet_leaf_273_clk _03274_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[448\]
+ sky130_fd_sc_hd__dfrtp_1
X_17490_ systolic_inst.B_outs\[10\]\[6\] systolic_inst.A_outs\[10\]\[6\] _11275_ systolic_inst.A_outs\[10\]\[5\]
+ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_186_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13653_ deser_B.word_buffer\[89\] deser_B.serial_word\[89\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__mux2_1
X_16441_ _03796_ _03801_ _03802_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__and3_1
X_28427_ clknet_leaf_21_clk _02225_ VGND VGND VPWR VPWR systolic_inst.A_shift\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25639_ systolic_inst.acc_wires\[3\]\[19\] C_out\[115\] net50 VGND VGND VPWR VPWR
+ _02941_ sky130_fd_sc_hd__mux2_1
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19160_ _06225_ _06224_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__and2b_1
X_16372_ _03747_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28358_ clknet_leaf_74_clk _02156_ VGND VGND VPWR VPWR systolic_inst.B_shift\[22\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13584_ deser_B.word_buffer\[20\] deser_B.serial_word\[20\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15323_ systolic_inst.acc_wires\[14\]\[24\] systolic_inst.acc_wires\[14\]\[25\] systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12411_ sky130_fd_sc_hd__o21a_1
X_18111_ _05297_ _05298_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27309_ clknet_leaf_300_clk _01107_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19091_ _06150_ _06158_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__nor2_1
XFILLER_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28289_ clknet_leaf_75_clk _02087_ VGND VGND VPWR VPWR systolic_inst.B_shift\[19\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_321_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_321_clk
+ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_2_2__f_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_2_2__leaf_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15254_ _12343_ _12351_ VGND VGND VPWR VPWR _12352_ sky130_fd_sc_hd__or2_1
XFILLER_9_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18042_ _05232_ _05231_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__nand2b_1
XFILLER_201_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_186_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14205_ _11392_ _11393_ VGND VGND VPWR VPWR _11394_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_186_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15185_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[14\]\[6\]
+ VGND VGND VPWR VPWR _12293_ sky130_fd_sc_hd__nand2_1
XFILLER_99_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14136_ systolic_inst.B_outs\[14\]\[4\] systolic_inst.B_outs\[10\]\[4\] net120 VGND
+ VGND VPWR VPWR _00958_ sky130_fd_sc_hd__mux2_1
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19993_ _06923_ _06965_ _06964_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__o21a_1
XFILLER_193_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_203_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14067_ deser_B.shift_reg\[101\] deser_B.shift_reg\[102\] net126 VGND VGND VPWR VPWR
+ _00893_ sky130_fd_sc_hd__mux2_1
X_18944_ _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__inv_2
XFILLER_234_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18875_ _05956_ _05960_ _05963_ _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__a211o_1
XFILLER_80_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17826_ _05017_ _05023_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__or2_1
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17757_ _04972_ _04976_ _04973_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__a21bo_1
X_14969_ _12047_ _12049_ _12088_ VGND VGND VPWR VPWR _12090_ sky130_fd_sc_hd__nand3_1
XFILLER_242_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16708_ _04028_ _04029_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__or2_1
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17688_ _04919_ _04920_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__nand2_1
XFILLER_222_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19427_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[7\]\[4\]
+ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__nand2_1
XFILLER_223_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16639_ _03952_ _03955_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_139_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19358_ _06415_ _06416_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__xor2_1
XFILLER_241_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18309_ _05469_ _05472_ _05471_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_171_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19289_ systolic_inst.A_outs\[7\]\[5\] systolic_inst.B_outs\[7\]\[6\] _11261_ systolic_inst.A_outs\[7\]\[4\]
+ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_312_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_312_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_241_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21320_ net63 _08173_ _08174_ systolic_inst.acc_wires\[4\]\[10\] _11258_ VGND VGND
+ VPWR VPWR _01692_ sky130_fd_sc_hd__a32o_1
XFILLER_50_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21251_ _11258_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] _08110_
+ _08116_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__a22o_1
Xmax_cap130 deser_A.receiving VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_12
XFILLER_11_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20202_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[28\]
+ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__nand2_1
XFILLER_143_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21182_ _08050_ _08026_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__nand2b_1
XFILLER_172_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20133_ net106 systolic_inst.acc_wires\[6\]\[17\] net62 _07108_ VGND VGND VPWR VPWR
+ _01571_ sky130_fd_sc_hd__a22o_1
X_25990_ systolic_inst.acc_wires\[14\]\[18\] ser_C.parallel_data\[466\] net25 VGND
+ VGND VPWR VPWR _03292_ sky130_fd_sc_hd__mux2_1
X_20064_ _07045_ _07046_ _07044_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__a21bo_1
XFILLER_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24941_ C_out\[297\] net102 net76 ser_C.shift_reg\[297\] _10940_ VGND VGND VPWR VPWR
+ _02547_ sky130_fd_sc_hd__a221o_1
XFILLER_213_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27660_ clknet_leaf_211_clk _01458_ net147 VGND VGND VPWR VPWR systolic_inst.A_outs\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_24872_ net110 ser_C.shift_reg\[264\] VGND VGND VPWR VPWR _10906_ sky130_fd_sc_hd__and2_1
XFILLER_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23823_ _10402_ _10407_ _10412_ _10416_ VGND VGND VPWR VPWR _10420_ sky130_fd_sc_hd__or4_1
X_26611_ clknet_leaf_16_B_in_serial_clk _00414_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27591_ clknet_leaf_223_clk _01389_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26542_ clknet_leaf_20_A_in_serial_clk _00345_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_29330_ clknet_leaf_220_clk _03128_ net139 VGND VGND VPWR VPWR C_out\[302\] sky130_fd_sc_hd__dfrtp_1
X_23754_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[0\]\[10\]
+ VGND VGND VPWR VPWR _10361_ sky130_fd_sc_hd__nand2_1
XFILLER_241_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20966_ systolic_inst.B_outs\[4\]\[7\] _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__xnor2_1
XFILLER_213_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22705_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.A_outs\[1\]\[1\] systolic_inst.B_outs\[1\]\[2\]
+ systolic_inst.B_outs\[1\]\[3\] VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__and4_1
X_29261_ clknet_leaf_198_clk _03059_ net146 VGND VGND VPWR VPWR C_out\[233\] sky130_fd_sc_hd__dfrtp_1
X_26473_ clknet_leaf_14_A_in_serial_clk _00276_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_23685_ net122 systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[14\] VGND
+ VGND VPWR VPWR _10304_ sky130_fd_sc_hd__nor2_1
XFILLER_81_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20897_ net108 systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[4\] _07771_
+ _07773_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__a22o_1
XFILLER_202_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28212_ clknet_leaf_72_clk _02010_ VGND VGND VPWR VPWR systolic_inst.B_shift\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25424_ _11181_ systolic_inst.A_shift\[0\]\[3\] net70 VGND VGND VPWR VPWR _02789_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22636_ net65 _09346_ _09347_ systolic_inst.acc_wires\[2\]\[25\] net109 VGND VGND
+ VPWR VPWR _01835_ sky130_fd_sc_hd__a32o_1
X_29192_ clknet_leaf_217_clk _02990_ net140 VGND VGND VPWR VPWR C_out\[164\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_230_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_230_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28143_ clknet_leaf_122_clk _01941_ net153 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_181_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25355_ ser_C.parallel_data\[504\] net98 net78 ser_C.shift_reg\[504\] _11147_ VGND
+ VGND VPWR VPWR _02754_ sky130_fd_sc_hd__a221o_1
XFILLER_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22567_ _09286_ _09288_ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_133_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_303_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_303_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_220_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24306_ _10626_ systolic_inst.A_shift\[10\]\[0\] net71 VGND VGND VPWR VPWR _02226_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28074_ clknet_leaf_119_clk _01872_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_21518_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[3\]
+ systolic_inst.A_outs\[3\]\[4\] VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_40_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25286_ net111 ser_C.shift_reg\[471\] VGND VGND VPWR VPWR _11113_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22498_ net65 _09228_ _09230_ systolic_inst.acc_wires\[2\]\[4\] net109 VGND VGND
+ VPWR VPWR _01814_ sky130_fd_sc_hd__a32o_1
XFILLER_177_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_125_Left_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27025_ clknet_leaf_19_B_in_serial_clk _00823_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24237_ systolic_inst.A_shift\[19\]\[2\] A_in\[66\] net59 VGND VGND VPWR VPWR _10604_
+ sky130_fd_sc_hd__mux2_1
XFILLER_181_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21449_ _08278_ _08281_ _08280_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__o21a_1
XFILLER_120_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24168_ _10585_ systolic_inst.A_shift\[27\]\[7\] net70 VGND VGND VPWR VPWR _02129_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23119_ _09780_ _09781_ _09779_ VGND VGND VPWR VPWR _09784_ sky130_fd_sc_hd__a21bo_1
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24099_ systolic_inst.B_shift\[23\]\[5\] B_in\[61\] _00008_ VGND VGND VPWR VPWR _10559_
+ sky130_fd_sc_hd__mux2_1
X_28976_ clknet_leaf_64_clk _02774_ VGND VGND VPWR VPWR systolic_inst.A_shift\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16990_ _04296_ _04297_ _04298_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__and3_1
XFILLER_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27927_ clknet_leaf_134_clk _01725_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_15941_ net107 systolic_inst.acc_wires\[13\]\[28\] net67 _12962_ VGND VGND VPWR VPWR
+ _01134_ sky130_fd_sc_hd__a22o_1
XFILLER_7_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _05786_ _05785_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__nand2b_1
X_15872_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[18\]
+ VGND VGND VPWR VPWR _12904_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27858_ clknet_leaf_35_clk _01656_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_134_Left_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17611_ _04854_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_237_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26809_ clknet_leaf_84_clk _00611_ net144 VGND VGND VPWR VPWR B_in\[81\] sky130_fd_sc_hd__dfrtp_1
X_14823_ _11942_ _11947_ VGND VGND VPWR VPWR _11948_ sky130_fd_sc_hd__nand2b_1
X_18591_ _05717_ _05718_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_237_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27789_ clknet_leaf_40_clk _01587_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_40_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29528_ clknet_leaf_262_clk _03326_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[500\]
+ sky130_fd_sc_hd__dfrtp_1
X_17542_ _04763_ _04768_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__o21ai_1
XFILLER_217_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14754_ systolic_inst.B_outs\[13\]\[6\] systolic_inst.B_outs\[9\]\[6\] net115 VGND
+ VGND VPWR VPWR _01024_ sky130_fd_sc_hd__mux2_1
XFILLER_205_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13705_ B_in\[12\] deser_B.word_buffer\[12\] net84 VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__mux2_1
XFILLER_204_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29459_ clknet_leaf_328_clk _03257_ net136 VGND VGND VPWR VPWR C_out\[431\] sky130_fd_sc_hd__dfrtp_1
X_14685_ _11832_ _11836_ _11839_ VGND VGND VPWR VPWR _11840_ sky130_fd_sc_hd__nand3_1
X_17473_ _04725_ _04726_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__nand2_1
XFILLER_229_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19212_ _06274_ _06275_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__or2_1
X_13636_ deser_B.word_buffer\[72\] deser_B.serial_word\[72\] net123 VGND VGND VPWR
+ VPWR _00473_ sky130_fd_sc_hd__mux2_1
X_16424_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[12\]\[8\]
+ _03790_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__and3_1
XFILLER_60_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_188_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19143_ systolic_inst.B_outs\[7\]\[3\] systolic_inst.A_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\]
+ systolic_inst.A_outs\[7\]\[4\] VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_188_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13567_ deser_B.word_buffer\[3\] deser_B.serial_word\[3\] net124 VGND VGND VPWR VPWR
+ _00404_ sky130_fd_sc_hd__mux2_1
XFILLER_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16355_ _03681_ _03686_ _03709_ _03710_ _03731_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__o311a_1
XFILLER_34_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_143_Left_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15306_ _12375_ _12382_ _12387_ _12392_ VGND VGND VPWR VPWR _12396_ sky130_fd_sc_hd__nand4_1
XFILLER_9_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19074_ net105 _06141_ _06142_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__or3_1
X_16286_ _03633_ _03635_ _03634_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_184_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13498_ deser_A.shift_reg\[62\] deser_A.shift_reg\[63\] net130 VGND VGND VPWR VPWR
+ _00335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_184_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18025_ _05180_ _05183_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__nand2_1
X_15237_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[14\]\[12\]
+ _12335_ VGND VGND VPWR VPWR _12338_ sky130_fd_sc_hd__and3_1
XFILLER_161_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15168_ _12278_ VGND VGND VPWR VPWR _12279_ sky130_fd_sc_hd__inv_2
XFILLER_154_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14119_ systolic_inst.A_shift\[21\]\[3\] net71 _11333_ A_in\[91\] VGND VGND VPWR
+ VPWR _00941_ sky130_fd_sc_hd__a22o_1
X_19976_ _06939_ _06941_ _06971_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__nor3_1
XFILLER_140_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15099_ _12214_ _12215_ VGND VGND VPWR VPWR _12216_ sky130_fd_sc_hd__nand2_1
XFILLER_140_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18927_ _06028_ _06029_ _06027_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__a21o_1
XFILLER_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_152_Left_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18858_ _05968_ _05969_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__or2_1
XFILLER_95_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17809_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.A_outs\[9\]\[2\] VGND VGND VPWR
+ VPWR _05008_ sky130_fd_sc_hd__nand2_1
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18789_ _05910_ _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__xor2_1
XFILLER_227_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20820_ _07715_ _07718_ VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__nand2_1
XFILLER_70_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20751_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[20\]
+ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_173_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23470_ _10091_ _10093_ _10050_ _10052_ VGND VGND VPWR VPWR _10095_ sky130_fd_sc_hd__o211a_1
XFILLER_56_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20682_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[5\]\[10\]
+ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__nand2_1
XFILLER_189_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22421_ _09159_ _09160_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__and2_1
XFILLER_195_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25140_ net110 ser_C.shift_reg\[398\] VGND VGND VPWR VPWR _11040_ sky130_fd_sc_hd__and2_1
X_22352_ systolic_inst.B_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\] VGND VGND VPWR
+ VPWR _09094_ sky130_fd_sc_hd__or2_1
XFILLER_148_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21303_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[4\]\[8\]
+ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__nand2_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25071_ C_out\[362\] net97 net77 ser_C.shift_reg\[362\] _11005_ VGND VGND VPWR VPWR
+ _02612_ sky130_fd_sc_hd__a221o_1
X_22283_ systolic_inst.B_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[5\]
+ systolic_inst.A_outs\[2\]\[6\] VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__and4_1
XFILLER_219_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24022_ systolic_inst.B_shift\[6\]\[5\] _11332_ net83 systolic_inst.B_shift\[10\]\[5\]
+ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__a22o_1
XFILLER_85_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21234_ _08069_ _08076_ _08099_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1003 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28830_ clknet_leaf_194_clk _02628_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[378\]
+ sky130_fd_sc_hd__dfrtp_1
X_21165_ systolic_inst.A_outs\[4\]\[6\] systolic_inst.B_outs\[4\]\[6\] VGND VGND VPWR
+ VPWR _08034_ sky130_fd_sc_hd__nand2_1
XFILLER_213_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20116_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[15\]
+ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__and2_1
XFILLER_132_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28761_ clknet_leaf_215_clk _02559_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[309\]
+ sky130_fd_sc_hd__dfrtp_1
X_21096_ _07963_ _07966_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__xnor2_1
X_25973_ systolic_inst.acc_wires\[14\]\[1\] ser_C.parallel_data\[449\] net24 VGND
+ VGND VPWR VPWR _03275_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27712_ clknet_leaf_192_clk _01510_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20047_ _07032_ _07033_ _07034_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__a21o_1
X_24924_ net111 ser_C.shift_reg\[290\] VGND VGND VPWR VPWR _10932_ sky130_fd_sc_hd__and2_1
X_28692_ clknet_leaf_193_clk _02490_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[240\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27643_ clknet_leaf_311_clk _01441_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_24855_ C_out\[254\] net99 net79 ser_C.shift_reg\[254\] _10897_ VGND VGND VPWR VPWR
+ _02504_ sky130_fd_sc_hd__a221o_1
XFILLER_233_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23806_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[17\]
+ VGND VGND VPWR VPWR _10406_ sky130_fd_sc_hd__xor2_2
XFILLER_215_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24786_ net113 ser_C.shift_reg\[221\] VGND VGND VPWR VPWR _10863_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_83_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27574_ clknet_leaf_304_clk _01372_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_233_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21998_ _08773_ _08777_ _08779_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__a21oi_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_232_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29313_ clknet_leaf_301_clk _03111_ net141 VGND VGND VPWR VPWR C_out\[285\] sky130_fd_sc_hd__dfrtp_1
X_23737_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[0\]\[7\]
+ VGND VGND VPWR VPWR _10347_ sky130_fd_sc_hd__or2_1
XFILLER_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26525_ clknet_leaf_4_A_in_serial_clk _00328_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_232_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20949_ _07822_ _07823_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_42_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29244_ clknet_leaf_187_clk _03042_ net148 VGND VGND VPWR VPWR C_out\[216\] sky130_fd_sc_hd__dfrtp_1
X_14470_ systolic_inst.A_outs\[15\]\[6\] _11273_ VGND VGND VPWR VPWR _11651_ sky130_fd_sc_hd__or2_1
X_23668_ systolic_inst.B_outs\[0\]\[7\] _11270_ _10120_ VGND VGND VPWR VPWR _10287_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_42_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26456_ clknet_leaf_10_clk _00263_ net132 VGND VGND VPWR VPWR A_in\[124\] sky130_fd_sc_hd__dfrtp_1
XFILLER_109_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13421_ deser_A.bit_idx\[1\] _11308_ VGND VGND VPWR VPWR _11309_ sky130_fd_sc_hd__and2_1
X_22619_ _09332_ VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__inv_2
X_25407_ systolic_inst.A_shift\[2\]\[3\] A_in\[11\] net59 VGND VGND VPWR VPWR _11173_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29175_ clknet_leaf_138_clk _02973_ net142 VGND VGND VPWR VPWR C_out\[147\] sky130_fd_sc_hd__dfrtp_1
X_26387_ clknet_leaf_15_clk _00194_ net133 VGND VGND VPWR VPWR A_in\[55\] sky130_fd_sc_hd__dfrtp_1
XFILLER_224_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23599_ _10145_ _10190_ _10189_ VGND VGND VPWR VPWR _10220_ sky130_fd_sc_hd__a21o_1
XFILLER_201_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16140_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[6\] VGND VGND
+ VPWR VPWR _03525_ sky130_fd_sc_hd__nand2_1
XFILLER_70_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28126_ clknet_leaf_50_clk _01924_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25338_ net112 ser_C.shift_reg\[497\] VGND VGND VPWR VPWR _11139_ sky130_fd_sc_hd__and2_1
X_13352_ A_in\[61\] deser_A.word_buffer\[61\] net91 VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_26_B_in_serial_clk clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_26_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_23_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16071_ _13063_ _13066_ VGND VGND VPWR VPWR _13067_ sky130_fd_sc_hd__xnor2_1
X_28057_ clknet_leaf_97_clk _01855_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_25269_ ser_C.parallel_data\[461\] net102 net74 ser_C.shift_reg\[461\] _11104_ VGND
+ VGND VPWR VPWR _02711_ sky130_fd_sc_hd__a221o_1
X_13283_ deser_A.word_buffer\[121\] deser_A.serial_word\[121\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__mux2_1
XFILLER_136_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15022_ _12031_ _12140_ VGND VGND VPWR VPWR _12141_ sky130_fd_sc_hd__or2_1
X_27008_ clknet_leaf_16_B_in_serial_clk _00806_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19830_ systolic_inst.A_outs\[6\]\[4\] systolic_inst.B_outs\[6\]\[5\] VGND VGND VPWR
+ VPWR _06830_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19761_ _06756_ _06762_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__nor2_1
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_239_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28959_ clknet_leaf_257_clk _02757_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[507\]
+ sky130_fd_sc_hd__dfrtp_1
X_16973_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[11\]\[1\]
+ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__nand2_1
XFILLER_89_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18712_ systolic_inst.A_outs\[8\]\[5\] systolic_inst.B_outs\[8\]\[6\] systolic_inst.A_outs\[8\]\[6\]
+ systolic_inst.B_outs\[8\]\[7\] VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__and4b_1
X_15924_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[26\]
+ VGND VGND VPWR VPWR _12948_ sky130_fd_sc_hd__nand2_1
XFILLER_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19692_ systolic_inst.A_outs\[6\]\[2\] systolic_inst.B_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\]
+ systolic_inst.A_outs\[6\]\[1\] VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__a22o_1
XFILLER_232_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18643_ _05735_ _05769_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_177_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _12880_ _12885_ _12889_ VGND VGND VPWR VPWR _12890_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14806_ net107 _11930_ _11931_ VGND VGND VPWR VPWR _11932_ sky130_fd_sc_hd__or3_1
X_18574_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[6\] VGND VGND VPWR
+ VPWR _05703_ sky130_fd_sc_hd__nand2_1
XFILLER_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15786_ _12830_ VGND VGND VPWR VPWR _12831_ sky130_fd_sc_hd__inv_2
X_17525_ _04744_ _04747_ _04775_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__or3_1
X_14737_ _11878_ _11882_ _11883_ VGND VGND VPWR VPWR _11884_ sky130_fd_sc_hd__a21oi_1
XFILLER_233_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_162_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17456_ _04602_ _04708_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__nand2_1
XFILLER_221_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14668_ _11823_ _11824_ _11821_ VGND VGND VPWR VPWR _11826_ sky130_fd_sc_hd__o21ai_2
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_215_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16407_ _03769_ _03772_ _03774_ _03776_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__o211a_1
XFILLER_20_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13619_ deser_B.word_buffer\[55\] deser_B.serial_word\[55\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__mux2_1
X_17387_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[7\] VGND VGND
+ VPWR VPWR _04643_ sky130_fd_sc_hd__nand2_4
XFILLER_242_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14599_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[15\]\[11\]
+ VGND VGND VPWR VPWR _11766_ sky130_fd_sc_hd__nor2_1
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19126_ _06190_ _06191_ _06168_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16338_ _03632_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__or2_1
XFILLER_145_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19057_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.A_outs\[7\]\[1\] systolic_inst.B_outs\[7\]\[3\]
+ systolic_inst.B_outs\[7\]\[4\] VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__nand4_1
X_16269_ _03613_ _03615_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__and3_1
XFILLER_103_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18008_ _05196_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_160_Left_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19959_ _06953_ _06954_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__nor2_1
XFILLER_101_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22970_ _09609_ _09611_ _09646_ VGND VGND VPWR VPWR _09648_ sky130_fd_sc_hd__a21o_1
XFILLER_228_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21921_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[3\]\[9\]
+ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_121_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24640_ net7 ser_C.shift_reg\[148\] VGND VGND VPWR VPWR _10790_ sky130_fd_sc_hd__and2_1
XFILLER_23_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21852_ _08584_ _08632_ _08631_ VGND VGND VPWR VPWR _08655_ sky130_fd_sc_hd__o21ba_1
XFILLER_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20803_ systolic_inst.acc_wires\[5\]\[26\] systolic_inst.acc_wires\[5\]\[27\] systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__o21a_1
XFILLER_212_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24571_ C_out\[112\] net100 net80 ser_C.shift_reg\[112\] _10755_ VGND VGND VPWR VPWR
+ _02362_ sky130_fd_sc_hd__a221o_1
XFILLER_82_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21783_ systolic_inst.A_outs\[3\]\[5\] systolic_inst.B_outs\[3\]\[6\] systolic_inst.A_outs\[3\]\[6\]
+ systolic_inst.B_outs\[3\]\[7\] VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__and4b_1
XFILLER_93_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_93_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23522_ systolic_inst.B_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[5\] _10025_ VGND
+ VGND VPWR VPWR _10145_ sky130_fd_sc_hd__and3_1
X_26310_ clknet_leaf_28_A_in_serial_clk _00118_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_169_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20734_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[17\]
+ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__xor2_2
X_27290_ clknet_leaf_319_clk _01088_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_223_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26241_ clknet_leaf_17_A_in_serial_clk _00049_ net143 VGND VGND VPWR VPWR deser_A.word_buffer\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23453_ systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[7\] VGND VGND VPWR
+ VPWR _10078_ sky130_fd_sc_hd__nand2b_1
XFILLER_11_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20665_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[5\]\[7\]
+ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_119_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22404_ _09091_ _09144_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__and2b_1
XFILLER_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26172_ deser_B.serial_word\[127\] deser_B.shift_reg\[127\] net56 VGND VGND VPWR
+ VPWR _03474_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23384_ _10008_ _10009_ VGND VGND VPWR VPWR _10011_ sky130_fd_sc_hd__xor2_1
X_20596_ _07525_ _07526_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_115_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25123_ C_out\[388\] net101 net73 ser_C.shift_reg\[388\] _11031_ VGND VGND VPWR VPWR
+ _02638_ sky130_fd_sc_hd__a221o_1
XFILLER_52_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22335_ _09024_ _09041_ _09039_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__o21a_1
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25054_ net112 ser_C.shift_reg\[355\] VGND VGND VPWR VPWR _10997_ sky130_fd_sc_hd__and2_1
X_22266_ _09008_ _09009_ VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__xor2_1
XFILLER_219_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24005_ systolic_inst.B_shift\[9\]\[6\] B_in\[14\] _00008_ VGND VGND VPWR VPWR _10528_
+ sky130_fd_sc_hd__mux2_1
X_21217_ _08083_ _08084_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__and2b_1
X_22197_ _08913_ _08943_ VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_221_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28813_ clknet_leaf_243_clk _02611_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[361\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_221_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21148_ _08015_ _08016_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_89_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28744_ clknet_leaf_297_clk _02542_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[292\]
+ sky130_fd_sc_hd__dfrtp_1
X_13970_ deser_B.shift_reg\[4\] deser_B.shift_reg\[5\] net125 VGND VGND VPWR VPWR
+ _00796_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25956_ systolic_inst.acc_wires\[13\]\[16\] C_out\[432\] net20 VGND VGND VPWR VPWR
+ _03258_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21079_ _07949_ _07950_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__xnor2_1
XFILLER_219_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24907_ C_out\[280\] net103 net75 ser_C.shift_reg\[280\] _10923_ VGND VGND VPWR VPWR
+ _02530_ sky130_fd_sc_hd__a221o_1
X_28675_ clknet_leaf_184_clk _02473_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[223\]
+ sky130_fd_sc_hd__dfrtp_1
X_25887_ systolic_inst.acc_wires\[11\]\[11\] C_out\[363\] net39 VGND VGND VPWR VPWR
+ _03189_ sky130_fd_sc_hd__mux2_1
XFILLER_219_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15640_ _12692_ _12693_ VGND VGND VPWR VPWR _12695_ sky130_fd_sc_hd__xnor2_1
X_27626_ clknet_leaf_311_clk _01424_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24838_ net113 ser_C.shift_reg\[247\] VGND VGND VPWR VPWR _10889_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_219_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15571_ _12625_ _12626_ VGND VGND VPWR VPWR _12628_ sky130_fd_sc_hd__xnor2_1
X_27557_ clknet_leaf_305_clk _01355_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24769_ C_out\[211\] net98 net78 ser_C.shift_reg\[211\] _10854_ VGND VGND VPWR VPWR
+ _02461_ sky130_fd_sc_hd__a221o_1
XFILLER_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_29_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17310_ _04538_ _04540_ _04566_ _04567_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__a211o_1
X_14522_ _11619_ _11680_ VGND VGND VPWR VPWR _11701_ sky130_fd_sc_hd__xnor2_1
X_26508_ clknet_leaf_17_A_in_serial_clk _00311_ net143 VGND VGND VPWR VPWR deser_A.shift_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _05454_ _05458_ _05459_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__nand3_1
XFILLER_186_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27488_ clknet_leaf_228_clk _01286_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29227_ clknet_leaf_211_clk _03025_ net147 VGND VGND VPWR VPWR C_out\[199\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17241_ _04483_ _04500_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__nor2_1
XFILLER_230_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26439_ clknet_leaf_0_clk _00246_ net132 VGND VGND VPWR VPWR A_in\[107\] sky130_fd_sc_hd__dfrtp_1
X_14453_ _11622_ _11634_ VGND VGND VPWR VPWR _11635_ sky130_fd_sc_hd__xor2_1
XFILLER_70_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13404_ A_in\[113\] deser_A.word_buffer\[113\] _00003_ VGND VGND VPWR VPWR _00252_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17172_ _04450_ _04453_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__or2_1
X_14384_ _11565_ _11566_ VGND VGND VPWR VPWR _11568_ sky130_fd_sc_hd__xnor2_1
X_29158_ clknet_leaf_309_clk _02956_ net142 VGND VGND VPWR VPWR C_out\[130\] sky130_fd_sc_hd__dfrtp_1
XFILLER_128_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_210_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_210_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28109_ clknet_leaf_57_clk _01907_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_127_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16123_ _13084_ _03507_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__xnor2_1
X_13335_ A_in\[44\] deser_A.word_buffer\[44\] net95 VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__mux2_1
XFILLER_122_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29089_ clknet_leaf_157_clk _02887_ net150 VGND VGND VPWR VPWR C_out\[61\] sky130_fd_sc_hd__dfrtp_1
XFILLER_116_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16054_ _13026_ _13049_ VGND VGND VPWR VPWR _13051_ sky130_fd_sc_hd__xnor2_1
X_13266_ deser_A.word_buffer\[104\] deser_A.serial_word\[104\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__mux2_1
XFILLER_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15005_ _12122_ _12123_ VGND VGND VPWR VPWR _12125_ sky130_fd_sc_hd__xor2_1
X_13197_ deser_A.word_buffer\[35\] deser_A.serial_word\[35\] net127 VGND VGND VPWR
+ VPWR _00045_ sky130_fd_sc_hd__mux2_1
XFILLER_194_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19813_ _06811_ _06812_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__and2_1
XFILLER_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19744_ _06744_ _06745_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16956_ _04268_ _04269_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15907_ _12925_ _12929_ _12932_ VGND VGND VPWR VPWR _12934_ sky130_fd_sc_hd__a21o_1
X_19675_ _06677_ _06678_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__xnor2_1
XFILLER_225_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16887_ systolic_inst.B_outs\[11\]\[5\] systolic_inst.A_outs\[11\]\[7\] VGND VGND
+ VPWR VPWR _04204_ sky130_fd_sc_hd__nand2_1
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18626_ _05753_ _05752_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__nand2b_1
X_15838_ _12869_ _12873_ VGND VGND VPWR VPWR _12875_ sky130_fd_sc_hd__nand2b_1
XFILLER_225_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18557_ _05655_ _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__and2b_1
XFILLER_75_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15769_ _12809_ _12810_ _12808_ VGND VGND VPWR VPWR _12816_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_44_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17508_ _04709_ _04759_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__xor2_1
XFILLER_178_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18488_ _05589_ _05591_ _05618_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__or3_1
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_14 systolic_inst.load_acc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _04642_ _04659_ _04657_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__o21a_1
XANTENNA_25 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_36 net153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 net153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20450_ _07359_ _07385_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19109_ systolic_inst.A_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[3\] systolic_inst.A_outs\[7\]\[3\]
+ systolic_inst.B_outs\[7\]\[4\] VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_168_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20381_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[7\] _07318_ net120
+ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__mux2_1
XFILLER_238_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22120_ _08855_ _08857_ _08868_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_110_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22051_ _08811_ _08816_ VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__nand2_1
XFILLER_138_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21002_ systolic_inst.A_outs\[4\]\[4\] systolic_inst.B_outs\[4\]\[4\] systolic_inst.A_outs\[4\]\[5\]
+ systolic_inst.B_outs\[4\]\[3\] VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__a22o_1
XFILLER_47_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25810_ systolic_inst.acc_wires\[8\]\[30\] C_out\[286\] net27 VGND VGND VPWR VPWR
+ _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_214_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26790_ clknet_leaf_74_clk _00592_ net153 VGND VGND VPWR VPWR B_in\[62\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25741_ systolic_inst.acc_wires\[6\]\[25\] C_out\[217\] net44 VGND VGND VPWR VPWR
+ _03043_ sky130_fd_sc_hd__mux2_1
X_22953_ _09629_ _09630_ VGND VGND VPWR VPWR _09631_ sky130_fd_sc_hd__or2_1
XFILLER_101_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap16 net32 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_8
XFILLER_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21904_ net68 _08697_ _08699_ systolic_inst.acc_wires\[3\]\[5\] net106 VGND VGND
+ VPWR VPWR _01751_ sky130_fd_sc_hd__a32o_1
Xmax_cap27 net28 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_4
X_28460_ clknet_leaf_97_clk _02258_ net153 VGND VGND VPWR VPWR ser_C.shift_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap38 net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_4
Xmax_cap49 net51 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_6
X_22884_ systolic_inst.A_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[6\] _11277_ systolic_inst.A_outs\[1\]\[2\]
+ VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__o2bb2a_1
X_25672_ systolic_inst.acc_wires\[4\]\[20\] C_out\[148\] net32 VGND VGND VPWR VPWR
+ _02974_ sky130_fd_sc_hd__mux2_1
XFILLER_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27411_ clknet_leaf_226_clk _01209_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_21835_ _08607_ _08612_ _08637_ net122 VGND VGND VPWR VPWR _08639_ sky130_fd_sc_hd__o31a_1
X_24623_ C_out\[138\] net103 net75 ser_C.shift_reg\[138\] _10781_ VGND VGND VPWR VPWR
+ _02388_ sky130_fd_sc_hd__a221o_1
XFILLER_58_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28391_ clknet_leaf_32_clk _02189_ VGND VGND VPWR VPWR systolic_inst.A_shift\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_203_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_35_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24554_ net113 ser_C.shift_reg\[105\] VGND VGND VPWR VPWR _10747_ sky130_fd_sc_hd__and2_1
XFILLER_145_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27342_ clknet_leaf_342_clk _01140_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_54_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21766_ _08571_ _08570_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__and2b_1
XFILLER_196_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20717_ _07629_ _07631_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__nand2_1
X_23505_ _10118_ _10126_ VGND VGND VPWR VPWR _10129_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_117_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24485_ C_out\[69\] _11302_ net81 ser_C.shift_reg\[69\] _10712_ VGND VGND VPWR VPWR
+ _02319_ sky130_fd_sc_hd__a221o_1
X_27273_ clknet_leaf_266_clk _01071_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21697_ _08502_ _08503_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29012_ clknet_leaf_103_clk _02810_ net151 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23436_ _10059_ _10060_ _10019_ _10021_ VGND VGND VPWR VPWR _10062_ sky130_fd_sc_hd__a211o_1
XFILLER_156_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26224_ clknet_leaf_6_A_in_serial_clk _00032_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_20648_ _07572_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__inv_2
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26155_ deser_B.serial_word\[110\] deser_B.shift_reg\[110\] _00001_ VGND VGND VPWR
+ VPWR _03457_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23367_ _09972_ _09992_ VGND VGND VPWR VPWR _09994_ sky130_fd_sc_hd__xnor2_1
X_20579_ _07508_ _07509_ VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__and2b_1
X_13120_ systolic_inst.B_outs\[5\]\[7\] VGND VGND VPWR VPWR _11276_ sky130_fd_sc_hd__inv_2
XFILLER_137_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22318_ systolic_inst.A_outs\[2\]\[6\] _09060_ _09059_ VGND VGND VPWR VPWR _09061_
+ sky130_fd_sc_hd__a21bo_1
X_25106_ net113 ser_C.shift_reg\[381\] VGND VGND VPWR VPWR _11023_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_223_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26086_ deser_B.serial_word\[41\] deser_B.shift_reg\[41\] net55 VGND VGND VPWR VPWR
+ _03388_ sky130_fd_sc_hd__mux2_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_223_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23298_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[2\] _09928_ net121
+ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__mux2_1
XFILLER_3_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25037_ C_out\[345\] net97 net77 ser_C.shift_reg\[345\] _10988_ VGND VGND VPWR VPWR
+ _02595_ sky130_fd_sc_hd__a221o_1
XFILLER_69_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22249_ _08992_ _08993_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16810_ _04057_ _04127_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17790_ systolic_inst.A_outs\[9\]\[5\] systolic_inst.A_outs\[8\]\[5\] net117 VGND
+ VGND VPWR VPWR _01335_ sky130_fd_sc_hd__mux2_1
XFILLER_232_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26988_ clknet_leaf_30_A_in_serial_clk _00786_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28727_ clknet_leaf_325_clk _02525_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[275\]
+ sky130_fd_sc_hd__dfrtp_1
X_16741_ systolic_inst.B_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[4\]
+ systolic_inst.A_outs\[11\]\[5\] VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__and4_1
X_25939_ systolic_inst.acc_wires\[12\]\[31\] C_out\[415\] net21 VGND VGND VPWR VPWR
+ _03241_ sky130_fd_sc_hd__mux2_1
X_13953_ deser_A.serial_word\[114\] deser_A.shift_reg\[114\] net57 VGND VGND VPWR
+ VPWR _00779_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19460_ _06502_ _06505_ _06507_ _06504_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__a211o_1
X_28658_ clknet_leaf_204_clk _02456_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[206\]
+ sky130_fd_sc_hd__dfrtp_1
X_16672_ systolic_inst.A_outs\[11\]\[2\] systolic_inst.B_outs\[11\]\[3\] systolic_inst.A_outs\[11\]\[3\]
+ systolic_inst.B_outs\[11\]\[4\] VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__nand4_2
XFILLER_98_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13884_ deser_A.serial_word\[45\] deser_A.shift_reg\[45\] net58 VGND VGND VPWR VPWR
+ _00710_ sky130_fd_sc_hd__mux2_1
XFILLER_207_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18411_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[3\]\[0\] net119 VGND
+ VGND VPWR VPWR _01402_ sky130_fd_sc_hd__mux2_1
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27609_ clknet_leaf_204_clk _01407_ net146 VGND VGND VPWR VPWR systolic_inst.B_outs\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_15623_ net107 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[10\] VGND
+ VGND VPWR VPWR _12679_ sky130_fd_sc_hd__and2_1
X_19391_ _06425_ _06449_ _06427_ _06401_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__a2bb2o_1
X_28589_ clknet_leaf_40_clk _02387_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[137\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
X_18342_ systolic_inst.acc_wires\[9\]\[20\] systolic_inst.acc_wires\[9\]\[21\] systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_191_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _12574_ _12580_ _12579_ VGND VGND VPWR VPWR _12611_ sky130_fd_sc_hd__a21o_1
XFILLER_199_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14505_ _11683_ _11684_ VGND VGND VPWR VPWR _11685_ sky130_fd_sc_hd__nor2_1
XFILLER_72_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_212_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[9\]\[12\]
+ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__or2_1
XFILLER_230_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15485_ _12543_ _12539_ VGND VGND VPWR VPWR _12544_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_13_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17224_ net107 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[3\] _04483_
+ _04485_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__a22o_1
XFILLER_30_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14436_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[7\] _11591_ _11558_
+ VGND VGND VPWR VPWR _11618_ sky130_fd_sc_hd__a31o_1
XFILLER_198_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17155_ _04424_ _04426_ _04438_ _04439_ _04432_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__a311oi_4
X_14367_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[9\] _11551_ net118
+ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__mux2_1
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16106_ systolic_inst.A_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[7\] VGND VGND
+ VPWR VPWR _03492_ sky130_fd_sc_hd__and2b_1
X_13318_ A_in\[27\] deser_A.word_buffer\[27\] net91 VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__mux2_1
XFILLER_116_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14298_ systolic_inst.B_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[5\]
+ systolic_inst.B_outs\[15\]\[3\] VGND VGND VPWR VPWR _11484_ sky130_fd_sc_hd__a22oi_1
X_17086_ _04381_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_208_Right_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16037_ _13011_ _13032_ VGND VGND VPWR VPWR _13034_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13249_ deser_A.word_buffer\[87\] deser_A.serial_word\[87\] net127 VGND VGND VPWR
+ VPWR _00097_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17988_ _05178_ _05179_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_144_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19727_ _06724_ _06728_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__xor2_1
XFILLER_211_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16939_ systolic_inst.B_outs\[11\]\[5\] systolic_inst.B_outs\[11\]\[6\] systolic_inst.A_outs\[11\]\[7\]
+ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_0_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19658_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[2\] VGND VGND VPWR
+ VPWR _06663_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18609_ systolic_inst.B_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[5\]
+ systolic_inst.A_outs\[8\]\[6\] VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_157_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19589_ _06602_ _06604_ _06616_ _06617_ _06610_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__a311oi_4
XFILLER_168_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
X_21620_ _08378_ _08379_ _08392_ _08391_ _08360_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__o32a_1
XFILLER_181_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21551_ _08362_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__inv_2
XFILLER_139_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20502_ systolic_inst.B_outs\[5\]\[5\] systolic_inst.A_outs\[5\]\[6\] VGND VGND VPWR
+ VPWR _07436_ sky130_fd_sc_hd__nand2_1
X_24270_ systolic_inst.B_shift\[17\]\[5\] net72 _11333_ B_in\[109\] VGND VGND VPWR
+ VPWR _02207_ sky130_fd_sc_hd__a22o_1
XFILLER_21_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21482_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.A_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\]
+ systolic_inst.A_outs\[3\]\[1\] VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__and4_1
XFILLER_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23221_ net65 _09870_ _09871_ systolic_inst.acc_wires\[1\]\[22\] net109 VGND VGND
+ VPWR VPWR _01896_ sky130_fd_sc_hd__a32o_1
XFILLER_119_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20433_ systolic_inst.A_outs\[5\]\[4\] systolic_inst.B_outs\[5\]\[5\] VGND VGND VPWR
+ VPWR _07369_ sky130_fd_sc_hd__nand2_1
XFILLER_88_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23152_ _09811_ _09812_ VGND VGND VPWR VPWR _09813_ sky130_fd_sc_hd__nor2_1
Xclkload250 clknet_leaf_126_clk VGND VGND VPWR VPWR clkload250/Y sky130_fd_sc_hd__clkinv_2
X_20364_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[7\] _07234_ _07267_
+ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__a211o_1
Xclkload261 clknet_leaf_104_clk VGND VGND VPWR VPWR clkload261/Y sky130_fd_sc_hd__clkinv_4
XFILLER_228_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload272 clknet_leaf_209_clk VGND VGND VPWR VPWR clkload272/Y sky130_fd_sc_hd__clkinv_2
X_22103_ _08852_ _08853_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__or2_1
Xclkload283 clknet_leaf_185_clk VGND VGND VPWR VPWR clkload283/Y sky130_fd_sc_hd__inv_8
XFILLER_175_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23083_ _09753_ VGND VGND VPWR VPWR _09754_ sky130_fd_sc_hd__inv_2
X_27960_ clknet_leaf_168_clk _01758_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload294 clknet_leaf_170_clk VGND VGND VPWR VPWR clkload294/Y sky130_fd_sc_hd__inv_8
XFILLER_175_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20295_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[5\] VGND VGND VPWR
+ VPWR _07235_ sky130_fd_sc_hd__nand2_1
XFILLER_88_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22034_ _08810_ _08809_ systolic_inst.acc_wires\[3\]\[24\] net106 VGND VGND VPWR
+ VPWR _01770_ sky130_fd_sc_hd__a2bb2o_1
X_26911_ clknet_leaf_18_A_in_serial_clk _00709_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27891_ clknet_leaf_38_clk _01689_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29630_ clknet_leaf_10_B_in_serial_clk _03425_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_26842_ clknet_leaf_73_clk _00644_ net144 VGND VGND VPWR VPWR B_in\[114\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29561_ clknet_leaf_15_B_in_serial_clk _03356_ net151 VGND VGND VPWR VPWR deser_B.serial_word\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_26773_ clknet_leaf_96_clk _00575_ net5 VGND VGND VPWR VPWR B_in\[45\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23985_ systolic_inst.B_shift\[12\]\[4\] B_in\[68\] _00008_ VGND VGND VPWR VPWR _10518_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28512_ clknet_leaf_157_clk _02310_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25724_ systolic_inst.acc_wires\[6\]\[8\] C_out\[200\] net47 VGND VGND VPWR VPWR
+ _03026_ sky130_fd_sc_hd__mux2_1
X_22936_ _09612_ _09613_ VGND VGND VPWR VPWR _09615_ sky130_fd_sc_hd__nand2_1
X_29492_ clknet_leaf_281_clk _03290_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[464\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_216_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28443_ clknet_leaf_25_clk _02241_ VGND VGND VPWR VPWR systolic_inst.A_shift\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_189_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25655_ systolic_inst.acc_wires\[4\]\[3\] C_out\[131\] net29 VGND VGND VPWR VPWR
+ _02957_ sky130_fd_sc_hd__mux2_1
X_22867_ _09508_ _09510_ _09507_ VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__a21oi_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire80 net82 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_12
XFILLER_188_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24606_ net110 ser_C.shift_reg\[131\] VGND VGND VPWR VPWR _10773_ sky130_fd_sc_hd__and2_1
X_21818_ _08620_ _08621_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__and2_1
X_28374_ clknet_leaf_33_clk _02172_ VGND VGND VPWR VPWR systolic_inst.A_shift\[19\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25586_ systolic_inst.acc_wires\[1\]\[30\] C_out\[62\] net34 VGND VGND VPWR VPWR
+ _02888_ sky130_fd_sc_hd__mux2_1
X_22798_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[6\] VGND VGND VPWR
+ VPWR _09480_ sky130_fd_sc_hd__nand2_1
XFILLER_197_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27325_ clknet_leaf_330_clk _01123_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_240_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24537_ C_out\[95\] net100 net82 ser_C.shift_reg\[95\] _10738_ VGND VGND VPWR VPWR
+ _02345_ sky130_fd_sc_hd__a221o_1
X_21749_ _08519_ _08554_ systolic_inst.A_outs\[3\]\[7\] VGND VGND VPWR VPWR _08555_
+ sky130_fd_sc_hd__and3b_1
XFILLER_145_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27256_ clknet_leaf_280_clk _01054_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15270_ _12364_ _12365_ VGND VGND VPWR VPWR _12366_ sky130_fd_sc_hd__nand2_1
X_24468_ net114 ser_C.shift_reg\[62\] VGND VGND VPWR VPWR _10704_ sky130_fd_sc_hd__and2_1
XFILLER_156_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26207_ clknet_leaf_15_A_in_serial_clk _00015_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14221_ _11404_ _11407_ VGND VGND VPWR VPWR _11409_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23419_ _10004_ _10043_ VGND VGND VPWR VPWR _10045_ sky130_fd_sc_hd__xnor2_1
X_24399_ C_out\[26\] _11302_ net82 ser_C.shift_reg\[26\] _10669_ VGND VGND VPWR VPWR
+ _02276_ sky130_fd_sc_hd__a221o_1
X_27187_ clknet_leaf_254_clk _00985_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14152_ _11336_ _11343_ VGND VGND VPWR VPWR _11344_ sky130_fd_sc_hd__or2_1
X_26138_ deser_B.serial_word\[93\] deser_B.shift_reg\[93\] net56 VGND VGND VPWR VPWR
+ _03440_ sky130_fd_sc_hd__mux2_1
XFILLER_125_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13103_ systolic_inst.B_outs\[8\]\[7\] VGND VGND VPWR VPWR _11259_ sky130_fd_sc_hd__inv_2
X_14083_ deser_B.shift_reg\[117\] deser_B.shift_reg\[118\] deser_B.receiving VGND
+ VGND VPWR VPWR _00909_ sky130_fd_sc_hd__mux2_1
X_18960_ net66 _06056_ _06057_ systolic_inst.acc_wires\[8\]\[23\] net108 VGND VGND
+ VPWR VPWR _01449_ sky130_fd_sc_hd__a32o_1
X_26069_ deser_B.serial_word\[24\] deser_B.shift_reg\[24\] net56 VGND VGND VPWR VPWR
+ _03371_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _05077_ _05103_ _05104_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__nor3_1
XFILLER_117_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18891_ _05991_ _05996_ _05997_ _05998_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__o211a_1
XFILLER_191_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17842_ _05019_ _05038_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__nor2_1
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_201_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17773_ systolic_inst.acc_wires\[10\]\[28\] systolic_inst.acc_wires\[10\]\[29\] systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__o21ai_1
XFILLER_232_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14985_ _12031_ _12104_ VGND VGND VPWR VPWR _12105_ sky130_fd_sc_hd__nor2_1
XFILLER_208_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19512_ _06540_ _06546_ _06547_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__o21ba_1
XFILLER_43_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16724_ _04043_ _04044_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__xnor2_1
X_13936_ deser_A.serial_word\[97\] deser_A.shift_reg\[97\] net57 VGND VGND VPWR VPWR
+ _00762_ sky130_fd_sc_hd__mux2_1
XFILLER_78_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_193_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19443_ _06492_ _06493_ _06485_ _06489_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__a211o_1
X_16655_ _03969_ _03977_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__xor2_1
X_13867_ deser_A.serial_word\[28\] deser_A.shift_reg\[28\] _00002_ VGND VGND VPWR
+ VPWR _00693_ sky130_fd_sc_hd__mux2_1
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15606_ _12620_ _12628_ _12627_ VGND VGND VPWR VPWR _12662_ sky130_fd_sc_hd__a21bo_1
X_19374_ _06430_ _06431_ _06432_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_18_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16586_ systolic_inst.B_outs\[10\]\[3\] systolic_inst.B_outs\[6\]\[3\] net120 VGND
+ VGND VPWR VPWR _01213_ sky130_fd_sc_hd__mux2_1
XFILLER_90_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13798_ B_in\[105\] deser_B.word_buffer\[105\] _00005_ VGND VGND VPWR VPWR _00635_
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18325_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[20\]
+ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__nand2_1
XFILLER_76_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15537_ _12586_ _12594_ VGND VGND VPWR VPWR _12595_ sky130_fd_sc_hd__xor2_1
XFILLER_176_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_A_in_serial_clk clknet_2_3__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_11_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_176_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18256_ _05429_ _05430_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__nand2_1
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15468_ _12525_ _12526_ _12514_ VGND VGND VPWR VPWR _12528_ sky130_fd_sc_hd__o21bai_1
XFILLER_191_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17207_ systolic_inst.A_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[2\] VGND VGND
+ VPWR VPWR _04470_ sky130_fd_sc_hd__and2_1
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14419_ _11593_ _11601_ VGND VGND VPWR VPWR _11602_ sky130_fd_sc_hd__nand2_1
X_18187_ _05371_ _05372_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__xnor2_1
XFILLER_239_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15399_ net107 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[3\] VGND
+ VGND VPWR VPWR _12462_ sky130_fd_sc_hd__nand2_1
XFILLER_102_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17138_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[25\]
+ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__xor2_2
XFILLER_239_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17069_ _04363_ _04366_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_6_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_146_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20080_ _07056_ _07062_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_146_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_191_Right_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23770_ _10351_ _10374_ _10364_ _10373_ VGND VGND VPWR VPWR _10375_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_211_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20982_ _07817_ _07855_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__and2_1
XFILLER_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22721_ _09404_ _09405_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__nand2_1
XFILLER_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25440_ systolic_inst.cycle_cnt\[1\] systolic_inst.cycle_cnt\[0\] systolic_inst.cycle_cnt\[3\]
+ systolic_inst.cycle_cnt\[2\] VGND VGND VPWR VPWR _11190_ sky130_fd_sc_hd__and4_1
X_22652_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[28\]
+ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__nand2_1
XFILLER_240_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21603_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[5\] VGND VGND VPWR
+ VPWR _08413_ sky130_fd_sc_hd__nand2_1
XFILLER_146_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22583_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[17\]
+ VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__xor2_2
X_25371_ systolic_inst.B_shift\[18\]\[1\] B_in\[49\] net59 VGND VGND VPWR VPWR _11155_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27110_ clknet_leaf_27_B_in_serial_clk _00908_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21534_ _08324_ _08326_ _08325_ VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__a21bo_1
XFILLER_167_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24322_ _10634_ systolic_inst.A_shift\[9\]\[0\] net70 VGND VGND VPWR VPWR _02234_
+ sky130_fd_sc_hd__mux2_1
X_28090_ clknet_leaf_113_clk _01888_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27041_ clknet_leaf_18_B_in_serial_clk _00839_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24253_ systolic_inst.A_shift\[17\]\[4\] net70 net83 systolic_inst.A_shift\[18\]\[4\]
+ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__a22o_1
X_21465_ systolic_inst.A_outs\[3\]\[1\] systolic_inst.A_outs\[2\]\[1\] net122 VGND
+ VGND VPWR VPWR _01715_ sky130_fd_sc_hd__mux2_1
XFILLER_239_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23204_ _09835_ _09856_ VGND VGND VPWR VPWR _09857_ sky130_fd_sc_hd__nor2_1
XFILLER_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20416_ _07352_ _07351_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_131_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24184_ systolic_inst.A_shift\[25\]\[7\] net70 _10505_ systolic_inst.A_shift\[26\]\[7\]
+ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__a22o_1
X_21396_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[21\]
+ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_131_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23135_ _09791_ _09797_ VGND VGND VPWR VPWR _09798_ sky130_fd_sc_hd__nand2_1
XFILLER_218_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20347_ _07263_ _07265_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_92_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28992_ clknet_leaf_58_clk _02790_ VGND VGND VPWR VPWR systolic_inst.A_shift\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_92_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_241_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27943_ clknet_leaf_148_clk _01741_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23066_ net122 _09730_ _09739_ VGND VGND VPWR VPWR _09740_ sky130_fd_sc_hd__and3_1
XFILLER_175_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_241_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20278_ _07217_ _07218_ _07199_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__o21ai_1
XFILLER_115_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_47_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22017_ _08794_ _08795_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__nor2_1
XFILLER_153_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27874_ clknet_leaf_38_clk _01672_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_26__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_26__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_29613_ clknet_leaf_2_B_in_serial_clk _03408_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_26825_ clknet_leaf_71_clk _00627_ net135 VGND VGND VPWR VPWR B_in\[97\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29544_ clknet_leaf_250_clk _03339_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_84_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26756_ clknet_leaf_53_clk _00558_ net143 VGND VGND VPWR VPWR B_in\[28\] sky130_fd_sc_hd__dfrtp_1
X_14770_ _11895_ _11896_ net118 VGND VGND VPWR VPWR _11898_ sky130_fd_sc_hd__o21a_1
X_23968_ _10509_ systolic_inst.B_shift\[9\]\[3\] _11332_ VGND VGND VPWR VPWR _02005_
+ sky130_fd_sc_hd__mux2_1
XFILLER_229_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25707_ systolic_inst.acc_wires\[5\]\[23\] C_out\[183\] net45 VGND VGND VPWR VPWR
+ _03009_ sky130_fd_sc_hd__mux2_1
X_13721_ B_in\[28\] deser_B.word_buffer\[28\] net85 VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__mux2_1
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22919_ _09562_ _09564_ _09563_ VGND VGND VPWR VPWR _09598_ sky130_fd_sc_hd__o21ba_1
X_29475_ clknet_leaf_279_clk _03273_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[447\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26687_ clknet_leaf_30_B_in_serial_clk _00490_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_23899_ _10482_ systolic_inst.B_shift\[13\]\[1\] net72 VGND VGND VPWR VPWR _01963_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16440_ _03805_ _03804_ systolic_inst.acc_wires\[12\]\[11\] net108 VGND VGND VPWR
+ VPWR _01181_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_15_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28426_ clknet_leaf_14_clk _02224_ VGND VGND VPWR VPWR systolic_inst.A_shift\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25638_ systolic_inst.acc_wires\[3\]\[18\] C_out\[114\] net49 VGND VGND VPWR VPWR
+ _02940_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13652_ deser_B.word_buffer\[88\] deser_B.serial_word\[88\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28357_ clknet_leaf_73_clk _02155_ VGND VGND VPWR VPWR systolic_inst.B_shift\[22\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16371_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[12\]\[0\]
+ _03744_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__and4_1
X_25569_ systolic_inst.acc_wires\[1\]\[13\] C_out\[45\] net35 VGND VGND VPWR VPWR
+ _02871_ sky130_fd_sc_hd__mux2_1
X_13583_ deser_B.word_buffer\[19\] deser_B.serial_word\[19\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__mux2_1
XFILLER_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18110_ _05298_ _05297_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__nand2b_1
X_15322_ _12408_ _12409_ VGND VGND VPWR VPWR _12410_ sky130_fd_sc_hd__nand2_1
X_27308_ clknet_leaf_291_clk _01106_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_19090_ _06156_ _06157_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__or2_1
X_28288_ clknet_leaf_54_clk _02086_ VGND VGND VPWR VPWR systolic_inst.B_shift\[19\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18041_ _05196_ _05198_ _05197_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__o21ba_1
XFILLER_240_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15253_ _12347_ _12348_ _12342_ VGND VGND VPWR VPWR _12351_ sky130_fd_sc_hd__or3b_1
X_27239_ clknet_leaf_278_clk _01037_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14204_ _11390_ _11391_ _11386_ VGND VGND VPWR VPWR _11393_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_186_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15184_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[14\]\[6\]
+ VGND VGND VPWR VPWR _12292_ sky130_fd_sc_hd__and2_1
XFILLER_193_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_207_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14135_ systolic_inst.B_outs\[14\]\[3\] systolic_inst.B_outs\[10\]\[3\] net120 VGND
+ VGND VPWR VPWR _00957_ sky130_fd_sc_hd__mux2_1
XFILLER_236_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19992_ _06923_ _06986_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_203_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14066_ deser_B.shift_reg\[100\] deser_B.shift_reg\[101\] net126 VGND VGND VPWR VPWR
+ _00892_ sky130_fd_sc_hd__mux2_1
XFILLER_165_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18943_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[21\]
+ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_199_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18874_ _05968_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__nand2_1
XFILLER_80_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17825_ _05021_ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__nand2_1
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17756_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[27\]
+ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14968_ _12047_ _12049_ _12088_ VGND VGND VPWR VPWR _12089_ sky130_fd_sc_hd__a21o_1
X_16707_ systolic_inst.A_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[4\]
+ systolic_inst.B_outs\[11\]\[3\] VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__a22oi_1
XFILLER_207_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13919_ deser_A.serial_word\[80\] deser_A.shift_reg\[80\] net57 VGND VGND VPWR VPWR
+ _00745_ sky130_fd_sc_hd__mux2_1
X_17687_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[16\]
+ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14899_ _11991_ _12020_ VGND VGND VPWR VPWR _12022_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19426_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[7\]\[4\]
+ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__and2_1
X_16638_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[4\] _03962_
+ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__a21bo_1
XFILLER_222_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19357_ _06415_ _06416_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__nand2b_1
XFILLER_241_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16569_ _03912_ _03915_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18308_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[17\]
+ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__xor2_1
XFILLER_241_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19288_ systolic_inst.A_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[5\] systolic_inst.B_outs\[7\]\[6\]
+ systolic_inst.B_outs\[7\]\[7\] VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__and4b_1
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18239_ _05408_ _05412_ _05414_ _05415_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__o211ai_2
XFILLER_175_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21250_ _08113_ _08114_ _08115_ _08104_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__a211oi_1
XFILLER_102_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap120 systolic_inst.ce_local VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_12
X_20201_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[28\]
+ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__or2_1
Xmax_cap131 net133 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_16
XFILLER_132_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap153 net5 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_16
XFILLER_137_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21181_ _08047_ _08048_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__xor2_1
XFILLER_102_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20132_ _07105_ _07107_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20063_ net68 _07047_ _07048_ systolic_inst.acc_wires\[6\]\[7\] net106 VGND VGND
+ VPWR VPWR _01561_ sky130_fd_sc_hd__a32o_1
X_24940_ net111 ser_C.shift_reg\[298\] VGND VGND VPWR VPWR _10940_ sky130_fd_sc_hd__and2_1
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24871_ C_out\[262\] net101 net73 ser_C.shift_reg\[262\] _10905_ VGND VGND VPWR VPWR
+ _02512_ sky130_fd_sc_hd__a221o_1
X_26610_ clknet_leaf_15_B_in_serial_clk _00413_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_23822_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[20\]
+ VGND VGND VPWR VPWR _10419_ sky130_fd_sc_hd__xor2_1
XFILLER_2_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27590_ clknet_leaf_223_clk _01388_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_A_in_serial_clk clknet_2_2__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_6_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26541_ clknet_leaf_20_A_in_serial_clk _00344_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23753_ _10356_ _10358_ _10360_ systolic_inst.acc_wires\[0\]\[9\] _11258_ VGND VGND
+ VPWR VPWR _01939_ sky130_fd_sc_hd__a32o_1
X_20965_ _07804_ _07837_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__xor2_1
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22704_ systolic_inst.A_outs\[1\]\[1\] systolic_inst.B_outs\[1\]\[2\] systolic_inst.B_outs\[1\]\[3\]
+ systolic_inst.A_outs\[1\]\[0\] VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__a22oi_1
X_29260_ clknet_leaf_198_clk _03058_ net146 VGND VGND VPWR VPWR C_out\[232\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26472_ clknet_leaf_14_A_in_serial_clk _00275_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23684_ _10299_ _10301_ VGND VGND VPWR VPWR _10303_ sky130_fd_sc_hd__xnor2_2
X_20896_ net108 _07772_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28211_ clknet_leaf_97_clk _02009_ VGND VGND VPWR VPWR systolic_inst.B_shift\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_81_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25423_ systolic_inst.A_shift\[1\]\[3\] A_in\[3\] net59 VGND VGND VPWR VPWR _11181_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22635_ _09341_ _09343_ _09345_ VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__o21ai_1
X_29191_ clknet_leaf_218_clk _02989_ net140 VGND VGND VPWR VPWR C_out\[163\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_230_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28142_ clknet_leaf_123_clk _01940_ net153 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_230_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22566_ _09286_ _09288_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_133_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25354_ net112 ser_C.shift_reg\[505\] VGND VGND VPWR VPWR _11147_ sky130_fd_sc_hd__and2_1
XFILLER_194_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21517_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.A_outs\[3\]\[4\] VGND VGND VPWR
+ VPWR _08330_ sky130_fd_sc_hd__nand2_1
XFILLER_155_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24305_ systolic_inst.A_shift\[11\]\[0\] A_in\[40\] net59 VGND VGND VPWR VPWR _10626_
+ sky130_fd_sc_hd__mux2_1
X_28073_ clknet_leaf_118_clk _01871_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22497_ _09229_ VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__inv_2
XFILLER_186_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25285_ ser_C.parallel_data\[469\] net102 net74 ser_C.shift_reg\[469\] _11112_ VGND
+ VGND VPWR VPWR _02719_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27024_ clknet_leaf_19_B_in_serial_clk _00822_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21448_ _08283_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__inv_2
X_24236_ _10603_ systolic_inst.A_shift\[18\]\[1\] net70 VGND VGND VPWR VPWR _02179_
+ sky130_fd_sc_hd__mux2_1
XFILLER_119_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24167_ systolic_inst.A_shift\[28\]\[7\] A_in\[103\] net59 VGND VGND VPWR VPWR _10585_
+ sky130_fd_sc_hd__mux2_1
X_21379_ _08224_ _08225_ _08223_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__a21o_1
XFILLER_163_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23118_ net64 _09782_ _09783_ systolic_inst.acc_wires\[1\]\[7\] net109 VGND VGND
+ VPWR VPWR _01881_ sky130_fd_sc_hd__a32o_1
XFILLER_123_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24098_ _10558_ systolic_inst.B_shift\[19\]\[4\] net71 VGND VGND VPWR VPWR _02086_
+ sky130_fd_sc_hd__mux2_1
X_28975_ clknet_leaf_63_clk _02773_ VGND VGND VPWR VPWR systolic_inst.A_shift\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23049_ _09655_ _09699_ _09698_ VGND VGND VPWR VPWR _09724_ sky130_fd_sc_hd__o21a_1
X_27926_ clknet_leaf_132_clk _01724_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_15940_ _12958_ _12961_ VGND VGND VPWR VPWR _12962_ sky130_fd_sc_hd__xor2_1
XFILLER_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15871_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[18\]
+ VGND VGND VPWR VPWR _12903_ sky130_fd_sc_hd__or2_1
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27857_ clknet_leaf_34_clk _01655_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_188_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _04850_ _04851_ _04852_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__and3_1
X_26808_ clknet_leaf_83_clk _00610_ net144 VGND VGND VPWR VPWR B_in\[80\] sky130_fd_sc_hd__dfrtp_1
X_14822_ _11943_ _11946_ VGND VGND VPWR VPWR _11947_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18590_ _05718_ _05717_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_237_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27788_ clknet_leaf_307_clk _01586_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_188_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29527_ clknet_leaf_264_clk _03325_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17541_ _04791_ _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__nor2_1
X_26739_ clknet_leaf_98_clk _00541_ net5 VGND VGND VPWR VPWR B_in\[11\] sky130_fd_sc_hd__dfrtp_1
X_14753_ systolic_inst.B_outs\[13\]\[5\] systolic_inst.B_outs\[9\]\[5\] net117 VGND
+ VGND VPWR VPWR _01023_ sky130_fd_sc_hd__mux2_1
XFILLER_229_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13704_ B_in\[11\] deser_B.word_buffer\[11\] net84 VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__mux2_1
XFILLER_205_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29458_ clknet_leaf_329_clk _03256_ net136 VGND VGND VPWR VPWR C_out\[430\] sky130_fd_sc_hd__dfrtp_1
X_17472_ _04685_ _04687_ _04724_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__nand3_1
X_14684_ _11838_ VGND VGND VPWR VPWR _11839_ sky130_fd_sc_hd__inv_2
XFILLER_225_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19211_ _06238_ _06273_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__and2_1
X_28409_ clknet_leaf_82_clk _02207_ VGND VGND VPWR VPWR systolic_inst.B_shift\[17\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16423_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[12\]\[8\]
+ _03786_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__a211o_1
XFILLER_232_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13635_ deser_B.word_buffer\[71\] deser_B.serial_word\[71\] net123 VGND VGND VPWR
+ VPWR _00472_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29389_ clknet_leaf_242_clk _03187_ net145 VGND VGND VPWR VPWR C_out\[361\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19142_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[5\] VGND VGND VPWR
+ VPWR _06208_ sky130_fd_sc_hd__nand2_1
XFILLER_201_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16354_ _03731_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__or2_1
XFILLER_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13566_ deser_B.word_buffer\[2\] deser_B.serial_word\[2\] net124 VGND VGND VPWR VPWR
+ _00403_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_188_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15305_ _11712_ _12394_ _12395_ systolic_inst.acc_wires\[14\]\[23\] net107 VGND VGND
+ VPWR VPWR _01065_ sky130_fd_sc_hd__a32o_1
XFILLER_201_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19073_ _06123_ _06139_ _06140_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__and3_1
XFILLER_146_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16285_ _03663_ _03664_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__xnor2_1
X_13497_ deser_A.shift_reg\[61\] deser_A.shift_reg\[62\] net130 VGND VGND VPWR VPWR
+ _00334_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_184_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18024_ _05213_ _05215_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__nand2_1
XFILLER_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15236_ _12331_ _12335_ VGND VGND VPWR VPWR _12337_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15167_ _12268_ _12272_ _12275_ _12276_ VGND VGND VPWR VPWR _12278_ sky130_fd_sc_hd__o211a_1
XFILLER_113_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14118_ systolic_inst.A_shift\[21\]\[2\] net71 _11333_ A_in\[90\] VGND VGND VPWR
+ VPWR _00940_ sky130_fd_sc_hd__a22o_1
XFILLER_236_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19975_ _06922_ _06970_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15098_ _12146_ _12213_ VGND VGND VPWR VPWR _12215_ sky130_fd_sc_hd__or2_1
XFILLER_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14049_ deser_B.shift_reg\[83\] deser_B.shift_reg\[84\] net125 VGND VGND VPWR VPWR
+ _00875_ sky130_fd_sc_hd__mux2_1
X_18926_ _06019_ _06021_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__nand2_1
XFILLER_136_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18857_ _05962_ _05964_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__nand2_1
XFILLER_227_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_230_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_230_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_209_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17808_ systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[1\] VGND VGND VPWR
+ VPWR _05007_ sky130_fd_sc_hd__nand2_1
X_18788_ _05856_ _05861_ _05885_ _05887_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__o31a_1
XFILLER_95_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17739_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[24\]
+ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_137_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20750_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[20\]
+ VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__or2_1
XFILLER_91_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19409_ _06464_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__inv_2
XFILLER_17_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20681_ _07596_ _07598_ _07600_ systolic_inst.acc_wires\[5\]\[9\] net109 VGND VGND
+ VPWR VPWR _01627_ sky130_fd_sc_hd__a32o_1
XFILLER_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22420_ _09128_ _09131_ _09158_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__or3_1
XFILLER_17_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22351_ _09091_ _09092_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__nand2_1
XFILLER_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_297_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_297_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_143_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21302_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[4\]\[8\]
+ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__or2_1
XFILLER_136_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25070_ net112 ser_C.shift_reg\[363\] VGND VGND VPWR VPWR _11005_ sky130_fd_sc_hd__and2_1
X_22282_ systolic_inst.B_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[5\] systolic_inst.A_outs\[2\]\[6\]
+ systolic_inst.B_outs\[2\]\[3\] VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__a22oi_1
XFILLER_164_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24021_ systolic_inst.B_shift\[6\]\[4\] _11332_ net83 systolic_inst.B_shift\[10\]\[4\]
+ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__a22o_1
XFILLER_219_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21233_ _08069_ _08076_ _08099_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__or3_1
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21164_ _08031_ _08032_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__nor2_1
XFILLER_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_B_in_serial_clk clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_13_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_132_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20115_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[15\]
+ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__nor2_1
X_28760_ clknet_leaf_217_clk _02558_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[308\]
+ sky130_fd_sc_hd__dfrtp_1
X_21095_ systolic_inst.A_outs\[4\]\[3\] _07852_ _07964_ VGND VGND VPWR VPWR _07966_
+ sky130_fd_sc_hd__o21a_1
X_25972_ systolic_inst.acc_wires\[14\]\[0\] ser_C.parallel_data\[448\] net24 VGND
+ VGND VPWR VPWR _03274_ sky130_fd_sc_hd__mux2_1
XFILLER_63_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27711_ clknet_leaf_193_clk _01509_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20046_ _07027_ _07028_ _07026_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__a21bo_1
X_24923_ C_out\[288\] net102 net74 ser_C.shift_reg\[288\] _10931_ VGND VGND VPWR VPWR
+ _02538_ sky130_fd_sc_hd__a221o_1
X_28691_ clknet_leaf_192_clk _02489_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[239\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_221_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_221_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27642_ clknet_leaf_311_clk _01440_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24854_ net113 ser_C.shift_reg\[255\] VGND VGND VPWR VPWR _10897_ sky130_fd_sc_hd__and2_1
XFILLER_234_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23805_ _11258_ systolic_inst.acc_wires\[0\]\[16\] _10403_ _10405_ VGND VGND VPWR
+ VPWR _01946_ sky130_fd_sc_hd__a22o_1
XFILLER_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27573_ clknet_leaf_304_clk _01371_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24785_ C_out\[219\] net98 net78 ser_C.shift_reg\[219\] _10862_ VGND VGND VPWR VPWR
+ _02469_ sky130_fd_sc_hd__a221o_1
X_21997_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[19\]
+ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__xnor2_1
XFILLER_215_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29312_ clknet_leaf_302_clk _03110_ net141 VGND VGND VPWR VPWR C_out\[284\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26524_ clknet_leaf_4_A_in_serial_clk _00327_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_232_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23736_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[0\]\[7\]
+ VGND VGND VPWR VPWR _10346_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_232_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20948_ _07786_ _07788_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__nand2_1
XFILLER_214_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29243_ clknet_leaf_187_clk _03041_ net148 VGND VGND VPWR VPWR C_out\[215\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26455_ clknet_leaf_346_clk _00262_ net132 VGND VGND VPWR VPWR A_in\[123\] sky130_fd_sc_hd__dfrtp_1
X_23667_ _10283_ _10285_ VGND VGND VPWR VPWR _10286_ sky130_fd_sc_hd__nand2_1
XFILLER_201_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _07754_ _07755_ VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__nor2_1
XFILLER_186_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25406_ _11172_ systolic_inst.A_shift\[1\]\[2\] net71 VGND VGND VPWR VPWR _02780_
+ sky130_fd_sc_hd__mux2_1
X_13420_ net130 deser_A.bit_idx\[0\] _11308_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__o21ba_1
X_22618_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[23\]
+ VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__xnor2_1
XFILLER_197_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29174_ clknet_leaf_41_clk _02972_ net142 VGND VGND VPWR VPWR C_out\[146\] sky130_fd_sc_hd__dfrtp_1
X_26386_ clknet_leaf_15_clk _00193_ net134 VGND VGND VPWR VPWR A_in\[54\] sky130_fd_sc_hd__dfrtp_1
XFILLER_201_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23598_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[11\] _10219_ systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__mux2_1
XFILLER_224_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28125_ clknet_leaf_50_clk _01923_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_288_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_288_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_31_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25337_ ser_C.parallel_data\[495\] net97 net77 ser_C.shift_reg\[495\] _11138_ VGND
+ VGND VPWR VPWR _02745_ sky130_fd_sc_hd__a221o_1
X_13351_ A_in\[60\] deser_A.word_buffer\[60\] net91 VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__mux2_1
X_22549_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[2\]\[12\]
+ VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28056_ clknet_leaf_125_clk _01854_ net144 VGND VGND VPWR VPWR systolic_inst.B_outs\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16070_ _13064_ _13065_ VGND VGND VPWR VPWR _13066_ sky130_fd_sc_hd__or2_1
XFILLER_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25268_ net111 ser_C.shift_reg\[462\] VGND VGND VPWR VPWR _11104_ sky130_fd_sc_hd__and2_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13282_ deser_A.word_buffer\[120\] deser_A.serial_word\[120\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__mux2_1
XFILLER_136_950 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27007_ clknet_leaf_16_B_in_serial_clk _00805_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_170_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15021_ systolic_inst.A_outs\[14\]\[6\] _12109_ _12110_ _12075_ VGND VGND VPWR VPWR
+ _12140_ sky130_fd_sc_hd__o2bb2a_1
X_24219_ systolic_inst.A_shift\[20\]\[1\] A_in\[73\] net59 VGND VGND VPWR VPWR _10595_
+ sky130_fd_sc_hd__mux2_1
X_25199_ C_out\[426\] net101 net73 ser_C.shift_reg\[426\] _11069_ VGND VGND VPWR VPWR
+ _02676_ sky130_fd_sc_hd__a221o_1
XFILLER_108_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19760_ _06727_ _06761_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16972_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[11\]\[1\]
+ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__and2_1
X_28958_ clknet_leaf_258_clk _02756_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[506\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15923_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[26\]
+ VGND VGND VPWR VPWR _12947_ sky130_fd_sc_hd__or2_1
XFILLER_42_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18711_ systolic_inst.B_outs\[8\]\[6\] systolic_inst.A_outs\[8\]\[6\] _11259_ systolic_inst.A_outs\[8\]\[5\]
+ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_231_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19691_ systolic_inst.A_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[2\] systolic_inst.B_outs\[6\]\[3\]
+ systolic_inst.B_outs\[6\]\[4\] VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__and4_1
X_27909_ clknet_leaf_44_clk _01707_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_118_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28889_ clknet_leaf_287_clk _02687_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[437\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_212_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_212_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18642_ systolic_inst.A_outs\[8\]\[6\] _05768_ _05767_ VGND VGND VPWR VPWR _05769_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_231_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _12887_ _12888_ VGND VGND VPWR VPWR _12889_ sky130_fd_sc_hd__or2_1
XFILLER_37_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14805_ _11911_ _11927_ _11929_ VGND VGND VPWR VPWR _11931_ sky130_fd_sc_hd__and3_1
X_18573_ _05700_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__nor2_1
X_15785_ _12826_ _12827_ _12828_ VGND VGND VPWR VPWR _12830_ sky130_fd_sc_hd__and3_1
XFILLER_206_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17524_ _04744_ _04747_ _04775_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__o21ai_1
X_14736_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[31\]
+ VGND VGND VPWR VPWR _11883_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17455_ _04602_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__or2_1
XFILLER_162_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14667_ _11821_ _11823_ _11824_ VGND VGND VPWR VPWR _11825_ sky130_fd_sc_hd__or3_1
XFILLER_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16406_ _03774_ _03776_ _03769_ _03772_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_215_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13618_ deser_B.word_buffer\[54\] deser_B.serial_word\[54\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__mux2_1
XFILLER_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17386_ _04640_ _04641_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__or2_1
XFILLER_158_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14598_ net105 systolic_inst.acc_wires\[15\]\[10\] net69 _11765_ VGND VGND VPWR VPWR
+ _00988_ sky130_fd_sc_hd__a22o_1
XFILLER_242_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19125_ _06168_ _06190_ _06191_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_279_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_279_clk
+ sky130_fd_sc_hd__clkbuf_8
X_16337_ systolic_inst.B_outs\[12\]\[5\] systolic_inst.B_outs\[12\]\[6\] systolic_inst.A_outs\[12\]\[7\]
+ _03715_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__a31o_1
X_13549_ deser_A.shift_reg\[113\] deser_A.shift_reg\[114\] net129 VGND VGND VPWR VPWR
+ _00386_ sky130_fd_sc_hd__mux2_1
XFILLER_146_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19056_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[2\] VGND VGND VPWR
+ VPWR _06125_ sky130_fd_sc_hd__and2_1
XFILLER_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16268_ _03590_ _03649_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18007_ _05197_ _05198_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__nor2_1
X_15219_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[14\]\[11\]
+ VGND VGND VPWR VPWR _12322_ sky130_fd_sc_hd__nand2_1
XFILLER_103_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16199_ _03582_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__inv_2
XFILLER_12_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19958_ _06951_ _06952_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_162_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_162_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18909_ _06012_ _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__and2_1
XFILLER_214_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19889_ _06885_ _06886_ _06884_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__o21ai_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_203_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_203_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_210_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21920_ _08712_ _08711_ systolic_inst.acc_wires\[3\]\[8\] net106 VGND VGND VPWR VPWR
+ _01754_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21851_ _08584_ _08653_ VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20802_ _07696_ _07700_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__nor2_1
X_24570_ net113 ser_C.shift_reg\[113\] VGND VGND VPWR VPWR _10755_ sky130_fd_sc_hd__and2_1
X_21782_ systolic_inst.B_outs\[3\]\[6\] systolic_inst.A_outs\[3\]\[6\] _11274_ systolic_inst.A_outs\[3\]\[5\]
+ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_230_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23521_ _10114_ _10116_ _10115_ VGND VGND VPWR VPWR _10144_ sky130_fd_sc_hd__o21ba_1
XFILLER_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20733_ net106 systolic_inst.acc_wires\[5\]\[16\] _07643_ _07645_ VGND VGND VPWR
+ VPWR _01634_ sky130_fd_sc_hd__a22o_1
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26240_ clknet_leaf_17_A_in_serial_clk _00048_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23452_ _10073_ _10076_ VGND VGND VPWR VPWR _10077_ sky130_fd_sc_hd__xnor2_1
X_20664_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[5\]\[7\]
+ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_119_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22403_ _09142_ _09143_ VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__nor2_1
XFILLER_108_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23383_ _10008_ _10009_ VGND VGND VPWR VPWR _10010_ sky130_fd_sc_hd__and2b_1
X_26171_ deser_B.serial_word\[126\] deser_B.shift_reg\[126\] net56 VGND VGND VPWR
+ VPWR _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20595_ _07435_ _07524_ VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25122_ net110 ser_C.shift_reg\[389\] VGND VGND VPWR VPWR _11031_ sky130_fd_sc_hd__and2_1
X_22334_ _09058_ _09076_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__xor2_1
XFILLER_192_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22265_ _09009_ _09008_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__nand2b_1
X_25053_ C_out\[353\] net97 net77 ser_C.shift_reg\[353\] _10996_ VGND VGND VPWR VPWR
+ _02603_ sky130_fd_sc_hd__a221o_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24004_ _10527_ systolic_inst.B_shift\[5\]\[5\] _11332_ VGND VGND VPWR VPWR _02023_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21216_ _08049_ _08051_ _08082_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_225_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22196_ _08941_ _08942_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__nor2_1
XFILLER_133_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21147_ _08016_ _08015_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__nand2b_1
X_28812_ clknet_leaf_243_clk _02610_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[360\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_221_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_221_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28743_ clknet_leaf_297_clk _02541_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_116_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25955_ systolic_inst.acc_wires\[13\]\[15\] C_out\[431\] net20 VGND VGND VPWR VPWR
+ _03257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21078_ _07907_ _07910_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__nor2_1
XFILLER_8_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20029_ net68 _07017_ _07019_ systolic_inst.acc_wires\[6\]\[2\] net106 VGND VGND
+ VPWR VPWR _01556_ sky130_fd_sc_hd__a32o_1
XFILLER_46_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24906_ net110 ser_C.shift_reg\[281\] VGND VGND VPWR VPWR _10923_ sky130_fd_sc_hd__and2_1
XFILLER_98_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28674_ clknet_leaf_184_clk _02472_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_150_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25886_ systolic_inst.acc_wires\[11\]\[10\] C_out\[362\] net39 VGND VGND VPWR VPWR
+ _03188_ sky130_fd_sc_hd__mux2_1
XFILLER_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27625_ clknet_leaf_316_clk _01423_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_24837_ C_out\[245\] net98 net78 ser_C.shift_reg\[245\] _10888_ VGND VGND VPWR VPWR
+ _02495_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_219_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15570_ _12626_ _12625_ VGND VGND VPWR VPWR _12627_ sky130_fd_sc_hd__nand2b_1
X_27556_ clknet_leaf_304_clk _01354_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_226_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24768_ net113 ser_C.shift_reg\[212\] VGND VGND VPWR VPWR _10854_ sky130_fd_sc_hd__and2_1
XFILLER_148_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14521_ _11622_ _11684_ _11683_ VGND VGND VPWR VPWR _11700_ sky130_fd_sc_hd__o21ba_1
X_26507_ clknet_leaf_17_A_in_serial_clk _00310_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_23719_ _10328_ _10329_ _10330_ VGND VGND VPWR VPWR _10332_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_29_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27487_ clknet_leaf_228_clk _01285_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_24699_ C_out\[176\] net100 net80 ser_C.shift_reg\[176\] _10819_ VGND VGND VPWR VPWR
+ _02426_ sky130_fd_sc_hd__a221o_1
XFILLER_186_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29226_ clknet_leaf_211_clk _03024_ net147 VGND VGND VPWR VPWR C_out\[198\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17240_ _04483_ _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__nand2_1
XFILLER_30_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26438_ clknet_leaf_1_clk _00245_ net134 VGND VGND VPWR VPWR A_in\[106\] sky130_fd_sc_hd__dfrtp_1
X_14452_ _11632_ _11633_ VGND VGND VPWR VPWR _11634_ sky130_fd_sc_hd__nand2_1
XFILLER_74_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13403_ A_in\[112\] deser_A.word_buffer\[112\] net96 VGND VGND VPWR VPWR _00251_
+ sky130_fd_sc_hd__mux2_1
X_17171_ _04450_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__nand2_1
X_29157_ clknet_leaf_311_clk _02955_ net142 VGND VGND VPWR VPWR C_out\[129\] sky130_fd_sc_hd__dfrtp_1
X_14383_ _11566_ _11565_ VGND VGND VPWR VPWR _11567_ sky130_fd_sc_hd__nand2b_1
X_26369_ clknet_leaf_27_clk _00176_ net137 VGND VGND VPWR VPWR A_in\[37\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_8_B_in_serial_clk clknet_2_2__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_8_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_200_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_210_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28108_ clknet_leaf_56_clk _01906_ net143 VGND VGND VPWR VPWR systolic_inst.A_outs\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_16122_ _13084_ _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__and2b_1
XFILLER_122_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13334_ A_in\[43\] deser_A.word_buffer\[43\] net95 VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__mux2_1
X_29088_ clknet_leaf_157_clk _02886_ net151 VGND VGND VPWR VPWR C_out\[60\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_210_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28039_ clknet_leaf_162_clk _01837_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16053_ _13026_ _13049_ VGND VGND VPWR VPWR _13050_ sky130_fd_sc_hd__nand2b_1
XFILLER_182_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13265_ deser_A.word_buffer\[103\] deser_A.serial_word\[103\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__mux2_1
XFILLER_108_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15004_ _12122_ _12123_ VGND VGND VPWR VPWR _12124_ sky130_fd_sc_hd__nand2b_1
XFILLER_237_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13196_ deser_A.word_buffer\[34\] deser_A.serial_word\[34\] net127 VGND VGND VPWR
+ VPWR _00044_ sky130_fd_sc_hd__mux2_1
XFILLER_9_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19812_ _06811_ _06812_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__nor2_1
XFILLER_155_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19743_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[6\]
+ systolic_inst.A_outs\[6\]\[7\] VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__nand4_1
XFILLER_42_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16955_ _04269_ _04268_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__nand2b_1
XFILLER_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15906_ _12925_ _12929_ _12932_ VGND VGND VPWR VPWR _12933_ sky130_fd_sc_hd__nand3_1
X_19674_ _06677_ _06678_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__nand2b_1
XFILLER_77_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16886_ _04201_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__nor2_1
XFILLER_133_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15837_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[13\]\[12\]
+ _12871_ _12873_ VGND VGND VPWR VPWR _12874_ sky130_fd_sc_hd__a211o_1
X_18625_ _05699_ _05716_ _05715_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__o21ba_1
XFILLER_18_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15768_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[13\]\[3\]
+ VGND VGND VPWR VPWR _12815_ sky130_fd_sc_hd__or2_1
X_18556_ _05656_ _05684_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14719_ _11867_ _11868_ VGND VGND VPWR VPWR _11869_ sky130_fd_sc_hd__nand2_1
X_17507_ _04709_ _04759_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__and2b_1
X_18487_ _05589_ _05591_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15699_ _12718_ _12721_ _12750_ VGND VGND VPWR VPWR _12752_ sky130_fd_sc_hd__or3_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17438_ _04674_ _04692_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_155_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_15 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 net153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_37 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17369_ _04571_ _04586_ _04585_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__o21a_1
XFILLER_242_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19108_ _06147_ _06174_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_168_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20380_ _07316_ _07317_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_168_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19039_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[2\] _06109_ VGND
+ VGND VPWR VPWR _06110_ sky130_fd_sc_hd__nand3_1
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22050_ _08823_ _08822_ systolic_inst.acc_wires\[3\]\[27\] net106 VGND VGND VPWR
+ VPWR _01773_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21001_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[5\] _07846_ _07845_
+ systolic_inst.B_outs\[4\]\[5\] VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__a32o_1
XFILLER_99_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_7__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_87_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25740_ systolic_inst.acc_wires\[6\]\[24\] C_out\[216\] net44 VGND VGND VPWR VPWR
+ _03042_ sky130_fd_sc_hd__mux2_1
XFILLER_96_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22952_ systolic_inst.A_outs\[1\]\[5\] systolic_inst.B_outs\[1\]\[6\] _11277_ systolic_inst.A_outs\[1\]\[4\]
+ VGND VGND VPWR VPWR _09630_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_108_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap17 net18 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_4
XFILLER_216_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21903_ _08698_ VGND VGND VPWR VPWR _08699_ sky130_fd_sc_hd__inv_2
Xmax_cap28 net29 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_4
X_25671_ systolic_inst.acc_wires\[4\]\[19\] C_out\[147\] net32 VGND VGND VPWR VPWR
+ _02973_ sky130_fd_sc_hd__mux2_1
XFILLER_16_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22883_ systolic_inst.A_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[6\]
+ systolic_inst.B_outs\[1\]\[7\] VGND VGND VPWR VPWR _09563_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_69_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap39 net40 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_8
XFILLER_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27410_ clknet_leaf_226_clk _01208_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_24622_ net110 ser_C.shift_reg\[139\] VGND VGND VPWR VPWR _10781_ sky130_fd_sc_hd__and2_1
X_21834_ _08607_ _08612_ _08637_ VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__o21ai_1
X_28390_ clknet_leaf_33_clk _02188_ VGND VGND VPWR VPWR systolic_inst.A_shift\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_203_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27341_ clknet_leaf_342_clk _01139_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24553_ C_out\[103\] net99 net79 ser_C.shift_reg\[103\] _10746_ VGND VGND VPWR VPWR
+ _02353_ sky130_fd_sc_hd__a221o_1
XFILLER_169_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21765_ _08517_ _08535_ _08534_ VGND VGND VPWR VPWR _08571_ sky130_fd_sc_hd__o21a_1
XFILLER_169_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23504_ _10118_ _10127_ VGND VGND VPWR VPWR _10128_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_117_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20716_ _07624_ _07630_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__nand2_1
X_27272_ clknet_leaf_266_clk _01070_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_24484_ net112 ser_C.shift_reg\[70\] VGND VGND VPWR VPWR _10712_ sky130_fd_sc_hd__and2_1
XFILLER_12_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21696_ _08503_ _08502_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__nand2b_1
X_29011_ clknet_leaf_103_clk _02809_ net151 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_211_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26223_ clknet_leaf_10_A_in_serial_clk _00031_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23435_ _10019_ _10021_ _10059_ _10060_ VGND VGND VPWR VPWR _10061_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_78_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20647_ _07568_ _07569_ _07570_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__and3_1
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_227_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26154_ deser_B.serial_word\[109\] deser_B.shift_reg\[109\] _00001_ VGND VGND VPWR
+ VPWR _03456_ sky130_fd_sc_hd__mux2_1
XFILLER_137_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20578_ _07509_ _07508_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__and2b_1
X_23366_ _09972_ _09992_ VGND VGND VPWR VPWR _09993_ sky130_fd_sc_hd__nand2_1
XFILLER_137_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25105_ C_out\[379\] net99 net79 ser_C.shift_reg\[379\] _11022_ VGND VGND VPWR VPWR
+ _02629_ sky130_fd_sc_hd__a221o_1
X_22317_ systolic_inst.B_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[7\]
+ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__and3_1
XFILLER_165_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_223_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26085_ deser_B.serial_word\[40\] deser_B.shift_reg\[40\] net55 VGND VGND VPWR VPWR
+ _03387_ sky130_fd_sc_hd__mux2_1
XFILLER_191_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23297_ _09919_ _09927_ VGND VGND VPWR VPWR _09928_ sky130_fd_sc_hd__xor2_1
XFILLER_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25036_ net112 ser_C.shift_reg\[346\] VGND VGND VPWR VPWR _10988_ sky130_fd_sc_hd__and2_1
XFILLER_3_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22248_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[6\] VGND VGND VPWR
+ VPWR _08993_ sky130_fd_sc_hd__nand2_1
XFILLER_180_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22179_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[4\] _08923_ _08924_
+ VGND VGND VPWR VPWR _08926_ sky130_fd_sc_hd__a22o_1
XFILLER_239_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26987_ clknet_leaf_30_A_in_serial_clk _00785_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16740_ _04054_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__xnor2_1
X_25938_ systolic_inst.acc_wires\[12\]\[30\] C_out\[414\] net21 VGND VGND VPWR VPWR
+ _03240_ sky130_fd_sc_hd__mux2_1
X_13952_ deser_A.serial_word\[113\] deser_A.shift_reg\[113\] net57 VGND VGND VPWR
+ VPWR _00778_ sky130_fd_sc_hd__mux2_1
X_28726_ clknet_leaf_314_clk _02524_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[274\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28657_ clknet_leaf_204_clk _02455_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[205\]
+ sky130_fd_sc_hd__dfrtp_1
X_16671_ _03966_ _03993_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__xor2_1
XFILLER_189_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25869_ systolic_inst.acc_wires\[10\]\[25\] C_out\[345\] net11 VGND VGND VPWR VPWR
+ _03171_ sky130_fd_sc_hd__mux2_1
XFILLER_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13883_ deser_A.serial_word\[44\] deser_A.shift_reg\[44\] net58 VGND VGND VPWR VPWR
+ _00709_ sky130_fd_sc_hd__mux2_1
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15622_ _12674_ _12676_ VGND VGND VPWR VPWR _12678_ sky130_fd_sc_hd__nand2_2
X_18410_ systolic_inst.A_outs\[8\]\[7\] systolic_inst.A_shift\[16\]\[7\] net121 VGND
+ VGND VPWR VPWR _01401_ sky130_fd_sc_hd__mux2_1
X_27608_ clknet_leaf_204_clk _01406_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_19390_ _06396_ _06426_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__nor2_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28588_ clknet_leaf_307_clk _02386_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[136\]
+ sky130_fd_sc_hd__dfrtp_1
X_18341_ _05502_ _05503_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__and2_1
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15553_ _12573_ _12602_ _12601_ VGND VGND VPWR VPWR _12610_ sky130_fd_sc_hd__a21o_1
X_27539_ clknet_leaf_311_clk _01337_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_226_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14504_ _11657_ _11659_ _11682_ VGND VGND VPWR VPWR _11684_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_212_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18272_ _05441_ _05444_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_212_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _11272_ _12542_ VGND VGND VPWR VPWR _12543_ sky130_fd_sc_hd__xnor2_1
XFILLER_230_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17223_ net107 _04484_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__nor2_1
X_29209_ clknet_leaf_181_clk _03007_ net146 VGND VGND VPWR VPWR C_out\[181\] sky130_fd_sc_hd__dfrtp_1
XFILLER_147_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[11\] _11617_ net118
+ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17154_ systolic_inst.acc_wires\[11\]\[26\] systolic_inst.acc_wires\[11\]\[27\] systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__o21a_1
XFILLER_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14366_ _11549_ _11550_ VGND VGND VPWR VPWR _11551_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16105_ systolic_inst.A_outs\[12\]\[2\] systolic_inst.B_outs\[12\]\[5\] VGND VGND
+ VPWR VPWR _13100_ sky130_fd_sc_hd__nand2_1
XFILLER_196_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13317_ A_in\[26\] deser_A.word_buffer\[26\] net91 VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__mux2_1
XFILLER_13_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17085_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[17\]
+ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14297_ systolic_inst.B_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[4\]
+ systolic_inst.A_outs\[15\]\[5\] VGND VGND VPWR VPWR _11483_ sky130_fd_sc_hd__and4_1
XFILLER_143_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16036_ _13011_ _13032_ VGND VGND VPWR VPWR _13033_ sky130_fd_sc_hd__nand2_1
XFILLER_131_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13248_ deser_A.word_buffer\[86\] deser_A.serial_word\[86\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__mux2_1
XFILLER_83_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13179_ deser_A.word_buffer\[17\] deser_A.serial_word\[17\] net128 VGND VGND VPWR
+ VPWR _00027_ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17987_ _05178_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__or2_2
XFILLER_111_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19726_ _06724_ _06725_ _06727_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__or3_1
XFILLER_133_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1092 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16938_ systolic_inst.B_outs\[11\]\[5\] systolic_inst.A_outs\[11\]\[7\] _04231_ _04230_
+ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__a31o_1
XFILLER_226_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19657_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[3\] _06662_ net119
+ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16869_ _04185_ _04186_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__nor2_1
XFILLER_25_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18608_ systolic_inst.B_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[5\] systolic_inst.A_outs\[8\]\[6\]
+ systolic_inst.B_outs\[8\]\[3\] VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__a22oi_1
XFILLER_203_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19588_ systolic_inst.acc_wires\[7\]\[26\] systolic_inst.acc_wires\[7\]\[27\] systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_157_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18539_ _05665_ _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21550_ _08353_ _08361_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20501_ _07364_ _07434_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__xnor2_4
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21481_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[0\] _08297_
+ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__a21o_1
XFILLER_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23220_ _09867_ _09868_ _09869_ VGND VGND VPWR VPWR _09871_ sky130_fd_sc_hd__or3_1
X_20432_ _07364_ _07367_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload240 clknet_leaf_91_clk VGND VGND VPWR VPWR clkload240/Y sky130_fd_sc_hd__clkinvlp_4
X_23151_ _09808_ _09809_ _09810_ VGND VGND VPWR VPWR _09812_ sky130_fd_sc_hd__a21oi_1
XFILLER_162_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20363_ systolic_inst.B_outs\[5\]\[5\] _07267_ systolic_inst.B_outs\[5\]\[7\] systolic_inst.A_outs\[5\]\[0\]
+ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__o211ai_1
XFILLER_179_1374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload251 clknet_leaf_127_clk VGND VGND VPWR VPWR clkload251/X sky130_fd_sc_hd__clkbuf_4
Xclkload262 clknet_leaf_105_clk VGND VGND VPWR VPWR clkload262/Y sky130_fd_sc_hd__clkinvlp_4
X_22102_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[1\]
+ systolic_inst.A_outs\[2\]\[2\] VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__and4_1
XFILLER_161_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload273 clknet_leaf_210_clk VGND VGND VPWR VPWR clkload273/Y sky130_fd_sc_hd__clkinv_4
X_23082_ _09749_ _09750_ _09751_ VGND VGND VPWR VPWR _09753_ sky130_fd_sc_hd__and3_1
Xclkload284 clknet_leaf_188_clk VGND VGND VPWR VPWR clkload284/Y sky130_fd_sc_hd__inv_4
Xclkload295 clknet_leaf_171_clk VGND VGND VPWR VPWR clkload295/Y sky130_fd_sc_hd__inv_6
X_20294_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[5\] VGND VGND VPWR
+ VPWR _07234_ sky130_fd_sc_hd__and2_1
X_22033_ _08805_ _08808_ net60 VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__a21o_1
XFILLER_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26910_ clknet_leaf_18_A_in_serial_clk _00708_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_27890_ clknet_leaf_38_clk _01688_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26841_ clknet_leaf_73_clk _00643_ net144 VGND VGND VPWR VPWR B_in\[113\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29560_ clknet_leaf_15_B_in_serial_clk _03355_ net152 VGND VGND VPWR VPWR deser_B.serial_word\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26772_ clknet_leaf_96_clk _00574_ net5 VGND VGND VPWR VPWR B_in\[44\] sky130_fd_sc_hd__dfrtp_1
X_23984_ _10517_ systolic_inst.B_shift\[8\]\[3\] net72 VGND VGND VPWR VPWR _02013_
+ sky130_fd_sc_hd__mux2_1
XFILLER_169_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28511_ clknet_leaf_157_clk _02309_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25723_ systolic_inst.acc_wires\[6\]\[7\] C_out\[199\] net47 VGND VGND VPWR VPWR
+ _03025_ sky130_fd_sc_hd__mux2_1
XFILLER_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22935_ _09612_ _09613_ VGND VGND VPWR VPWR _09614_ sky130_fd_sc_hd__or2_2
X_29491_ clknet_leaf_282_clk _03289_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_216_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28442_ clknet_leaf_35_clk _02240_ VGND VGND VPWR VPWR systolic_inst.A_shift\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25654_ systolic_inst.acc_wires\[4\]\[2\] C_out\[130\] net29 VGND VGND VPWR VPWR
+ _02956_ sky130_fd_sc_hd__mux2_1
X_22866_ _09544_ _09545_ VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24605_ C_out\[129\] net103 net75 ser_C.shift_reg\[129\] _10772_ VGND VGND VPWR VPWR
+ _02379_ sky130_fd_sc_hd__a221o_1
X_21817_ _08588_ _08591_ _08619_ VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__or3_1
X_28373_ clknet_leaf_27_clk _02171_ VGND VGND VPWR VPWR systolic_inst.A_shift\[19\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25585_ systolic_inst.acc_wires\[1\]\[29\] C_out\[61\] net52 VGND VGND VPWR VPWR
+ _02887_ sky130_fd_sc_hd__mux2_1
X_22797_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.A_outs\[1\]\[7\] VGND VGND VPWR
+ VPWR _09479_ sky130_fd_sc_hd__nand2_1
XFILLER_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27324_ clknet_leaf_330_clk _01122_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_24536_ net114 ser_C.shift_reg\[96\] VGND VGND VPWR VPWR _10738_ sky130_fd_sc_hd__and2_1
X_21748_ systolic_inst.B_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\] VGND VGND VPWR
+ VPWR _08554_ sky130_fd_sc_hd__or2_1
XFILLER_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27255_ clknet_leaf_278_clk _01053_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_24467_ C_out\[60\] net100 net82 ser_C.shift_reg\[60\] _10703_ VGND VGND VPWR VPWR
+ _02310_ sky130_fd_sc_hd__a221o_1
XFILLER_200_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21679_ systolic_inst.B_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[5\]
+ systolic_inst.A_outs\[3\]\[6\] VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__and4_1
XFILLER_156_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26206_ clknet_leaf_15_A_in_serial_clk _00014_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14220_ _11407_ _11404_ VGND VGND VPWR VPWR _11408_ sky130_fd_sc_hd__and2b_1
X_23418_ _10004_ _10043_ VGND VGND VPWR VPWR _10044_ sky130_fd_sc_hd__nand2_1
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27186_ clknet_leaf_253_clk _00984_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24398_ net114 ser_C.shift_reg\[27\] VGND VGND VPWR VPWR _10669_ sky130_fd_sc_hd__and2_1
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26137_ deser_B.serial_word\[92\] deser_B.shift_reg\[92\] net56 VGND VGND VPWR VPWR
+ _03439_ sky130_fd_sc_hd__mux2_1
XFILLER_153_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14151_ _11341_ _11342_ VGND VGND VPWR VPWR _11343_ sky130_fd_sc_hd__nor2_1
X_23349_ _09974_ _09975_ _09949_ VGND VGND VPWR VPWR _09977_ sky130_fd_sc_hd__o21a_1
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13102_ net116 VGND VGND VPWR VPWR _11258_ sky130_fd_sc_hd__clkinv_16
X_14082_ deser_B.shift_reg\[116\] deser_B.shift_reg\[117\] deser_B.receiving VGND
+ VGND VPWR VPWR _00908_ sky130_fd_sc_hd__mux2_1
X_26068_ deser_B.serial_word\[23\] deser_B.shift_reg\[23\] net55 VGND VGND VPWR VPWR
+ _03370_ sky130_fd_sc_hd__mux2_1
XFILLER_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25019_ C_out\[336\] net97 net80 ser_C.shift_reg\[336\] _10979_ VGND VGND VPWR VPWR
+ _02586_ sky130_fd_sc_hd__a221o_1
X_17910_ _05103_ _05104_ _05077_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__o21ai_1
XFILLER_121_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18890_ _05989_ _05995_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__or2_1
XFILLER_117_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17841_ _05016_ _05037_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14984_ _12075_ _12076_ _12077_ VGND VGND VPWR VPWR _12104_ sky130_fd_sc_hd__o21ba_1
X_17772_ net105 systolic_inst.acc_wires\[10\]\[29\] net62 _04991_ VGND VGND VPWR VPWR
+ _01327_ sky130_fd_sc_hd__a22o_1
XFILLER_208_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19511_ _06528_ _06536_ _06550_ _06551_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__o31a_1
XFILLER_130_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28709_ clknet_leaf_325_clk _02507_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[257\]
+ sky130_fd_sc_hd__dfrtp_1
X_13935_ deser_A.serial_word\[96\] deser_A.shift_reg\[96\] net57 VGND VGND VPWR VPWR
+ _00761_ sky130_fd_sc_hd__mux2_1
X_16723_ _04044_ _04043_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__nand2b_1
X_29689_ clknet_leaf_8_clk _03484_ VGND VGND VPWR VPWR systolic_inst.A_shift\[30\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_193_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_193_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19442_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[7\]\[6\]
+ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__or2_1
X_16654_ _03969_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__nor2_1
XFILLER_90_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13866_ deser_A.serial_word\[27\] deser_A.shift_reg\[27\] net58 VGND VGND VPWR VPWR
+ _00692_ sky130_fd_sc_hd__mux2_1
XFILLER_35_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15605_ _12659_ _12660_ VGND VGND VPWR VPWR _12661_ sky130_fd_sc_hd__nand2_1
XFILLER_234_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19373_ _11261_ systolic_inst.A_outs\[7\]\[7\] _06380_ _06404_ VGND VGND VPWR VPWR
+ _06432_ sky130_fd_sc_hd__o211a_1
X_16585_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.B_outs\[6\]\[2\] net120 VGND
+ VGND VPWR VPWR _01212_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13797_ B_in\[104\] deser_B.word_buffer\[104\] _00005_ VGND VGND VPWR VPWR _00634_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_241_Right_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18324_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[20\]
+ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__or2_1
XFILLER_37_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15536_ _12591_ _12592_ VGND VGND VPWR VPWR _12594_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_152_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18255_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[9\]\[10\]
+ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__nand2_1
XFILLER_163_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15467_ _12525_ _12526_ _12514_ VGND VGND VPWR VPWR _12527_ sky130_fd_sc_hd__or3b_1
XFILLER_198_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17206_ _04460_ _04467_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__xnor2_1
X_14418_ _11598_ _11599_ VGND VGND VPWR VPWR _11601_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18186_ _05289_ _05351_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__xnor2_1
X_15398_ _12446_ _12448_ _12459_ VGND VGND VPWR VPWR _12461_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17137_ _04425_ _04424_ systolic_inst.acc_wires\[11\]\[24\] net105 VGND VGND VPWR
+ VPWR _01258_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_156_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14349_ systolic_inst.A_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[5\] _11491_ _11490_
+ VGND VGND VPWR VPWR _11534_ sky130_fd_sc_hd__a31o_1
XFILLER_128_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17068_ _04363_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__nand2_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16019_ _13009_ _13015_ VGND VGND VPWR VPWR _13017_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_146_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19709_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[3\] _06696_ _06695_
+ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__a31o_1
XFILLER_226_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20981_ _07849_ _07854_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22720_ systolic_inst.A_outs\[1\]\[1\] systolic_inst.B_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\]
+ systolic_inst.A_outs\[1\]\[0\] VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__a22o_1
XFILLER_168_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22651_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[28\]
+ VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__or2_1
XFILLER_213_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21602_ _08375_ _08411_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25370_ _11154_ systolic_inst.B_shift\[14\]\[0\] _11332_ VGND VGND VPWR VPWR _02762_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22582_ net109 systolic_inst.acc_wires\[2\]\[16\] _09300_ _09302_ VGND VGND VPWR
+ VPWR _01826_ sky130_fd_sc_hd__a22o_1
XFILLER_240_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24321_ systolic_inst.A_shift\[10\]\[0\] A_in\[32\] net59 VGND VGND VPWR VPWR _10634_
+ sky130_fd_sc_hd__mux2_1
X_21533_ _08311_ _08332_ _08334_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27040_ clknet_leaf_12_B_in_serial_clk _00838_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24252_ systolic_inst.A_shift\[17\]\[3\] net70 net83 systolic_inst.A_shift\[18\]\[3\]
+ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__a22o_1
X_21464_ systolic_inst.A_outs\[3\]\[0\] systolic_inst.A_outs\[2\]\[0\] net122 VGND
+ VGND VPWR VPWR _01714_ sky130_fd_sc_hd__mux2_1
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23203_ _09836_ _09841_ _09846_ _09850_ VGND VGND VPWR VPWR _09856_ sky130_fd_sc_hd__or4_1
X_20415_ _07310_ _07312_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_96_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21395_ net63 _08238_ _08239_ systolic_inst.acc_wires\[4\]\[20\] _11258_ VGND VGND
+ VPWR VPWR _01702_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_131_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24183_ systolic_inst.A_shift\[25\]\[6\] net70 _10505_ systolic_inst.A_shift\[26\]\[6\]
+ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__a22o_1
XFILLER_190_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23134_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[1\]\[9\]
+ _09792_ VGND VGND VPWR VPWR _09797_ sky130_fd_sc_hd__a21oi_1
XFILLER_190_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20346_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[6\] _07284_ net120
+ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28991_ clknet_leaf_58_clk _02789_ VGND VGND VPWR VPWR systolic_inst.A_shift\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_92_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_241_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27942_ clknet_leaf_148_clk _01740_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_23065_ _09735_ _09738_ VGND VGND VPWR VPWR _09739_ sky130_fd_sc_hd__xnor2_1
X_20277_ _07214_ _07216_ _07197_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_241_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22016_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[22\]
+ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__and2_1
XFILLER_62_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27873_ clknet_leaf_38_clk _01671_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29612_ clknet_leaf_33_B_in_serial_clk _03407_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_26824_ clknet_leaf_71_clk _00626_ net135 VGND VGND VPWR VPWR B_in\[96\] sky130_fd_sc_hd__dfrtp_1
XFILLER_153_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26755_ clknet_leaf_56_clk _00557_ net137 VGND VGND VPWR VPWR B_in\[27\] sky130_fd_sc_hd__dfrtp_1
X_29543_ clknet_leaf_250_clk _03338_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_23967_ systolic_inst.B_shift\[13\]\[3\] B_in\[43\] _00008_ VGND VGND VPWR VPWR _10509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25706_ systolic_inst.acc_wires\[5\]\[22\] C_out\[182\] net45 VGND VGND VPWR VPWR
+ _03008_ sky130_fd_sc_hd__mux2_1
X_13720_ B_in\[27\] deser_B.word_buffer\[27\] net85 VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__mux2_1
X_22918_ _09593_ _09596_ VGND VGND VPWR VPWR _09597_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26686_ clknet_leaf_29_B_in_serial_clk _00489_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_29474_ clknet_leaf_285_clk _03272_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23898_ systolic_inst.B_shift\[17\]\[1\] B_in\[73\] _00008_ VGND VGND VPWR VPWR _10482_
+ sky130_fd_sc_hd__mux2_1
XFILLER_216_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25637_ systolic_inst.acc_wires\[3\]\[17\] C_out\[113\] net49 VGND VGND VPWR VPWR
+ _02939_ sky130_fd_sc_hd__mux2_1
X_13651_ deser_B.word_buffer\[87\] deser_B.serial_word\[87\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28425_ clknet_leaf_22_clk _02223_ VGND VGND VPWR VPWR systolic_inst.A_shift\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22849_ _09489_ _09529_ VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28356_ clknet_leaf_84_clk _02154_ VGND VGND VPWR VPWR systolic_inst.B_shift\[22\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16370_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[12\]\[1\]
+ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__or2_1
X_25568_ systolic_inst.acc_wires\[1\]\[12\] C_out\[44\] net35 VGND VGND VPWR VPWR
+ _02870_ sky130_fd_sc_hd__mux2_1
X_13582_ deser_B.word_buffer\[18\] deser_B.serial_word\[18\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__mux2_1
XFILLER_213_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27307_ clknet_leaf_329_clk _01105_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15321_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[26\]
+ VGND VGND VPWR VPWR _12409_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24519_ C_out\[86\] net100 net82 ser_C.shift_reg\[86\] _10729_ VGND VGND VPWR VPWR
+ _02336_ sky130_fd_sc_hd__a221o_1
X_28287_ clknet_leaf_56_clk _02085_ VGND VGND VPWR VPWR systolic_inst.B_shift\[19\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25499_ _11228_ _11229_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__nor2_1
XFILLER_8_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18040_ _05227_ _05230_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15252_ net67 _12349_ _12350_ systolic_inst.acc_wires\[14\]\[15\] net107 VGND VGND
+ VPWR VPWR _01057_ sky130_fd_sc_hd__a32o_1
X_27238_ clknet_leaf_278_clk _01036_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_200_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ _11386_ _11390_ _11391_ VGND VGND VPWR VPWR _11392_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_186_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15183_ _11712_ _12289_ _12291_ systolic_inst.acc_wires\[14\]\[5\] net107 VGND VGND
+ VPWR VPWR _01047_ sky130_fd_sc_hd__a32o_1
X_27169_ clknet_leaf_253_clk _00967_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_186_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_207_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14134_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.B_outs\[10\]\[2\] net120 VGND
+ VGND VPWR VPWR _00956_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_207_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19991_ _06984_ _06985_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__nor2_1
XFILLER_235_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14065_ deser_B.shift_reg\[99\] deser_B.shift_reg\[100\] net126 VGND VGND VPWR VPWR
+ _00891_ sky130_fd_sc_hd__mux2_1
XFILLER_165_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18942_ net66 _06041_ _06042_ systolic_inst.acc_wires\[8\]\[20\] net108 VGND VGND
+ VPWR VPWR _01446_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_203_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18873_ _05974_ _05979_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__nor2_1
XFILLER_121_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17824_ _05019_ _05020_ _05009_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__a21o_1
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14967_ _12079_ _12087_ VGND VGND VPWR VPWR _12088_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17755_ net105 systolic_inst.acc_wires\[10\]\[26\] net69 _04977_ VGND VGND VPWR VPWR
+ _01324_ sky130_fd_sc_hd__a22o_1
XFILLER_208_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16706_ systolic_inst.B_outs\[11\]\[3\] systolic_inst.A_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\]
+ systolic_inst.A_outs\[11\]\[4\] VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__and4_1
X_13918_ deser_A.serial_word\[79\] deser_A.shift_reg\[79\] net57 VGND VGND VPWR VPWR
+ _00744_ sky130_fd_sc_hd__mux2_1
X_14898_ _11991_ _12020_ VGND VGND VPWR VPWR _12021_ sky130_fd_sc_hd__nand2b_1
X_17686_ _04917_ _04918_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__and2_1
XFILLER_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19425_ net62 _06476_ _06478_ systolic_inst.acc_wires\[7\]\[3\] net105 VGND VGND
+ VPWR VPWR _01493_ sky130_fd_sc_hd__a32o_1
X_13849_ deser_A.serial_word\[10\] deser_A.shift_reg\[10\] net58 VGND VGND VPWR VPWR
+ _00675_ sky130_fd_sc_hd__mux2_1
XFILLER_23_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16637_ net105 _03960_ _03961_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__or3_1
XFILLER_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19356_ _06348_ _06384_ _06383_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__a21bo_1
X_16568_ _03913_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__nand2_1
XFILLER_222_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18307_ net106 systolic_inst.acc_wires\[9\]\[16\] _05473_ _05475_ VGND VGND VPWR
+ VPWR _01378_ sky130_fd_sc_hd__a22o_1
XFILLER_52_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15519_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[7\]
+ VGND VGND VPWR VPWR _12577_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_171_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19287_ systolic_inst.B_outs\[7\]\[5\] systolic_inst.A_outs\[7\]\[6\] VGND VGND VPWR
+ VPWR _06349_ sky130_fd_sc_hd__nand2_1
X_16499_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[19\]
+ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18238_ _05414_ _05415_ _05408_ _05412_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_21_B_in_serial_clk clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_21_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_102_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18169_ _05354_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__nor2_1
XFILLER_172_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap110 net7 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_12
Xmax_cap121 systolic_inst.ce_local VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_12
X_20200_ _07149_ _07151_ _07163_ _07164_ _07157_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__a311oi_4
XFILLER_85_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21180_ _08048_ _08047_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__nand2b_1
XFILLER_239_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20131_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[16\]
+ _07103_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__a21oi_1
XFILLER_132_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20062_ _07044_ _07045_ _07046_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__nand3_1
XFILLER_98_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24870_ net110 ser_C.shift_reg\[263\] VGND VGND VPWR VPWR _10905_ sky130_fd_sc_hd__and2_1
XFILLER_61_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23821_ _11258_ systolic_inst.acc_wires\[0\]\[19\] net64 _10418_ VGND VGND VPWR VPWR
+ _01949_ sky130_fd_sc_hd__a22o_1
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26540_ clknet_leaf_21_A_in_serial_clk _00343_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_23752_ _11713_ _10359_ VGND VGND VPWR VPWR _10360_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20964_ _07804_ _07837_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__or2_1
XFILLER_226_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22703_ net122 _09388_ _09389_ _09382_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_85_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26471_ clknet_leaf_13_A_in_serial_clk _00274_ net143 VGND VGND VPWR VPWR deser_A.shift_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_23683_ _10299_ _10301_ VGND VGND VPWR VPWR _10302_ sky130_fd_sc_hd__nor2_1
XFILLER_242_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20895_ _07748_ _07770_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__and2_1
X_28210_ clknet_leaf_97_clk _02008_ VGND VGND VPWR VPWR systolic_inst.B_shift\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25422_ _11180_ systolic_inst.A_shift\[0\]\[2\] net71 VGND VGND VPWR VPWR _02788_
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22634_ _09341_ _09343_ _09345_ VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__or3_1
XFILLER_213_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29190_ clknet_leaf_306_clk _02988_ net140 VGND VGND VPWR VPWR C_out\[162\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28141_ clknet_leaf_124_clk _01939_ net153 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_181_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25353_ ser_C.parallel_data\[503\] net98 net78 ser_C.shift_reg\[503\] _11146_ VGND
+ VGND VPWR VPWR _02753_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_230_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22565_ _09281_ _09287_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__nand2_1
XFILLER_167_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_230_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24304_ _10625_ systolic_inst.A_shift\[11\]\[7\] net71 VGND VGND VPWR VPWR _02225_
+ sky130_fd_sc_hd__mux2_1
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28072_ clknet_leaf_119_clk _01870_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_21516_ _08328_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__inv_2
X_25284_ net111 ser_C.shift_reg\[470\] VGND VGND VPWR VPWR _11112_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22496_ _09225_ _09226_ _09227_ VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__and3_1
XFILLER_155_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27023_ clknet_leaf_19_B_in_serial_clk _00821_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24235_ systolic_inst.A_shift\[19\]\[1\] A_in\[65\] net59 VGND VGND VPWR VPWR _10603_
+ sky130_fd_sc_hd__mux2_1
X_21447_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[29\]
+ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__xor2_1
XFILLER_33_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24166_ _10584_ systolic_inst.A_shift\[27\]\[6\] net70 VGND VGND VPWR VPWR _02128_
+ sky130_fd_sc_hd__mux2_1
X_21378_ _08216_ _08218_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__nand2_1
XFILLER_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23117_ _09779_ _09780_ _09781_ VGND VGND VPWR VPWR _09783_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_9_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20329_ systolic_inst.A_outs\[5\]\[1\] systolic_inst.B_outs\[5\]\[5\] systolic_inst.B_outs\[5\]\[6\]
+ systolic_inst.A_outs\[5\]\[0\] VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24097_ systolic_inst.B_shift\[23\]\[4\] B_in\[60\] _00008_ VGND VGND VPWR VPWR _10558_
+ sky130_fd_sc_hd__mux2_1
X_28974_ clknet_leaf_60_clk _02772_ VGND VGND VPWR VPWR systolic_inst.A_shift\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23048_ _09655_ _09722_ VGND VGND VPWR VPWR _09723_ sky130_fd_sc_hd__xnor2_1
X_27925_ clknet_leaf_131_clk _01723_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15870_ net108 systolic_inst.acc_wires\[13\]\[17\] net67 _12902_ VGND VGND VPWR VPWR
+ _01123_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27856_ clknet_leaf_35_clk _01654_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_34_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14821_ _11944_ _11945_ VGND VGND VPWR VPWR _11946_ sky130_fd_sc_hd__and2b_1
X_26807_ clknet_leaf_83_clk _00609_ net144 VGND VGND VPWR VPWR B_in\[79\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27787_ clknet_leaf_184_clk _01585_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24999_ C_out\[326\] net97 net80 ser_C.shift_reg\[326\] _10969_ VGND VGND VPWR VPWR
+ _02576_ sky130_fd_sc_hd__a221o_1
XFILLER_91_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29526_ clknet_leaf_264_clk _03324_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[498\]
+ sky130_fd_sc_hd__dfrtp_1
X_14752_ systolic_inst.B_outs\[13\]\[4\] systolic_inst.B_outs\[9\]\[4\] net115 VGND
+ VGND VPWR VPWR _01022_ sky130_fd_sc_hd__mux2_1
X_17540_ _04758_ _04760_ _04790_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__o21a_1
X_26738_ clknet_leaf_94_clk _00540_ net152 VGND VGND VPWR VPWR B_in\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13703_ B_in\[10\] deser_B.word_buffer\[10\] net84 VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _04685_ _04687_ _04724_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__a21o_1
X_26669_ clknet_leaf_8_B_in_serial_clk _00472_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_29457_ clknet_leaf_329_clk _03255_ net136 VGND VGND VPWR VPWR C_out\[429\] sky130_fd_sc_hd__dfrtp_1
X_14683_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[23\]
+ VGND VGND VPWR VPWR _11838_ sky130_fd_sc_hd__xor2_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19210_ _06238_ _06273_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__nor2_1
XFILLER_242_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28408_ clknet_leaf_82_clk _02206_ VGND VGND VPWR VPWR systolic_inst.B_shift\[17\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13634_ deser_B.word_buffer\[70\] deser_B.serial_word\[70\] net123 VGND VGND VPWR
+ VPWR _00471_ sky130_fd_sc_hd__mux2_1
X_16422_ _03788_ _03789_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__nor2_1
XFILLER_32_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29388_ clknet_leaf_243_clk _03186_ net145 VGND VGND VPWR VPWR C_out\[360\] sky130_fd_sc_hd__dfrtp_1
X_19141_ _06171_ _06206_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__xnor2_1
X_16353_ _03681_ _03686_ _03709_ _03710_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__o31a_1
XFILLER_201_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13565_ deser_B.word_buffer\[1\] deser_B.serial_word\[1\] net124 VGND VGND VPWR VPWR
+ _00402_ sky130_fd_sc_hd__mux2_1
X_28339_ clknet_leaf_342_clk _02137_ VGND VGND VPWR VPWR systolic_inst.A_shift\[26\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15304_ _12386_ _12390_ _12393_ VGND VGND VPWR VPWR _12395_ sky130_fd_sc_hd__a21o_1
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19072_ _06139_ _06140_ _06123_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__a21oi_1
X_16284_ systolic_inst.B_outs\[12\]\[5\] systolic_inst.A_outs\[12\]\[7\] _03663_ VGND
+ VGND VPWR VPWR _03665_ sky130_fd_sc_hd__and3_1
X_13496_ deser_A.shift_reg\[60\] deser_A.shift_reg\[61\] net130 VGND VGND VPWR VPWR
+ _00333_ sky130_fd_sc_hd__mux2_1
XFILLER_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15235_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[14\]\[12\]
+ _12333_ _12335_ VGND VGND VPWR VPWR _12336_ sky130_fd_sc_hd__a211o_1
X_18023_ _05214_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__inv_2
XFILLER_201_1153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15166_ _12275_ _12276_ _12268_ _12272_ VGND VGND VPWR VPWR _12277_ sky130_fd_sc_hd__a211o_1
XFILLER_236_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14117_ systolic_inst.A_shift\[21\]\[1\] net71 _11333_ A_in\[89\] VGND VGND VPWR
+ VPWR _00939_ sky130_fd_sc_hd__a22o_1
X_19974_ _06968_ _06969_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__nor2_1
X_15097_ _12146_ _12213_ VGND VGND VPWR VPWR _12214_ sky130_fd_sc_hd__nand2_1
X_14048_ deser_B.shift_reg\[82\] deser_B.shift_reg\[83\] net125 VGND VGND VPWR VPWR
+ _00874_ sky130_fd_sc_hd__mux2_1
XFILLER_45_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18925_ systolic_inst.acc_wires\[8\]\[16\] systolic_inst.acc_wires\[8\]\[17\] systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__o21ai_1
XFILLER_192_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18856_ _05966_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__and2b_1
XFILLER_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17807_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[1\] _05004_
+ _05006_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__a22o_1
XFILLER_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18787_ _05907_ _05908_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__xnor2_1
X_15999_ _12996_ _12997_ VGND VGND VPWR VPWR _12998_ sky130_fd_sc_hd__nand2_1
XFILLER_94_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17738_ _04942_ _04962_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__nor2_1
XFILLER_224_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_207_Left_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17669_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[10\]\[14\]
+ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__or2_1
XFILLER_224_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19408_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[7\]\[0\]
+ _06462_ _06463_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__and4_1
XFILLER_1_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20680_ _11713_ _07599_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19339_ _06335_ _06339_ _06369_ _06368_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__o31a_1
XFILLER_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22350_ _08985_ _09090_ VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__nand2_1
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21301_ net63 _08157_ _08158_ systolic_inst.acc_wires\[4\]\[7\] net108 VGND VGND
+ VPWR VPWR _01689_ sky130_fd_sc_hd__a32o_1
X_22281_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[7\] VGND VGND VPWR
+ VPWR _09025_ sky130_fd_sc_hd__nand2_4
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24020_ systolic_inst.B_shift\[6\]\[3\] _11332_ net83 systolic_inst.B_shift\[10\]\[3\]
+ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__a22o_1
XFILLER_145_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21232_ _08097_ _08098_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__and2_1
XFILLER_219_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21163_ systolic_inst.A_outs\[4\]\[5\] _07852_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__nor2_1
XFILLER_176_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20114_ net68 _07091_ _07092_ systolic_inst.acc_wires\[6\]\[14\] net106 VGND VGND
+ VPWR VPWR _01568_ sky130_fd_sc_hd__a32o_1
XFILLER_49_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21094_ systolic_inst.A_outs\[4\]\[3\] _07852_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__nor2_1
XFILLER_115_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25971_ systolic_inst.acc_wires\[13\]\[31\] ser_C.parallel_data\[447\] net26 VGND
+ VGND VPWR VPWR _03273_ sky130_fd_sc_hd__mux2_1
XFILLER_59_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27710_ clknet_leaf_194_clk _01508_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_20045_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[6\]\[5\]
+ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_126_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24922_ net111 ser_C.shift_reg\[289\] VGND VGND VPWR VPWR _10931_ sky130_fd_sc_hd__and2_1
X_28690_ clknet_leaf_192_clk _02488_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24853_ C_out\[253\] net98 net78 ser_C.shift_reg\[253\] _10896_ VGND VGND VPWR VPWR
+ _02503_ sky130_fd_sc_hd__a221o_1
XFILLER_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27641_ clknet_leaf_316_clk _01439_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23804_ _11713_ _10404_ VGND VGND VPWR VPWR _10405_ sky130_fd_sc_hd__nor2_1
XFILLER_100_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27572_ clknet_leaf_304_clk _01370_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24784_ net113 ser_C.shift_reg\[220\] VGND VGND VPWR VPWR _10862_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_83_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21996_ net65 _08777_ _08778_ systolic_inst.acc_wires\[3\]\[18\] net109 VGND VGND
+ VPWR VPWR _01764_ sky130_fd_sc_hd__a32o_1
XFILLER_96_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29311_ clknet_leaf_302_clk _03109_ net141 VGND VGND VPWR VPWR C_out\[283\] sky130_fd_sc_hd__dfrtp_1
X_26523_ clknet_leaf_4_A_in_serial_clk _00326_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23735_ net63 _10343_ _10345_ systolic_inst.acc_wires\[0\]\[6\] _11258_ VGND VGND
+ VPWR VPWR _01936_ sky130_fd_sc_hd__a32o_1
XFILLER_27_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20947_ _07809_ _07821_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_232_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_232_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29242_ clknet_leaf_176_clk _03040_ net148 VGND VGND VPWR VPWR C_out\[214\] sky130_fd_sc_hd__dfrtp_1
X_26454_ clknet_leaf_346_clk _00261_ net132 VGND VGND VPWR VPWR A_in\[122\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23666_ _10154_ _10195_ _10222_ VGND VGND VPWR VPWR _10285_ sky130_fd_sc_hd__or3b_1
XFILLER_241_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20878_ _07741_ _07753_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__and2_1
XFILLER_224_1120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25405_ systolic_inst.A_shift\[2\]\[2\] A_in\[10\] net59 VGND VGND VPWR VPWR _11172_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22617_ net65 _09330_ _09331_ systolic_inst.acc_wires\[2\]\[22\] net109 VGND VGND
+ VPWR VPWR _01832_ sky130_fd_sc_hd__a32o_1
X_29173_ clknet_leaf_41_clk _02971_ net141 VGND VGND VPWR VPWR C_out\[145\] sky130_fd_sc_hd__dfrtp_1
XFILLER_70_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26385_ clknet_leaf_12_clk _00192_ net132 VGND VGND VPWR VPWR A_in\[53\] sky130_fd_sc_hd__dfrtp_1
X_23597_ _10184_ _10218_ VGND VGND VPWR VPWR _10219_ sky130_fd_sc_hd__xnor2_1
XFILLER_197_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28124_ clknet_leaf_124_clk _01922_ net144 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25336_ net112 ser_C.shift_reg\[496\] VGND VGND VPWR VPWR _11138_ sky130_fd_sc_hd__and2_1
X_13350_ A_in\[59\] deser_A.word_buffer\[59\] net91 VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__mux2_1
XFILLER_224_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22548_ _09258_ _09264_ _09266_ VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__o21a_1
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28055_ clknet_leaf_125_clk _01853_ net144 VGND VGND VPWR VPWR systolic_inst.B_outs\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_127_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25267_ ser_C.parallel_data\[460\] net102 net74 ser_C.shift_reg\[460\] _11103_ VGND
+ VGND VPWR VPWR _02710_ sky130_fd_sc_hd__a221o_1
X_13281_ deser_A.word_buffer\[119\] deser_A.serial_word\[119\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__mux2_1
X_22479_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[2\]\[2\]
+ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__or2_1
X_27006_ clknet_leaf_15_B_in_serial_clk _00804_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_170_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15020_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[10\] _12139_ net118
+ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__mux2_1
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24218_ _10594_ systolic_inst.A_shift\[19\]\[0\] net70 VGND VGND VPWR VPWR _02170_
+ sky130_fd_sc_hd__mux2_1
X_25198_ net111 ser_C.shift_reg\[427\] VGND VGND VPWR VPWR _11069_ sky130_fd_sc_hd__and2_1
XFILLER_151_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24149_ systolic_inst.A_shift\[29\]\[6\] A_in\[110\] net59 VGND VGND VPWR VPWR _10576_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28957_ clknet_leaf_258_clk _02755_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[505\]
+ sky130_fd_sc_hd__dfrtp_1
X_16971_ net118 _04282_ _04283_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18710_ _05833_ _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__nand2_2
X_27908_ clknet_leaf_43_clk _01706_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_15922_ net67 _12945_ _12946_ systolic_inst.acc_wires\[13\]\[25\] net107 VGND VGND
+ VPWR VPWR _01131_ sky130_fd_sc_hd__a32o_1
X_19690_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[3\] VGND VGND VPWR
+ VPWR _06694_ sky130_fd_sc_hd__nand2_1
X_28888_ clknet_leaf_287_clk _02686_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[436\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_231_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18641_ systolic_inst.B_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[7\]
+ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_177_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27839_ clknet_leaf_205_clk _01637_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_15853_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[15\]
+ VGND VGND VPWR VPWR _12888_ sky130_fd_sc_hd__and2_1
XFILLER_76_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_177_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14804_ _11927_ _11929_ _11911_ VGND VGND VPWR VPWR _11930_ sky130_fd_sc_hd__a21oi_1
XFILLER_206_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18572_ systolic_inst.B_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[5\]
+ systolic_inst.B_outs\[8\]\[3\] VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__a22oi_1
XFILLER_218_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15784_ _12826_ _12827_ _12828_ VGND VGND VPWR VPWR _12829_ sky130_fd_sc_hd__a21o_1
XFILLER_217_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29509_ clknet_leaf_265_clk _03307_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[481\]
+ sky130_fd_sc_hd__dfrtp_1
X_17523_ _04746_ _04773_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14735_ net69 _11881_ _11882_ systolic_inst.acc_wires\[15\]\[30\] net105 VGND VGND
+ VPWR VPWR _01008_ sky130_fd_sc_hd__a32o_1
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14666_ systolic_inst.acc_wires\[15\]\[16\] systolic_inst.acc_wires\[15\]\[17\] systolic_inst.acc_wires\[15\]\[18\]
+ systolic_inst.acc_wires\[15\]\[19\] systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _11824_ sky130_fd_sc_hd__o41a_1
X_17454_ systolic_inst.A_outs\[10\]\[6\] _04676_ _04677_ _04643_ VGND VGND VPWR VPWR
+ _04708_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13617_ deser_B.word_buffer\[53\] deser_B.serial_word\[53\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__mux2_1
X_16405_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[12\]\[6\]
+ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_215_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14597_ _11762_ _11764_ VGND VGND VPWR VPWR _11765_ sky130_fd_sc_hd__xor2_1
X_17385_ _04602_ _04639_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__and2_1
XFILLER_41_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19124_ _06188_ _06189_ _06159_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__a21o_1
XFILLER_119_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16336_ systolic_inst.A_outs\[12\]\[6\] _11260_ _03689_ _03692_ _03714_ VGND VGND
+ VPWR VPWR _03715_ sky130_fd_sc_hd__o311a_1
X_13548_ deser_A.shift_reg\[112\] deser_A.shift_reg\[113\] net129 VGND VGND VPWR VPWR
+ _00385_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19055_ net105 _06122_ _06123_ _06124_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__o31ai_1
X_16267_ _03646_ _03647_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__xnor2_1
X_13479_ deser_A.shift_reg\[43\] deser_A.shift_reg\[44\] net130 VGND VGND VPWR VPWR
+ _00316_ sky130_fd_sc_hd__mux2_1
XFILLER_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15218_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[14\]\[11\]
+ VGND VGND VPWR VPWR _12321_ sky130_fd_sc_hd__or2_1
X_18006_ systolic_inst.A_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[6\] _11263_ systolic_inst.A_outs\[9\]\[2\]
+ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_127_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16198_ _03542_ _03544_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15149_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[14\]\[1\]
+ VGND VGND VPWR VPWR _12262_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_166_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19957_ _06951_ _06952_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__and2_1
XFILLER_102_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18908_ _06001_ _06007_ _06008_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__o21ba_1
X_19888_ _06884_ _06885_ _06886_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__or3_1
XFILLER_132_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18839_ _05946_ _05950_ _05952_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__o211ai_2
XFILLER_132_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21850_ _08651_ _08652_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__nor2_1
XFILLER_110_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20801_ net106 systolic_inst.acc_wires\[5\]\[27\] net68 _07702_ VGND VGND VPWR VPWR
+ _01645_ sky130_fd_sc_hd__a22o_1
XFILLER_184_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21781_ _08585_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__inv_2
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23520_ net121 systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[9\] _10142_
+ _10143_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__o22a_1
XFILLER_211_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20732_ net60 _07644_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__nor2_1
XFILLER_223_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_186_Right_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23451_ _10074_ _10075_ VGND VGND VPWR VPWR _10076_ sky130_fd_sc_hd__nor2_1
X_20663_ net64 _07583_ _07585_ systolic_inst.acc_wires\[5\]\[6\] net109 VGND VGND
+ VPWR VPWR _01624_ sky130_fd_sc_hd__a32o_1
XFILLER_52_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_83_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22402_ _09140_ _09141_ VGND VGND VPWR VPWR _09143_ sky130_fd_sc_hd__and2b_1
XFILLER_195_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26170_ deser_B.serial_word\[125\] deser_B.shift_reg\[125\] net56 VGND VGND VPWR
+ VPWR _03472_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23382_ _09973_ _09977_ _09976_ VGND VGND VPWR VPWR _10009_ sky130_fd_sc_hd__o21bai_1
XFILLER_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20594_ _07435_ _07524_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__nor2_1
XFILLER_177_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25121_ C_out\[387\] net101 net73 ser_C.shift_reg\[387\] _11030_ VGND VGND VPWR VPWR
+ _02637_ sky130_fd_sc_hd__a221o_1
X_22333_ _09073_ _09074_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_115_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25052_ net112 ser_C.shift_reg\[354\] VGND VGND VPWR VPWR _10996_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22264_ _08954_ _08969_ _08968_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__o21a_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_225_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24003_ systolic_inst.B_shift\[9\]\[5\] B_in\[13\] _00008_ VGND VGND VPWR VPWR _10527_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_225_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21215_ _08049_ _08051_ _08082_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_225_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22195_ _08939_ _08940_ _08908_ _08910_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__o211a_1
XFILLER_191_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28811_ clknet_leaf_243_clk _02609_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[359\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_221_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21146_ _07959_ _07974_ _07973_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_221_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_221_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28742_ clknet_leaf_297_clk _02540_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[290\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_238_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25954_ systolic_inst.acc_wires\[13\]\[14\] C_out\[430\] net20 VGND VGND VPWR VPWR
+ _03256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21077_ _07946_ _07947_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20028_ _07018_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__inv_2
X_24905_ C_out\[279\] net103 net75 ser_C.shift_reg\[279\] _10922_ VGND VGND VPWR VPWR
+ _02529_ sky130_fd_sc_hd__a221o_1
XFILLER_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28673_ clknet_leaf_184_clk _02471_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[221\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25885_ systolic_inst.acc_wires\[11\]\[9\] C_out\[361\] net39 VGND VGND VPWR VPWR
+ _03187_ sky130_fd_sc_hd__mux2_1
XFILLER_73_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27624_ clknet_leaf_316_clk _01422_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24836_ net113 ser_C.shift_reg\[246\] VGND VGND VPWR VPWR _10888_ sky130_fd_sc_hd__and2_1
XFILLER_55_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_219_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24767_ C_out\[210\] net98 net78 ser_C.shift_reg\[210\] _10853_ VGND VGND VPWR VPWR
+ _02460_ sky130_fd_sc_hd__a221o_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27555_ clknet_leaf_304_clk _01353_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_21979_ _08759_ _08763_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__or2_1
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14520_ _11620_ _11689_ _11688_ VGND VGND VPWR VPWR _11699_ sky130_fd_sc_hd__a21o_1
XFILLER_215_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23718_ _10328_ _10329_ _10330_ VGND VGND VPWR VPWR _10331_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_29_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26506_ clknet_leaf_16_A_in_serial_clk _00309_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27486_ clknet_leaf_295_clk _01284_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24698_ net112 ser_C.shift_reg\[177\] VGND VGND VPWR VPWR _10819_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_29_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29225_ clknet_leaf_212_clk _03023_ net147 VGND VGND VPWR VPWR C_out\[197\] sky130_fd_sc_hd__dfrtp_1
X_14451_ _11600_ _11602_ _11631_ VGND VGND VPWR VPWR _11633_ sky130_fd_sc_hd__nand3_1
XFILLER_109_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23649_ _10222_ _10268_ VGND VGND VPWR VPWR _10269_ sky130_fd_sc_hd__nor2_1
X_26437_ clknet_leaf_8_clk _00244_ net134 VGND VGND VPWR VPWR A_in\[105\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13402_ A_in\[111\] deser_A.word_buffer\[111\] _00003_ VGND VGND VPWR VPWR _00250_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17170_ _04451_ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__nand2_1
XFILLER_122_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14382_ systolic_inst.A_outs\[15\]\[4\] systolic_inst.B_outs\[15\]\[5\] _11532_ _11531_
+ VGND VGND VPWR VPWR _11566_ sky130_fd_sc_hd__a31oi_2
XFILLER_70_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29156_ clknet_leaf_311_clk _02954_ net142 VGND VGND VPWR VPWR C_out\[128\] sky130_fd_sc_hd__dfrtp_1
X_26368_ clknet_leaf_26_clk _00175_ net137 VGND VGND VPWR VPWR A_in\[36\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16121_ _13085_ _03505_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__xnor2_1
X_28107_ clknet_leaf_155_clk _01905_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25319_ ser_C.parallel_data\[486\] net97 net77 ser_C.shift_reg\[486\] _11129_ VGND
+ VGND VPWR VPWR _02736_ sky130_fd_sc_hd__a221o_1
X_13333_ A_in\[42\] deser_A.word_buffer\[42\] net93 VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29087_ clknet_leaf_157_clk _02885_ net151 VGND VGND VPWR VPWR C_out\[59\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_210_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_130_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
X_26299_ clknet_leaf_22_A_in_serial_clk _00107_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_16052_ _13047_ _13048_ VGND VGND VPWR VPWR _13049_ sky130_fd_sc_hd__and2_1
X_28038_ clknet_leaf_163_clk _01836_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13264_ deser_A.word_buffer\[102\] deser_A.serial_word\[102\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__mux2_1
XFILLER_109_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15003_ _12079_ _12087_ _12086_ VGND VGND VPWR VPWR _12123_ sky130_fd_sc_hd__a21bo_1
X_13195_ deser_A.word_buffer\[33\] deser_A.serial_word\[33\] net127 VGND VGND VPWR
+ VPWR _00043_ sky130_fd_sc_hd__mux2_1
XFILLER_123_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19811_ _06770_ _06772_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__and2_1
XFILLER_123_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19742_ systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[6\] systolic_inst.A_outs\[6\]\[7\]
+ systolic_inst.B_outs\[6\]\[0\] VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__a22o_1
X_16954_ _04198_ _04245_ _04244_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__o21ba_1
XFILLER_238_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15905_ _12931_ VGND VGND VPWR VPWR _12932_ sky130_fd_sc_hd__inv_2
X_19673_ _06652_ _06658_ _06656_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_197_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_197_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16885_ systolic_inst.A_outs\[11\]\[5\] systolic_inst.B_outs\[11\]\[6\] systolic_inst.A_outs\[11\]\[6\]
+ systolic_inst.B_outs\[11\]\[7\] VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__and4b_1
XFILLER_65_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18624_ _05734_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__xor2_1
X_15836_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[13\]\[13\]
+ VGND VGND VPWR VPWR _12873_ sky130_fd_sc_hd__xor2_1
XFILLER_64_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18555_ _05656_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__nand2b_1
XFILLER_209_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15767_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[13\]\[3\]
+ VGND VGND VPWR VPWR _12814_ sky130_fd_sc_hd__nand2_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17506_ _04756_ _04757_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__xnor2_1
X_14718_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[28\]
+ VGND VGND VPWR VPWR _11868_ sky130_fd_sc_hd__nand2_1
X_18486_ _05594_ _05616_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__xor2_1
X_15698_ _12718_ _12721_ _12750_ VGND VGND VPWR VPWR _12751_ sky130_fd_sc_hd__o21ai_1
XFILLER_220_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17437_ _04689_ _04690_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_155_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14649_ net107 systolic_inst.acc_wires\[15\]\[17\] net69 _11809_ VGND VGND VPWR VPWR
+ _00995_ sky130_fd_sc_hd__a22o_1
XANTENNA_16 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_27 systolic_inst.A_outs\[1\]\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_38 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17368_ _04606_ _04623_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__xor2_1
XFILLER_140_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19107_ _06169_ _06172_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16319_ _03697_ _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_121_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_168_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17299_ _04556_ _04557_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_168_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19038_ _06101_ _06107_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_149_Left_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21000_ systolic_inst.B_outs\[4\]\[7\] _07839_ _07838_ VGND VGND VPWR VPWR _07873_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_173_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22951_ systolic_inst.A_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[5\] systolic_inst.B_outs\[1\]\[6\]
+ systolic_inst.B_outs\[1\]\[7\] VGND VGND VPWR VPWR _09629_ sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_188_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_188_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_96_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21902_ _08688_ _08692_ _08695_ _08696_ VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__o211a_1
X_25670_ systolic_inst.acc_wires\[4\]\[18\] C_out\[146\] net16 VGND VGND VPWR VPWR
+ _02972_ sky130_fd_sc_hd__mux2_1
Xmax_cap18 net21 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_6
XFILLER_56_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22882_ systolic_inst.A_outs\[1\]\[4\] systolic_inst.B_outs\[1\]\[5\] VGND VGND VPWR
+ VPWR _09562_ sky130_fd_sc_hd__nand2_1
XFILLER_44_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24621_ C_out\[137\] net103 net75 ser_C.shift_reg\[137\] _10780_ VGND VGND VPWR VPWR
+ _02387_ sky130_fd_sc_hd__a221o_1
XFILLER_71_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21833_ _08635_ _08636_ VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__nor2_1
XFILLER_83_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27340_ clknet_leaf_319_clk _01138_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_65_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24552_ net113 ser_C.shift_reg\[104\] VGND VGND VPWR VPWR _10746_ sky130_fd_sc_hd__and2_1
XFILLER_184_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21764_ _08553_ _08569_ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__xor2_1
XFILLER_180_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23503_ _10126_ VGND VGND VPWR VPWR _10127_ sky130_fd_sc_hd__inv_2
XFILLER_51_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20715_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[5\]\[13\]
+ _07625_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__a21oi_1
X_27271_ clknet_leaf_266_clk _01069_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24483_ C_out\[68\] _11302_ net81 ser_C.shift_reg\[68\] _10711_ VGND VGND VPWR VPWR
+ _02318_ sky130_fd_sc_hd__a221o_1
X_21695_ _08462_ _08463_ _08465_ VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__o21a_1
X_29010_ clknet_leaf_103_clk _02808_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_221_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26222_ clknet_leaf_8_A_in_serial_clk _00030_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23434_ _10056_ _10057_ _10015_ _10017_ VGND VGND VPWR VPWR _10060_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_78_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20646_ _07568_ _07569_ _07570_ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_24_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26153_ deser_B.serial_word\[108\] deser_B.shift_reg\[108\] _00001_ VGND VGND VPWR
+ VPWR _03455_ sky130_fd_sc_hd__mux2_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_227_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23365_ _09990_ _09991_ VGND VGND VPWR VPWR _09992_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_112_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20577_ _07464_ _07478_ _07476_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__o21a_1
XFILLER_221_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25104_ net113 ser_C.shift_reg\[380\] VGND VGND VPWR VPWR _11022_ sky130_fd_sc_hd__and2_1
X_22316_ systolic_inst.B_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[6\] systolic_inst.A_outs\[2\]\[7\]
+ systolic_inst.B_outs\[2\]\[3\] VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__a22o_1
XFILLER_180_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26084_ deser_B.serial_word\[39\] deser_B.shift_reg\[39\] net55 VGND VGND VPWR VPWR
+ _03386_ sky130_fd_sc_hd__mux2_1
X_23296_ _09924_ _09926_ VGND VGND VPWR VPWR _09927_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_223_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25035_ C_out\[344\] net97 net77 ser_C.shift_reg\[344\] _10987_ VGND VGND VPWR VPWR
+ _02594_ sky130_fd_sc_hd__a221o_1
X_22247_ _08990_ _08991_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__nor2_1
XFILLER_191_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22178_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[4\] _08923_ _08924_
+ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__nand4_2
XFILLER_152_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21129_ systolic_inst.A_outs\[4\]\[6\] _07884_ _07998_ VGND VGND VPWR VPWR _07999_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26986_ clknet_leaf_0_A_in_serial_clk _00784_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28725_ clknet_leaf_312_clk _02523_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[273\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_179_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_179_clk
+ sky130_fd_sc_hd__clkbuf_8
X_25937_ systolic_inst.acc_wires\[12\]\[29\] C_out\[413\] net21 VGND VGND VPWR VPWR
+ _03239_ sky130_fd_sc_hd__mux2_1
X_13951_ deser_A.serial_word\[112\] deser_A.shift_reg\[112\] net57 VGND VGND VPWR
+ VPWR _00777_ sky130_fd_sc_hd__mux2_1
XFILLER_232_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_222_Right_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28656_ clknet_leaf_204_clk _02454_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[204\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16670_ _03988_ _03991_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__xnor2_1
X_13882_ deser_A.serial_word\[43\] deser_A.shift_reg\[43\] net58 VGND VGND VPWR VPWR
+ _00708_ sky130_fd_sc_hd__mux2_1
X_25868_ systolic_inst.acc_wires\[10\]\[24\] C_out\[344\] net11 VGND VGND VPWR VPWR
+ _03170_ sky130_fd_sc_hd__mux2_1
XFILLER_100_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27607_ clknet_leaf_204_clk _01405_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_15621_ _12674_ _12676_ VGND VGND VPWR VPWR _12677_ sky130_fd_sc_hd__or2_1
X_24819_ C_out\[236\] net99 net79 ser_C.shift_reg\[236\] _10879_ VGND VGND VPWR VPWR
+ _02486_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28587_ clknet_leaf_308_clk _02385_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[135\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25799_ systolic_inst.acc_wires\[8\]\[19\] C_out\[275\] net22 VGND VGND VPWR VPWR
+ _03101_ sky130_fd_sc_hd__mux2_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18340_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[22\]
+ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__nand2_1
X_15552_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[8\] _12609_ net115
+ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__mux2_1
X_27538_ clknet_leaf_311_clk _01336_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_187_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_191_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_191_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14503_ _11657_ _11659_ _11682_ VGND VGND VPWR VPWR _11683_ sky130_fd_sc_hd__a21oi_1
X_15483_ _12540_ _12541_ VGND VGND VPWR VPWR _12542_ sky130_fd_sc_hd__nand2_1
X_18271_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[9\]\[11\]
+ _05439_ _05442_ _05443_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_212_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27469_ clknet_leaf_298_clk _01267_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_212_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29208_ clknet_leaf_205_clk _03006_ net146 VGND VGND VPWR VPWR C_out\[180\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _04481_ _04482_ _04468_ _04471_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__o211a_1
XFILLER_202_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14434_ _11586_ _11616_ VGND VGND VPWR VPWR _11617_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29139_ clknet_leaf_167_clk _02937_ net152 VGND VGND VPWR VPWR C_out\[111\] sky130_fd_sc_hd__dfrtp_1
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17153_ _04431_ _04435_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__nor2_1
XFILLER_122_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14365_ _11508_ _11510_ VGND VGND VPWR VPWR _11550_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_103_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_200_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13316_ A_in\[25\] deser_A.word_buffer\[25\] net91 VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__mux2_1
X_16104_ _13095_ _13098_ VGND VGND VPWR VPWR _13099_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17084_ net105 systolic_inst.acc_wires\[11\]\[16\] _04378_ _04380_ VGND VGND VPWR
+ VPWR _01250_ sky130_fd_sc_hd__a22o_1
XFILLER_171_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14296_ _11475_ _11481_ VGND VGND VPWR VPWR _11482_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16035_ _13027_ _13030_ VGND VGND VPWR VPWR _13032_ sky130_fd_sc_hd__xnor2_1
X_13247_ deser_A.word_buffer\[85\] deser_A.serial_word\[85\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13178_ deser_A.word_buffer\[16\] deser_A.serial_word\[16\] net128 VGND VGND VPWR
+ VPWR _00026_ sky130_fd_sc_hd__mux2_1
XFILLER_123_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17986_ _05137_ _05139_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__and2_1
XFILLER_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19725_ _06725_ _06727_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__nor2_1
XFILLER_81_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16937_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[13\] _04252_ net119
+ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__mux2_1
XFILLER_226_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19656_ _06659_ _06660_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16868_ _04183_ _04184_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_0_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18607_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[7\] VGND VGND VPWR
+ VPWR _05735_ sky130_fd_sc_hd__nand2_4
XFILLER_93_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15819_ net108 systolic_inst.acc_wires\[13\]\[10\] net67 _12858_ VGND VGND VPWR VPWR
+ _01116_ sky130_fd_sc_hd__a22o_1
XFILLER_20_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19587_ _06609_ _06613_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_157_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16799_ _04116_ _04117_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_103_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18538_ _05666_ _05667_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__or2_1
XFILLER_181_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18469_ _05581_ _05583_ _05582_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__a21bo_1
XFILLER_61_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_342_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_342_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_60_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20500_ _07398_ _07433_ systolic_inst.A_outs\[5\]\[7\] VGND VGND VPWR VPWR _07434_
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_60_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21480_ net122 systolic_inst.B_outs\[3\]\[0\] systolic_inst.A_outs\[3\]\[0\] VGND
+ VGND VPWR VPWR _08297_ sky130_fd_sc_hd__and3_1
XFILLER_14_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20431_ _07365_ _07366_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__nor2_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_157_Left_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23150_ _09808_ _09809_ _09810_ VGND VGND VPWR VPWR _09811_ sky130_fd_sc_hd__and3_1
XFILLER_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload230 clknet_leaf_77_clk VGND VGND VPWR VPWR clkload230/Y sky130_fd_sc_hd__clkinvlp_4
X_20362_ _07295_ _07299_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__xnor2_1
Xclkload241 clknet_leaf_51_clk VGND VGND VPWR VPWR clkload241/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload252 clknet_leaf_131_clk VGND VGND VPWR VPWR clkload252/Y sky130_fd_sc_hd__inv_6
XFILLER_162_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload263 clknet_leaf_106_clk VGND VGND VPWR VPWR clkload263/X sky130_fd_sc_hd__clkbuf_8
XFILLER_228_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22101_ systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[2\]
+ systolic_inst.B_outs\[2\]\[0\] VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__a22oi_1
XFILLER_179_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload274 clknet_leaf_132_clk VGND VGND VPWR VPWR clkload274/Y sky130_fd_sc_hd__clkinv_2
XFILLER_162_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23081_ _09749_ _09750_ _09751_ VGND VGND VPWR VPWR _09752_ sky130_fd_sc_hd__a21o_1
Xclkload285 clknet_leaf_189_clk VGND VGND VPWR VPWR clkload285/Y sky130_fd_sc_hd__inv_6
X_20293_ _07216_ _07232_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__xor2_1
Xclkload296 clknet_leaf_176_clk VGND VGND VPWR VPWR clkload296/Y sky130_fd_sc_hd__inv_6
XFILLER_216_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22032_ _08805_ _08808_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26840_ clknet_leaf_83_clk _00642_ net144 VGND VGND VPWR VPWR B_in\[112\] sky130_fd_sc_hd__dfrtp_1
XFILLER_88_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26771_ clknet_leaf_94_clk _00573_ net152 VGND VGND VPWR VPWR B_in\[43\] sky130_fd_sc_hd__dfrtp_1
X_23983_ systolic_inst.B_shift\[12\]\[3\] B_in\[67\] _00008_ VGND VGND VPWR VPWR _10517_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28510_ clknet_leaf_157_clk _02308_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22934_ _09552_ _09578_ _09577_ VGND VGND VPWR VPWR _09613_ sky130_fd_sc_hd__a21boi_1
X_25722_ systolic_inst.acc_wires\[6\]\[6\] C_out\[198\] net47 VGND VGND VPWR VPWR
+ _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_5_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29490_ clknet_leaf_284_clk _03288_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_228_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28441_ clknet_leaf_34_clk _02239_ VGND VGND VPWR VPWR systolic_inst.A_shift\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_216_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22865_ _09545_ _09544_ VGND VGND VPWR VPWR _09546_ sky130_fd_sc_hd__nand2b_1
XFILLER_186_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25653_ systolic_inst.acc_wires\[4\]\[1\] C_out\[129\] net29 VGND VGND VPWR VPWR
+ _02955_ sky130_fd_sc_hd__mux2_1
XFILLER_231_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21816_ _08588_ _08591_ _08619_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__o21ai_1
X_24604_ net110 ser_C.shift_reg\[130\] VGND VGND VPWR VPWR _10772_ sky130_fd_sc_hd__and2_1
X_25584_ systolic_inst.acc_wires\[1\]\[28\] C_out\[60\] net52 VGND VGND VPWR VPWR
+ _02886_ sky130_fd_sc_hd__mux2_1
Xwire71 _11332_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_16
X_28372_ clknet_leaf_30_clk _02170_ VGND VGND VPWR VPWR systolic_inst.A_shift\[19\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22796_ _09457_ _09459_ VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__nand2_1
XFILLER_197_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24535_ C_out\[94\] net100 net82 ser_C.shift_reg\[94\] _10737_ VGND VGND VPWR VPWR
+ _02344_ sky130_fd_sc_hd__a221o_1
XFILLER_184_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27323_ clknet_leaf_329_clk _01121_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_240_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21747_ _08551_ _08552_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__nand2_1
XFILLER_196_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_333_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_333_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24466_ net114 ser_C.shift_reg\[61\] VGND VGND VPWR VPWR _10703_ sky130_fd_sc_hd__and2_1
XFILLER_200_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27254_ clknet_leaf_281_clk _01052_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_21678_ systolic_inst.B_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[5\] systolic_inst.A_outs\[3\]\[6\]
+ systolic_inst.B_outs\[3\]\[3\] VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__a22oi_1
XFILLER_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23417_ _10039_ _10042_ VGND VGND VPWR VPWR _10043_ sky130_fd_sc_hd__xor2_1
X_26205_ clknet_leaf_15_A_in_serial_clk _00013_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20629_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[5\]\[2\]
+ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__nand2_1
XFILLER_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27185_ clknet_leaf_253_clk _00983_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24397_ C_out\[25\] _11302_ net82 ser_C.shift_reg\[25\] _10668_ VGND VGND VPWR VPWR
+ _02275_ sky130_fd_sc_hd__a221o_1
XFILLER_123_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26136_ deser_B.serial_word\[91\] deser_B.shift_reg\[91\] net56 VGND VGND VPWR VPWR
+ _03438_ sky130_fd_sc_hd__mux2_1
X_14150_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[2\] _11339_ _11340_
+ VGND VGND VPWR VPWR _11342_ sky130_fd_sc_hd__a22oi_1
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23348_ _09949_ _09974_ _09975_ VGND VGND VPWR VPWR _09976_ sky130_fd_sc_hd__nor3_1
XFILLER_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13101_ systolic_inst.cycle_cnt\[2\] VGND VGND VPWR VPWR _11257_ sky130_fd_sc_hd__inv_2
XFILLER_98_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14081_ deser_B.shift_reg\[115\] deser_B.shift_reg\[116\] deser_B.receiving VGND
+ VGND VPWR VPWR _00907_ sky130_fd_sc_hd__mux2_1
X_26067_ deser_B.serial_word\[22\] deser_B.shift_reg\[22\] net55 VGND VGND VPWR VPWR
+ _03369_ sky130_fd_sc_hd__mux2_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23279_ systolic_inst.A_outs\[0\]\[2\] systolic_inst.A_shift\[0\]\[2\] net121 VGND
+ VGND VPWR VPWR _01908_ sky130_fd_sc_hd__mux2_1
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25018_ net111 ser_C.shift_reg\[337\] VGND VGND VPWR VPWR _10979_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_56_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17840_ _05018_ _05035_ _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_205_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17771_ _04988_ _04990_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_197_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14983_ _12103_ _12102_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[9\]
+ net107 VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__a2bb2o_1
X_26969_ clknet_leaf_23_A_in_serial_clk _00767_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_201_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19510_ _06542_ _06550_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__or2_1
XFILLER_120_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28708_ clknet_leaf_325_clk _02506_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[256\]
+ sky130_fd_sc_hd__dfrtp_1
X_16722_ _04005_ _04007_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_1_A_in_serial_clk clknet_2_0__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_1_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_207_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13934_ deser_A.serial_word\[95\] deser_A.shift_reg\[95\] net57 VGND VGND VPWR VPWR
+ _00760_ sky130_fd_sc_hd__mux2_1
X_29688_ clknet_leaf_106_clk _03483_ net151 VGND VGND VPWR VPWR ser_C.bit_idx\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_193_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19441_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[7\]\[6\]
+ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_193_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28639_ clknet_leaf_179_clk _02437_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[187\]
+ sky130_fd_sc_hd__dfrtp_1
X_16653_ _03975_ _03976_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__or2_1
X_13865_ deser_A.serial_word\[26\] deser_A.shift_reg\[26\] net58 VGND VGND VPWR VPWR
+ _00691_ sky130_fd_sc_hd__mux2_1
XFILLER_235_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15604_ _12650_ _12658_ VGND VGND VPWR VPWR _12660_ sky130_fd_sc_hd__or2_1
X_19372_ systolic_inst.B_outs\[7\]\[5\] systolic_inst.B_outs\[7\]\[6\] systolic_inst.A_outs\[7\]\[7\]
+ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__nand3_1
X_16584_ systolic_inst.B_outs\[10\]\[1\] systolic_inst.B_outs\[6\]\[1\] net120 VGND
+ VGND VPWR VPWR _01211_ sky130_fd_sc_hd__mux2_1
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13796_ B_in\[103\] deser_B.word_buffer\[103\] _00005_ VGND VGND VPWR VPWR _00633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_215_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18323_ _05488_ _05487_ systolic_inst.acc_wires\[9\]\[19\] net106 VGND VGND VPWR
+ VPWR _01381_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_152_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _12591_ _12592_ VGND VGND VPWR VPWR _12593_ sky130_fd_sc_hd__and2_1
XFILLER_206_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_324_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_324_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18254_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[9\]\[10\]
+ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__or2_1
X_15466_ _12523_ _12524_ _12494_ VGND VGND VPWR VPWR _12526_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17205_ _04461_ _04467_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__or2_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14417_ _11599_ _11598_ VGND VGND VPWR VPWR _11600_ sky130_fd_sc_hd__nand2b_1
XFILLER_30_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18185_ _05292_ _05356_ _05354_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__a21oi_1
X_15397_ _12446_ _12448_ _12459_ VGND VGND VPWR VPWR _12460_ sky130_fd_sc_hd__and3_1
XFILLER_200_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17136_ _04418_ _04420_ _04423_ net60 VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__a31o_1
XFILLER_239_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14348_ _11528_ _11532_ VGND VGND VPWR VPWR _11533_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14279_ _11465_ _11464_ VGND VGND VPWR VPWR _11466_ sky130_fd_sc_hd__and2b_1
X_17067_ _04358_ _04365_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__nand2_1
X_16018_ _13009_ _13015_ VGND VGND VPWR VPWR _13016_ sky130_fd_sc_hd__nor2_1
XFILLER_98_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_999 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17969_ systolic_inst.A_outs\[9\]\[2\] systolic_inst.B_outs\[9\]\[6\] _11263_ systolic_inst.A_outs\[9\]\[1\]
+ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19708_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[5\] _06710_
+ _06711_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__a22o_1
X_20980_ _07850_ _07851_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19639_ _06638_ _06644_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_101_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22650_ _09343_ _09345_ _09357_ _09358_ _09351_ VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__a311oi_4
XTAP_TAPCELL_ROW_62_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21601_ _08409_ _08410_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__nor2_1
XFILLER_179_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22581_ net60 _09301_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__nor2_1
XFILLER_55_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_315_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_315_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_142_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24320_ _10633_ systolic_inst.A_shift\[10\]\[7\] net71 VGND VGND VPWR VPWR _02233_
+ sky130_fd_sc_hd__mux2_1
X_21532_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[5\] VGND
+ VGND VPWR VPWR _08344_ sky130_fd_sc_hd__and2_1
XFILLER_181_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24251_ systolic_inst.A_shift\[17\]\[2\] net70 net83 systolic_inst.A_shift\[18\]\[2\]
+ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__a22o_1
X_21463_ _08296_ _08295_ systolic_inst.acc_wires\[4\]\[31\] _11258_ VGND VGND VPWR
+ VPWR _01713_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_135_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23202_ _09853_ _09854_ VGND VGND VPWR VPWR _09855_ sky130_fd_sc_hd__and2_1
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20414_ _07319_ _07349_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24182_ systolic_inst.A_shift\[25\]\[5\] net70 _10505_ systolic_inst.A_shift\[26\]\[5\]
+ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21394_ _08236_ _08237_ _08233_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_96_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23133_ _09794_ _09795_ VGND VGND VPWR VPWR _09796_ sky130_fd_sc_hd__and2_1
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20345_ _07252_ _07283_ VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28990_ clknet_leaf_57_clk _02788_ VGND VGND VPWR VPWR systolic_inst.A_shift\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_92_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27941_ clknet_leaf_170_clk _01739_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_23064_ _09736_ _09737_ VGND VGND VPWR VPWR _09738_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20276_ _07197_ _07214_ _07216_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__and3_1
XFILLER_118_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_241_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_241_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22015_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[22\]
+ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__nor2_1
X_27872_ clknet_leaf_38_clk _01670_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29611_ clknet_leaf_24_B_in_serial_clk _03406_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26823_ clknet_leaf_71_clk _00625_ net135 VGND VGND VPWR VPWR B_in\[95\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29542_ clknet_leaf_105_clk _00000_ net152 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_4
XFILLER_124_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26754_ clknet_leaf_61_clk _00556_ net143 VGND VGND VPWR VPWR B_in\[26\] sky130_fd_sc_hd__dfrtp_1
X_23966_ _10508_ systolic_inst.B_shift\[9\]\[2\] net72 VGND VGND VPWR VPWR _02004_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25705_ systolic_inst.acc_wires\[5\]\[21\] C_out\[181\] net45 VGND VGND VPWR VPWR
+ _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_72_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22917_ _09594_ _09595_ VGND VGND VPWR VPWR _09596_ sky130_fd_sc_hd__nor2_1
X_29473_ clknet_leaf_284_clk _03271_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[445\]
+ sky130_fd_sc_hd__dfrtp_1
X_23897_ _10481_ systolic_inst.B_shift\[13\]\[0\] net72 VGND VGND VPWR VPWR _01962_
+ sky130_fd_sc_hd__mux2_1
X_26685_ clknet_leaf_28_B_in_serial_clk _00488_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_205_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28424_ clknet_leaf_14_clk _02222_ VGND VGND VPWR VPWR systolic_inst.A_shift\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_231_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25636_ systolic_inst.acc_wires\[3\]\[16\] C_out\[112\] net49 VGND VGND VPWR VPWR
+ _02938_ sky130_fd_sc_hd__mux2_1
X_22848_ _09526_ _09527_ VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__xnor2_1
X_13650_ deser_B.word_buffer\[86\] deser_B.serial_word\[86\] net124 VGND VGND VPWR
+ VPWR _00487_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13581_ deser_B.word_buffer\[17\] deser_B.serial_word\[17\] net124 VGND VGND VPWR
+ VPWR _00418_ sky130_fd_sc_hd__mux2_1
XFILLER_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28355_ clknet_leaf_342_clk _02153_ VGND VGND VPWR VPWR systolic_inst.A_shift\[24\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25567_ systolic_inst.acc_wires\[1\]\[11\] C_out\[43\] net36 VGND VGND VPWR VPWR
+ _02869_ sky130_fd_sc_hd__mux2_1
X_22779_ systolic_inst.A_outs\[1\]\[1\] systolic_inst.B_outs\[1\]\[5\] systolic_inst.B_outs\[1\]\[6\]
+ systolic_inst.A_outs\[1\]\[0\] VGND VGND VPWR VPWR _09462_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_306_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_306_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27306_ clknet_leaf_329_clk _01104_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_15320_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[26\]
+ VGND VGND VPWR VPWR _12408_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24518_ net114 ser_C.shift_reg\[87\] VGND VGND VPWR VPWR _10729_ sky130_fd_sc_hd__and2_1
XFILLER_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25498_ systolic_inst.cycle_cnt\[22\] _11279_ _11225_ systolic_inst.cycle_cnt\[21\]
+ VGND VGND VPWR VPWR _11229_ sky130_fd_sc_hd__a22oi_1
XFILLER_169_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28286_ clknet_leaf_61_clk _02084_ VGND VGND VPWR VPWR systolic_inst.B_shift\[19\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15251_ _12341_ _12345_ _12347_ _12348_ VGND VGND VPWR VPWR _12350_ sky130_fd_sc_hd__a211o_1
XFILLER_8_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27237_ clknet_leaf_278_clk _01035_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24449_ C_out\[51\] _11302_ net81 ser_C.shift_reg\[51\] _10694_ VGND VGND VPWR VPWR
+ _02301_ sky130_fd_sc_hd__a221o_1
XFILLER_201_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14202_ _11388_ _11389_ _11387_ VGND VGND VPWR VPWR _11391_ sky130_fd_sc_hd__o21ai_1
X_15182_ _12290_ VGND VGND VPWR VPWR _12291_ sky130_fd_sc_hd__inv_2
XFILLER_201_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27168_ clknet_leaf_253_clk _00966_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_186_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14133_ systolic_inst.B_outs\[14\]\[1\] systolic_inst.B_outs\[10\]\[1\] net120 VGND
+ VGND VPWR VPWR _00955_ sky130_fd_sc_hd__mux2_1
X_26119_ deser_B.serial_word\[74\] deser_B.shift_reg\[74\] _00001_ VGND VGND VPWR
+ VPWR _03421_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_207_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19990_ _06958_ _06960_ _06983_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__and3_1
X_27099_ clknet_leaf_7_B_in_serial_clk _00897_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14064_ deser_B.shift_reg\[98\] deser_B.shift_reg\[99\] net126 VGND VGND VPWR VPWR
+ _00890_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18941_ _06039_ _06040_ _06037_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_203_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18872_ _05981_ _05980_ systolic_inst.acc_wires\[8\]\[11\] net108 VGND VGND VPWR
+ VPWR _01437_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_141_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17823_ _05009_ _05019_ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_141_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17754_ _04974_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14966_ _12084_ _12085_ VGND VGND VPWR VPWR _12087_ sky130_fd_sc_hd__xnor2_1
X_16705_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[5\] VGND VGND
+ VPWR VPWR _04027_ sky130_fd_sc_hd__nand2_1
X_13917_ deser_A.serial_word\[78\] deser_A.shift_reg\[78\] net57 VGND VGND VPWR VPWR
+ _00743_ sky130_fd_sc_hd__mux2_1
XFILLER_169_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17685_ _04905_ _04912_ _04913_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__o21ba_1
XFILLER_74_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14897_ _12017_ _12018_ VGND VGND VPWR VPWR _12020_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19424_ _06477_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__inv_2
XFILLER_39_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16636_ _03942_ _03958_ _03959_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__and3_1
XFILLER_78_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13848_ deser_A.serial_word\[9\] deser_A.shift_reg\[9\] net58 VGND VGND VPWR VPWR
+ _00674_ sky130_fd_sc_hd__mux2_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19355_ _06413_ _06414_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__nand2_1
XFILLER_62_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16567_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[30\]
+ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__or2_1
X_13779_ B_in\[86\] deser_B.word_buffer\[86\] net85 VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__mux2_1
XFILLER_95_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18306_ net60 _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__nor2_1
X_15518_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[7\]
+ VGND VGND VPWR VPWR _12576_ sky130_fd_sc_hd__o21a_1
X_19286_ _06277_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__xnor2_4
XFILLER_128_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16498_ net67 _03855_ _03856_ systolic_inst.acc_wires\[12\]\[18\] net108 VGND VGND
+ VPWR VPWR _01188_ sky130_fd_sc_hd__a32o_1
XFILLER_200_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18237_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[9\]\[7\]
+ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__or2_1
X_15449_ systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[5\] systolic_inst.A_outs\[13\]\[6\]
+ systolic_inst.B_outs\[13\]\[0\] VGND VGND VPWR VPWR _12509_ sky130_fd_sc_hd__a22oi_1
XFILLER_164_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18168_ _05327_ _05329_ _05353_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__and3_1
Xmax_cap100 _11302_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_12
XFILLER_11_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap122 systolic_inst.ce_local VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_12
X_17119_ _04401_ _04402_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__nor2_1
Xmax_cap133 net134 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_16
Xmax_cap144 net153 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_16
XFILLER_171_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18099_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[7\] _05260_ _05224_
+ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__a31o_1
XFILLER_176_1356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20130_ _07105_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__inv_2
XFILLER_116_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20061_ _07044_ _07045_ _07046_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__a21o_1
XFILLER_219_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23820_ _10416_ _10417_ VGND VGND VPWR VPWR _10418_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23751_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[0\]\[8\]
+ _10355_ VGND VGND VPWR VPWR _10359_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_124_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20963_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.A_outs\[4\]\[4\] VGND VGND VPWR
+ VPWR _07837_ sky130_fd_sc_hd__nand2_1
XFILLER_199_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_92_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_93_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22702_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[2\] _09387_ VGND
+ VGND VPWR VPWR _09389_ sky130_fd_sc_hd__a21o_1
XFILLER_183_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23682_ _10253_ _10280_ _10300_ VGND VGND VPWR VPWR _10301_ sky130_fd_sc_hd__a21oi_2
X_26470_ clknet_leaf_57_clk net94 net137 VGND VGND VPWR VPWR A_in_valid sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_85_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20894_ _07748_ _07770_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__or2_1
X_22633_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[25\]
+ VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__xor2_2
X_25421_ systolic_inst.A_shift\[1\]\[2\] A_in\[2\] net59 VGND VGND VPWR VPWR _11180_
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28140_ clknet_leaf_124_clk _01938_ net153 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_25352_ net112 ser_C.shift_reg\[504\] VGND VGND VPWR VPWR _11146_ sky130_fd_sc_hd__and2_1
X_22564_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[2\]\[13\]
+ _09282_ VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_230_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_230_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21515_ _08324_ _08327_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24303_ systolic_inst.A_shift\[12\]\[7\] A_in\[55\] net59 VGND VGND VPWR VPWR _10625_
+ sky130_fd_sc_hd__mux2_1
X_28071_ clknet_leaf_119_clk _01869_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_25283_ ser_C.parallel_data\[468\] net102 net74 ser_C.shift_reg\[468\] _11111_ VGND
+ VGND VPWR VPWR _02718_ sky130_fd_sc_hd__a221o_1
X_22495_ _09225_ _09226_ _09227_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__a21o_1
XFILLER_186_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27022_ clknet_leaf_25_B_in_serial_clk _00820_ net143 VGND VGND VPWR VPWR deser_B.shift_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_24234_ _10602_ systolic_inst.A_shift\[18\]\[0\] net70 VGND VGND VPWR VPWR _02178_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21446_ _11258_ systolic_inst.acc_wires\[4\]\[28\] net63 _08282_ VGND VGND VPWR VPWR
+ _01710_ sky130_fd_sc_hd__a22o_1
XFILLER_148_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24165_ systolic_inst.A_shift\[28\]\[6\] A_in\[102\] net59 VGND VGND VPWR VPWR _10584_
+ sky130_fd_sc_hd__mux2_1
X_21377_ systolic_inst.acc_wires\[4\]\[16\] systolic_inst.acc_wires\[4\]\[17\] systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__o21ai_1
X_23116_ _09779_ _09780_ _09781_ VGND VGND VPWR VPWR _09782_ sky130_fd_sc_hd__a21o_1
X_20328_ systolic_inst.A_outs\[5\]\[1\] systolic_inst.B_outs\[5\]\[6\] VGND VGND VPWR
+ VPWR _07267_ sky130_fd_sc_hd__nand2_1
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24096_ _10557_ systolic_inst.B_shift\[19\]\[3\] net71 VGND VGND VPWR VPWR _02085_
+ sky130_fd_sc_hd__mux2_1
X_28973_ clknet_leaf_63_clk _02771_ VGND VGND VPWR VPWR systolic_inst.A_shift\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27924_ clknet_leaf_123_clk _01722_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_23047_ _09720_ _09721_ VGND VGND VPWR VPWR _09722_ sky130_fd_sc_hd__nor2_1
XFILLER_66_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20259_ _07190_ _07199_ _07200_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_38_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27855_ clknet_leaf_35_clk _01653_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_27_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26806_ clknet_leaf_82_clk _00608_ net153 VGND VGND VPWR VPWR B_in\[78\] sky130_fd_sc_hd__dfrtp_1
X_14820_ systolic_inst.A_outs\[14\]\[2\] systolic_inst.B_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\]
+ systolic_inst.A_outs\[14\]\[1\] VGND VGND VPWR VPWR _11945_ sky130_fd_sc_hd__a22o_1
X_27786_ clknet_leaf_183_clk _01584_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_24998_ net111 ser_C.shift_reg\[327\] VGND VGND VPWR VPWR _10969_ sky130_fd_sc_hd__and2_1
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29525_ clknet_leaf_261_clk _03323_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26737_ clknet_leaf_103_clk _00539_ net151 VGND VGND VPWR VPWR B_in\[9\] sky130_fd_sc_hd__dfrtp_1
X_14751_ systolic_inst.B_outs\[13\]\[3\] systolic_inst.B_outs\[9\]\[3\] net115 VGND
+ VGND VPWR VPWR _01021_ sky130_fd_sc_hd__mux2_1
XFILLER_229_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23949_ _10503_ systolic_inst.B_shift\[10\]\[6\] net70 VGND VGND VPWR VPWR _01992_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_83_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
X_13702_ B_in\[9\] deser_B.word_buffer\[9\] net84 VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29456_ clknet_leaf_288_clk _03254_ net136 VGND VGND VPWR VPWR C_out\[428\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17470_ _04714_ _04722_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__xnor2_1
XFILLER_229_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26668_ clknet_leaf_8_B_in_serial_clk _00471_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_14682_ net69 _11836_ _11837_ systolic_inst.acc_wires\[15\]\[22\] net107 VGND VGND
+ VPWR VPWR _01000_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_103_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28407_ clknet_leaf_88_clk _02205_ VGND VGND VPWR VPWR systolic_inst.B_shift\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16421_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[12\]\[9\]
+ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__and2_1
XFILLER_38_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25619_ systolic_inst.acc_wires\[2\]\[31\] C_out\[95\] net50 VGND VGND VPWR VPWR
+ _02921_ sky130_fd_sc_hd__mux2_1
X_13633_ deser_B.word_buffer\[69\] deser_B.serial_word\[69\] net123 VGND VGND VPWR
+ VPWR _00470_ sky130_fd_sc_hd__mux2_1
XFILLER_60_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29387_ clknet_leaf_243_clk _03185_ net145 VGND VGND VPWR VPWR C_out\[359\] sky130_fd_sc_hd__dfrtp_1
XFILLER_242_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26599_ clknet_leaf_3_B_in_serial_clk _00402_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_125_1200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19140_ _06200_ _06204_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16352_ _03728_ _03729_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__xnor2_1
X_28338_ clknet_leaf_2_clk _02136_ VGND VGND VPWR VPWR systolic_inst.A_shift\[26\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13564_ deser_B.word_buffer\[0\] deser_B.serial_word\[0\] net124 VGND VGND VPWR VPWR
+ _00401_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15303_ _12386_ _12390_ _12393_ VGND VGND VPWR VPWR _12394_ sky130_fd_sc_hd__nand3_1
X_19071_ _06137_ _06138_ _06117_ _06120_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__o211ai_2
XFILLER_201_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28269_ clknet_leaf_48_clk _02067_ VGND VGND VPWR VPWR systolic_inst.B_shift\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16283_ systolic_inst.B_outs\[12\]\[5\] systolic_inst.A_outs\[12\]\[7\] VGND VGND
+ VPWR VPWR _03664_ sky130_fd_sc_hd__nand2_1
X_13495_ deser_A.shift_reg\[59\] deser_A.shift_reg\[60\] net130 VGND VGND VPWR VPWR
+ _00332_ sky130_fd_sc_hd__mux2_1
XFILLER_200_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18022_ _05175_ _05177_ _05212_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__and3_1
X_15234_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[14\]\[13\]
+ VGND VGND VPWR VPWR _12335_ sky130_fd_sc_hd__xor2_1
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15165_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[14\]\[3\]
+ VGND VGND VPWR VPWR _12276_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_112_Left_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14116_ systolic_inst.A_shift\[21\]\[0\] net71 _11333_ A_in\[88\] VGND VGND VPWR
+ VPWR _00938_ sky130_fd_sc_hd__a22o_1
X_19973_ _06966_ _06967_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__and2b_1
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15096_ _12211_ _12212_ VGND VGND VPWR VPWR _12213_ sky130_fd_sc_hd__and2_1
XFILLER_119_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18924_ _06025_ _06026_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nand2_1
X_14047_ deser_B.shift_reg\[81\] deser_B.shift_reg\[82\] deser_B.receiving VGND VGND
+ VPWR VPWR _00873_ sky130_fd_sc_hd__mux2_1
XFILLER_136_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18855_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[8\]\[9\]
+ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__nand2_1
XFILLER_227_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17806_ net116 _05005_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__and2_1
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18786_ _05908_ _05907_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__nand2b_1
XFILLER_227_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ _12994_ _12995_ _12983_ VGND VGND VPWR VPWR _12997_ sky130_fd_sc_hd__a21o_1
XFILLER_67_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17737_ systolic_inst.acc_wires\[10\]\[20\] systolic_inst.acc_wires\[10\]\[21\] systolic_inst.acc_wires\[10\]\[22\]
+ systolic_inst.acc_wires\[10\]\[23\] systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__o41a_1
XPHY_EDGE_ROW_121_Left_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14949_ _12028_ _12034_ _12033_ VGND VGND VPWR VPWR _12070_ sky130_fd_sc_hd__a21o_1
XFILLER_224_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_36_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17668_ _04899_ _04901_ _04903_ systolic_inst.acc_wires\[10\]\[13\] net105 VGND VGND
+ VPWR VPWR _01311_ sky130_fd_sc_hd__a32o_1
XFILLER_235_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_888 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19407_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[7\]\[1\]
+ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_173_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16619_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[2\] VGND VGND
+ VPWR VPWR _03944_ sky130_fd_sc_hd__and2_1
XFILLER_223_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17599_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[10\]\[4\]
+ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_98_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19338_ _06398_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__inv_2
XFILLER_17_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_3_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_17_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19269_ _06274_ _06330_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_132_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21300_ _08155_ _08156_ _08149_ _08153_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__a211o_1
X_22280_ _09022_ _09023_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__or2_1
XFILLER_178_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_130_Left_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21231_ _08074_ _08096_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__nand2_1
XFILLER_117_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21162_ systolic_inst.A_outs\[4\]\[5\] _11271_ _07850_ VGND VGND VPWR VPWR _08031_
+ sky130_fd_sc_hd__o21a_1
XFILLER_105_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20113_ _07087_ _07090_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__or2_1
XFILLER_160_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21093_ systolic_inst.A_outs\[4\]\[3\] _11271_ _07850_ VGND VGND VPWR VPWR _07964_
+ sky130_fd_sc_hd__o21ai_1
X_25970_ systolic_inst.acc_wires\[13\]\[30\] ser_C.parallel_data\[446\] net26 VGND
+ VGND VPWR VPWR _03272_ sky130_fd_sc_hd__mux2_1
XFILLER_131_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20044_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[6\]\[5\]
+ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_126_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24921_ C_out\[287\] net103 net75 ser_C.shift_reg\[287\] _10930_ VGND VGND VPWR VPWR
+ _02537_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27640_ clknet_leaf_316_clk _01438_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24852_ net113 ser_C.shift_reg\[254\] VGND VGND VPWR VPWR _10896_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23803_ _10401_ _10402_ VGND VGND VPWR VPWR _10404_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27571_ clknet_leaf_304_clk _01369_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_236_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _08774_ _08775_ _08776_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__nand3_1
X_24783_ C_out\[218\] net98 net78 ser_C.shift_reg\[218\] _10861_ VGND VGND VPWR VPWR
+ _02468_ sky130_fd_sc_hd__a221o_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29310_ clknet_leaf_302_clk _03108_ net141 VGND VGND VPWR VPWR C_out\[282\] sky130_fd_sc_hd__dfrtp_1
X_26522_ clknet_leaf_4_A_in_serial_clk _00325_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_23734_ _10344_ VGND VGND VPWR VPWR _10345_ sky130_fd_sc_hd__inv_2
XFILLER_96_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20946_ _07784_ _07819_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__xnor2_1
XFILLER_214_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_232_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_232_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29241_ clknet_leaf_176_clk _03039_ net148 VGND VGND VPWR VPWR C_out\[213\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26453_ clknet_leaf_346_clk _00260_ net132 VGND VGND VPWR VPWR A_in\[121\] sky130_fd_sc_hd__dfrtp_1
XFILLER_214_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23665_ _10283_ VGND VGND VPWR VPWR _10284_ sky130_fd_sc_hd__inv_2
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20877_ _07741_ _07753_ VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__nor2_1
XFILLER_242_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25404_ _11171_ systolic_inst.A_shift\[1\]\[1\] net71 VGND VGND VPWR VPWR _02779_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22616_ _09327_ _09328_ _09329_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__or3_1
XFILLER_224_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29172_ clknet_leaf_42_clk _02970_ net141 VGND VGND VPWR VPWR C_out\[144\] sky130_fd_sc_hd__dfrtp_1
X_23596_ _10215_ _10216_ VGND VGND VPWR VPWR _10218_ sky130_fd_sc_hd__nor2_1
X_26384_ clknet_leaf_14_clk _00191_ net133 VGND VGND VPWR VPWR A_in\[52\] sky130_fd_sc_hd__dfrtp_1
XFILLER_195_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28123_ clknet_leaf_125_clk _01921_ net144 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22547_ _09248_ _09271_ _09261_ _09270_ VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__o2bb2a_1
X_25335_ ser_C.parallel_data\[494\] net97 net77 ser_C.shift_reg\[494\] _11137_ VGND
+ VGND VPWR VPWR _02744_ sky130_fd_sc_hd__a221o_1
XFILLER_182_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28054_ clknet_leaf_51_clk _01852_ net143 VGND VGND VPWR VPWR systolic_inst.B_outs\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_10_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13280_ deser_A.word_buffer\[118\] deser_A.serial_word\[118\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__mux2_1
X_22478_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[2\]\[2\]
+ VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__nand2_1
XFILLER_212_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25266_ net111 ser_C.shift_reg\[461\] VGND VGND VPWR VPWR _11103_ sky130_fd_sc_hd__and2_1
XFILLER_108_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27005_ clknet_leaf_15_B_in_serial_clk _00803_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_21429_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[26\]
+ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__nand2_1
XFILLER_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24217_ systolic_inst.A_shift\[20\]\[0\] A_in\[72\] net59 VGND VGND VPWR VPWR _10594_
+ sky130_fd_sc_hd__mux2_1
X_25197_ C_out\[425\] net102 net74 ser_C.shift_reg\[425\] _11068_ VGND VGND VPWR VPWR
+ _02675_ sky130_fd_sc_hd__a221o_1
XFILLER_120_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24148_ _10575_ systolic_inst.A_shift\[28\]\[5\] net71 VGND VGND VPWR VPWR _02119_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24079_ systolic_inst.B_shift\[3\]\[6\] _11332_ net83 systolic_inst.B_shift\[7\]\[6\]
+ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__a22o_1
X_28956_ clknet_leaf_259_clk _02754_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[504\]
+ sky130_fd_sc_hd__dfrtp_1
X_16970_ net118 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[11\]\[0\]
+ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__a21oi_1
XFILLER_77_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27907_ clknet_leaf_136_clk _01705_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_15921_ _12940_ _12942_ _12944_ VGND VGND VPWR VPWR _12946_ sky130_fd_sc_hd__o21ai_1
XFILLER_103_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28887_ clknet_leaf_331_clk _02685_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[435\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18640_ systolic_inst.B_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[6\] systolic_inst.A_outs\[8\]\[7\]
+ systolic_inst.B_outs\[8\]\[3\] VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__a22o_1
XFILLER_231_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27838_ clknet_leaf_207_clk _01636_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_15852_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[15\]
+ VGND VGND VPWR VPWR _12887_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_177_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _11905_ _11908_ _11926_ VGND VGND VPWR VPWR _11929_ sky130_fd_sc_hd__nand3_1
XFILLER_92_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18571_ systolic_inst.B_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[4\]
+ systolic_inst.A_outs\[8\]\[5\] VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__and4_1
X_27769_ clknet_leaf_207_clk _01567_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_15783_ _12821_ _12822_ _12820_ VGND VGND VPWR VPWR _12828_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29508_ clknet_leaf_272_clk _03306_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17522_ _04746_ _04773_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__nand2b_1
X_14734_ _11877_ _11880_ VGND VGND VPWR VPWR _11882_ sky130_fd_sc_hd__or2_1
XFILLER_217_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29439_ clknet_leaf_332_clk _03237_ net131 VGND VGND VPWR VPWR C_out\[411\] sky130_fd_sc_hd__dfrtp_1
X_17453_ net118 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[11\] VGND
+ VGND VPWR VPWR _04707_ sky130_fd_sc_hd__or2_1
X_14665_ _11801_ _11822_ VGND VGND VPWR VPWR _11823_ sky130_fd_sc_hd__nor2_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16404_ _03774_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__inv_2
XFILLER_189_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13616_ deser_B.word_buffer\[52\] deser_B.serial_word\[52\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__mux2_1
XFILLER_158_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17384_ _04602_ _04639_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__nor2_1
X_14596_ _11757_ _11763_ VGND VGND VPWR VPWR _11764_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_215_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19123_ _06159_ _06188_ _06189_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__nand3_1
X_16335_ _11260_ systolic_inst.A_outs\[12\]\[7\] _03664_ _03689_ VGND VGND VPWR VPWR
+ _03714_ sky130_fd_sc_hd__o211ai_1
X_13547_ deser_A.shift_reg\[111\] deser_A.shift_reg\[112\] net129 VGND VGND VPWR VPWR
+ _00384_ sky130_fd_sc_hd__mux2_1
XFILLER_9_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19054_ net105 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[3\] VGND
+ VGND VPWR VPWR _06124_ sky130_fd_sc_hd__nand2_1
X_16266_ _03647_ _03646_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__and2b_1
XFILLER_139_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13478_ deser_A.shift_reg\[42\] deser_A.shift_reg\[43\] net130 VGND VGND VPWR VPWR
+ _00315_ sky130_fd_sc_hd__mux2_1
XFILLER_195_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18005_ systolic_inst.A_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[6\]
+ systolic_inst.B_outs\[9\]\[7\] VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__and4b_1
X_15217_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[14\]\[11\]
+ VGND VGND VPWR VPWR _12320_ sky130_fd_sc_hd__nor2_1
XFILLER_103_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16197_ _03555_ _03580_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15148_ net118 _12260_ _12261_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_236_Right_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19956_ systolic_inst.A_outs\[6\]\[6\] _11278_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__or2_1
X_15079_ _12141_ _12195_ VGND VGND VPWR VPWR _12197_ sky130_fd_sc_hd__xor2_1
XFILLER_141_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18907_ _05997_ _06003_ _06011_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__a21o_1
XFILLER_228_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19887_ _06813_ _06847_ _06848_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__o21ba_1
XFILLER_228_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18838_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[8\]\[6\]
+ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__or2_1
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18769_ systolic_inst.B_outs\[8\]\[5\] systolic_inst.A_outs\[8\]\[7\] _05868_ _05867_
+ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__a31o_1
XFILLER_110_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
X_20800_ _07700_ _07701_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__xnor2_1
X_21780_ _08583_ _08584_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__nand2_2
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20731_ _07641_ _07642_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__nor2_1
XFILLER_24_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23450_ systolic_inst.B_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[5\]
+ systolic_inst.B_outs\[0\]\[3\] VGND VGND VPWR VPWR _10075_ sky130_fd_sc_hd__a22oi_1
XFILLER_149_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20662_ _07584_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__inv_2
XFILLER_177_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22401_ _09141_ _09140_ VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__and2b_1
XFILLER_52_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23381_ _10002_ _10007_ VGND VGND VPWR VPWR _10008_ sky130_fd_sc_hd__xnor2_1
X_20593_ systolic_inst.B_outs\[5\]\[5\] systolic_inst.B_outs\[5\]\[6\] systolic_inst.A_outs\[5\]\[7\]
+ _07523_ VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__a31o_1
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22332_ _09073_ _09074_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__nand2b_1
XFILLER_192_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25120_ net110 ser_C.shift_reg\[388\] VGND VGND VPWR VPWR _11030_ sky130_fd_sc_hd__and2_1
XFILLER_17_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25051_ C_out\[352\] net97 net77 ser_C.shift_reg\[352\] _10995_ VGND VGND VPWR VPWR
+ _02602_ sky130_fd_sc_hd__a221o_1
X_22263_ _08989_ _09006_ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__xor2_1
XFILLER_117_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24002_ _10526_ systolic_inst.B_shift\[5\]\[4\] _11332_ VGND VGND VPWR VPWR _02022_
+ sky130_fd_sc_hd__mux2_1
X_21214_ _08028_ _08080_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_225_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22194_ _08908_ _08910_ _08939_ _08940_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_225_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_203_Right_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28810_ clknet_leaf_244_clk _02608_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[358\]
+ sky130_fd_sc_hd__dfrtp_1
X_21145_ _07997_ _08014_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__xor2_1
XFILLER_219_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_221_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_221_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28741_ clknet_leaf_296_clk _02539_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[289\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25953_ systolic_inst.acc_wires\[13\]\[13\] C_out\[429\] net19 VGND VGND VPWR VPWR
+ _03255_ sky130_fd_sc_hd__mux2_1
XFILLER_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21076_ _07947_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_238_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20027_ _07014_ _07015_ _07016_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__and3_1
X_24904_ net110 ser_C.shift_reg\[280\] VGND VGND VPWR VPWR _10922_ sky130_fd_sc_hd__and2_1
X_28672_ clknet_leaf_184_clk _02470_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25884_ systolic_inst.acc_wires\[11\]\[8\] C_out\[360\] net39 VGND VGND VPWR VPWR
+ _03186_ sky130_fd_sc_hd__mux2_1
XFILLER_86_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27623_ clknet_leaf_317_clk _01421_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_24835_ C_out\[244\] net98 net78 ser_C.shift_reg\[244\] _10887_ VGND VGND VPWR VPWR
+ _02494_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_38_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_189_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27554_ clknet_leaf_304_clk _01352_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24766_ net113 ser_C.shift_reg\[211\] VGND VGND VPWR VPWR _10853_ sky130_fd_sc_hd__and2_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21978_ _08762_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__inv_2
XFILLER_226_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26505_ clknet_leaf_16_A_in_serial_clk _00308_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23717_ _10323_ _10324_ _10322_ VGND VGND VPWR VPWR _10330_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_29_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27485_ clknet_leaf_296_clk _01283_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_20929_ systolic_inst.A_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\] VGND VGND VPWR
+ VPWR _07804_ sky130_fd_sc_hd__nand2_1
X_24697_ C_out\[175\] net104 net76 ser_C.shift_reg\[175\] _10818_ VGND VGND VPWR VPWR
+ _02425_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_29_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29224_ clknet_leaf_211_clk _03022_ net147 VGND VGND VPWR VPWR C_out\[196\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26436_ clknet_leaf_4_clk _00243_ net131 VGND VGND VPWR VPWR A_in\[104\] sky130_fd_sc_hd__dfrtp_1
X_14450_ _11600_ _11602_ _11631_ VGND VGND VPWR VPWR _11632_ sky130_fd_sc_hd__a21o_1
X_23648_ systolic_inst.A_outs\[0\]\[6\] _10195_ _10154_ VGND VGND VPWR VPWR _10268_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_186_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13401_ A_in\[110\] deser_A.word_buffer\[110\] net95 VGND VGND VPWR VPWR _00249_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_226_Left_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29155_ clknet_leaf_168_clk _02953_ net148 VGND VGND VPWR VPWR C_out\[127\] sky130_fd_sc_hd__dfrtp_1
XFILLER_186_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14381_ _11561_ _11564_ VGND VGND VPWR VPWR _11565_ sky130_fd_sc_hd__xnor2_1
X_26367_ clknet_leaf_26_clk _00174_ net137 VGND VGND VPWR VPWR A_in\[35\] sky130_fd_sc_hd__dfrtp_1
X_23579_ _10199_ _10200_ VGND VGND VPWR VPWR _10201_ sky130_fd_sc_hd__and2_1
XFILLER_22_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28106_ clknet_leaf_156_clk _01904_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16120_ _13085_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__nand2b_1
XFILLER_122_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25318_ net112 ser_C.shift_reg\[487\] VGND VGND VPWR VPWR _11129_ sky130_fd_sc_hd__and2_1
X_13332_ A_in\[41\] deser_A.word_buffer\[41\] net93 VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__mux2_1
X_29086_ clknet_leaf_111_clk _02884_ net151 VGND VGND VPWR VPWR C_out\[58\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_210_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26298_ clknet_leaf_22_A_in_serial_clk _00106_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_210_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28037_ clknet_leaf_159_clk _01835_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16051_ _13016_ _13046_ VGND VGND VPWR VPWR _13048_ sky130_fd_sc_hd__or2_1
X_25249_ ser_C.parallel_data\[451\] net102 net74 ser_C.shift_reg\[451\] _11094_ VGND
+ VGND VPWR VPWR _02701_ sky130_fd_sc_hd__a221o_1
X_13263_ deser_A.word_buffer\[101\] deser_A.serial_word\[101\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15002_ _12120_ _12121_ VGND VGND VPWR VPWR _12122_ sky130_fd_sc_hd__nand2_1
X_13194_ deser_A.word_buffer\[32\] deser_A.serial_word\[32\] net127 VGND VGND VPWR
+ VPWR _00042_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19810_ _06779_ _06809_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__xor2_1
XFILLER_151_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_235_Left_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19741_ _06720_ _06722_ _06721_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__o21ba_1
X_16953_ _04198_ _04267_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28939_ clknet_leaf_260_clk _02737_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15904_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[23\]
+ VGND VGND VPWR VPWR _12931_ sky130_fd_sc_hd__xor2_1
X_19672_ _06675_ _06676_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__or2_1
XFILLER_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16884_ systolic_inst.B_outs\[11\]\[6\] systolic_inst.A_outs\[11\]\[6\] _11262_ systolic_inst.A_outs\[11\]\[5\]
+ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_238_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18623_ _05748_ _05749_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__xor2_1
X_15835_ net108 systolic_inst.acc_wires\[13\]\[12\] net67 _12872_ VGND VGND VPWR VPWR
+ _01118_ sky130_fd_sc_hd__a22o_1
XFILLER_92_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_218_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18554_ _05681_ _05682_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__xnor2_1
X_15766_ net66 _12811_ _12813_ systolic_inst.acc_wires\[13\]\[2\] net107 VGND VGND
+ VPWR VPWR _01108_ sky130_fd_sc_hd__a32o_1
XFILLER_209_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17505_ _04757_ _04756_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__and2b_1
X_14717_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[28\]
+ VGND VGND VPWR VPWR _11867_ sky130_fd_sc_hd__or2_1
XFILLER_178_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18485_ _05594_ _05616_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__nand2_1
XFILLER_127_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15697_ _12720_ _12748_ VGND VGND VPWR VPWR _12750_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17436_ _04689_ _04690_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__nand2b_1
XFILLER_220_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14648_ _11806_ _11808_ VGND VGND VPWR VPWR _11809_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_155_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_221_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_17 net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_28 systolic_inst.A_outs\[8\]\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17367_ _04606_ _04623_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__or2_1
XFILLER_14_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14579_ net69 _11748_ _11749_ systolic_inst.acc_wires\[15\]\[7\] net105 VGND VGND
+ VPWR VPWR _00985_ sky130_fd_sc_hd__a32o_1
XFILLER_105_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19106_ _06172_ _06169_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__and2b_1
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16318_ _03632_ _03696_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__or2_1
X_17298_ _04554_ _04555_ _04523_ _04525_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_168_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19037_ _06105_ _06106_ _06101_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__or3b_1
XFILLER_173_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16249_ _03594_ _03630_ systolic_inst.A_outs\[12\]\[7\] VGND VGND VPWR VPWR _03631_
+ sky130_fd_sc_hd__and3b_1
XFILLER_161_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19939_ _06934_ _06935_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__nand2_1
XFILLER_102_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22950_ systolic_inst.B_outs\[1\]\[5\] systolic_inst.A_outs\[1\]\[6\] VGND VGND VPWR
+ VPWR _09628_ sky130_fd_sc_hd__nand2_1
XFILLER_229_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21901_ _08695_ _08696_ _08688_ _08692_ VGND VGND VPWR VPWR _08697_ sky130_fd_sc_hd__a211o_1
XFILLER_56_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap19 net20 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_8
X_22881_ _09557_ _09560_ VGND VGND VPWR VPWR _09561_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_69_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24620_ net110 ser_C.shift_reg\[138\] VGND VGND VPWR VPWR _10780_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21832_ _08602_ _08604_ _08634_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__o21a_1
XFILLER_24_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24551_ C_out\[102\] net99 net79 ser_C.shift_reg\[102\] _10745_ VGND VGND VPWR VPWR
+ _02352_ sky130_fd_sc_hd__a221o_1
X_21763_ _08567_ _08568_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20714_ _07627_ _07628_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__and2_1
X_23502_ _10123_ _10124_ VGND VGND VPWR VPWR _10126_ sky130_fd_sc_hd__xnor2_1
X_27270_ clknet_leaf_267_clk _01068_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_24482_ net112 ser_C.shift_reg\[69\] VGND VGND VPWR VPWR _10711_ sky130_fd_sc_hd__and2_1
X_21694_ _08484_ _08501_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__xor2_1
XFILLER_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26221_ clknet_leaf_8_A_in_serial_clk _00029_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_23433_ _10015_ _10017_ _10056_ _10057_ VGND VGND VPWR VPWR _10059_ sky130_fd_sc_hd__a211o_1
X_20645_ _07563_ _07564_ _07562_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_24_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_227_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26152_ deser_B.serial_word\[107\] deser_B.shift_reg\[107\] _00001_ VGND VGND VPWR
+ VPWR _03454_ sky130_fd_sc_hd__mux2_1
X_23364_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[5\]
+ systolic_inst.A_outs\[0\]\[6\] VGND VGND VPWR VPWR _09991_ sky130_fd_sc_hd__and4_1
X_20576_ _07465_ _07507_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_227_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25103_ C_out\[378\] net98 net78 ser_C.shift_reg\[378\] _11021_ VGND VGND VPWR VPWR
+ _02628_ sky130_fd_sc_hd__a221o_1
X_22315_ _09056_ _09057_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__or2_1
XFILLER_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26083_ deser_B.serial_word\[38\] deser_B.shift_reg\[38\] net55 VGND VGND VPWR VPWR
+ _03385_ sky130_fd_sc_hd__mux2_1
XFILLER_192_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23295_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[2\] _09922_ _09923_
+ VGND VGND VPWR VPWR _09926_ sky130_fd_sc_hd__a22oi_1
XFILLER_164_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22246_ systolic_inst.B_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[5\]
+ systolic_inst.B_outs\[2\]\[3\] VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__a22oi_1
XFILLER_180_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25034_ net112 ser_C.shift_reg\[345\] VGND VGND VPWR VPWR _10987_ sky130_fd_sc_hd__and2_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22177_ systolic_inst.B_outs\[2\]\[3\] systolic_inst.A_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\]
+ systolic_inst.A_outs\[2\]\[2\] VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__a22o_1
XFILLER_191_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21128_ systolic_inst.B_outs\[4\]\[5\] systolic_inst.A_outs\[4\]\[6\] systolic_inst.A_outs\[4\]\[7\]
+ systolic_inst.B_outs\[4\]\[1\] VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__a22o_1
XFILLER_105_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26985_ clknet_leaf_0_A_in_serial_clk _00783_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28724_ clknet_leaf_312_clk _02522_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[272\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21059_ _07927_ _07930_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__xnor2_1
X_25936_ systolic_inst.acc_wires\[12\]\[28\] C_out\[412\] net21 VGND VGND VPWR VPWR
+ _03238_ sky130_fd_sc_hd__mux2_1
X_13950_ deser_A.serial_word\[111\] deser_A.shift_reg\[111\] net57 VGND VGND VPWR
+ VPWR _00776_ sky130_fd_sc_hd__mux2_1
XFILLER_4_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28655_ clknet_leaf_204_clk _02453_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[203\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13881_ deser_A.serial_word\[42\] deser_A.shift_reg\[42\] net58 VGND VGND VPWR VPWR
+ _00707_ sky130_fd_sc_hd__mux2_1
X_25867_ systolic_inst.acc_wires\[10\]\[23\] C_out\[343\] net11 VGND VGND VPWR VPWR
+ _03169_ sky130_fd_sc_hd__mux2_1
XFILLER_35_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27606_ clknet_leaf_203_clk _01404_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_28_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15620_ _12608_ _12640_ _12675_ VGND VGND VPWR VPWR _12676_ sky130_fd_sc_hd__a21o_1
X_24818_ net113 ser_C.shift_reg\[237\] VGND VGND VPWR VPWR _10879_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28586_ clknet_leaf_308_clk _02384_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[134\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_195_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25798_ systolic_inst.acc_wires\[8\]\[18\] C_out\[274\] net22 VGND VGND VPWR VPWR
+ _03100_ sky130_fd_sc_hd__mux2_1
X_15551_ _12606_ _12607_ VGND VGND VPWR VPWR _12609_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27537_ clknet_leaf_317_clk _01335_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_226_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24749_ C_out\[201\] net97 net80 ser_C.shift_reg\[201\] _10844_ VGND VGND VPWR VPWR
+ _02451_ sky130_fd_sc_hd__a221o_1
XFILLER_188_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_191_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14502_ _11680_ _11681_ VGND VGND VPWR VPWR _11682_ sky130_fd_sc_hd__nand2_1
XFILLER_230_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[9\]\[10\]
+ _05434_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__and3_1
XFILLER_15_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15482_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[6\]
+ systolic_inst.A_outs\[13\]\[7\] VGND VGND VPWR VPWR _12541_ sky130_fd_sc_hd__nand4_1
X_27468_ clknet_leaf_297_clk _01266_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_212_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29207_ clknet_leaf_205_clk _03005_ net146 VGND VGND VPWR VPWR C_out\[179\] sky130_fd_sc_hd__dfrtp_1
X_17221_ _04468_ _04471_ _04481_ _04482_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__a211o_1
X_14433_ _11613_ _11614_ VGND VGND VPWR VPWR _11616_ sky130_fd_sc_hd__or2_1
XFILLER_74_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26419_ clknet_leaf_6_clk _00226_ net133 VGND VGND VPWR VPWR A_in\[87\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27399_ clknet_leaf_332_clk _01197_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29138_ clknet_leaf_167_clk _02936_ net148 VGND VGND VPWR VPWR C_out\[110\] sky130_fd_sc_hd__dfrtp_1
X_17152_ net105 systolic_inst.acc_wires\[11\]\[27\] net62 _04437_ VGND VGND VPWR VPWR
+ _01261_ sky130_fd_sc_hd__a22o_1
XFILLER_122_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14364_ _11546_ _11548_ VGND VGND VPWR VPWR _11549_ sky130_fd_sc_hd__or2_1
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16103_ _13096_ _13097_ VGND VGND VPWR VPWR _13098_ sky130_fd_sc_hd__or2_1
XFILLER_183_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13315_ A_in\[24\] deser_A.word_buffer\[24\] net91 VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__mux2_1
XFILLER_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29069_ clknet_leaf_118_clk _02867_ net152 VGND VGND VPWR VPWR C_out\[41\] sky130_fd_sc_hd__dfrtp_1
X_17083_ net60 _04379_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__nor2_1
X_14295_ _11476_ _11480_ VGND VGND VPWR VPWR _11481_ sky130_fd_sc_hd__xnor2_1
X_16034_ _13030_ _13027_ VGND VGND VPWR VPWR _13031_ sky130_fd_sc_hd__nand2b_1
X_13246_ deser_A.word_buffer\[84\] deser_A.serial_word\[84\] net127 VGND VGND VPWR
+ VPWR _00094_ sky130_fd_sc_hd__mux2_1
XFILLER_124_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13177_ deser_A.word_buffer\[15\] deser_A.serial_word\[15\] net128 VGND VGND VPWR
+ VPWR _00025_ sky130_fd_sc_hd__mux2_1
XFILLER_123_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17985_ _05146_ _05176_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__xor2_1
XFILLER_97_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19724_ _06693_ _06726_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_144_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16936_ _04250_ _04251_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__xor2_1
XFILLER_238_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19655_ _06659_ _06660_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__and2b_1
X_16867_ _04184_ _04183_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_0_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15818_ _12855_ _12857_ VGND VGND VPWR VPWR _12858_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18606_ _05732_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__or2_1
X_19586_ net106 systolic_inst.acc_wires\[7\]\[27\] net62 _06615_ VGND VGND VPWR VPWR
+ _01517_ sky130_fd_sc_hd__a22o_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16798_ _04117_ _04116_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_103_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18537_ systolic_inst.A_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\] systolic_inst.A_outs\[8\]\[4\]
+ systolic_inst.B_outs\[8\]\[3\] VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__a22oi_1
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15749_ net108 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] _12792_
+ _12799_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__a22o_1
XFILLER_234_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18468_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[4\] _05600_
+ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__a21bo_1
XFILLER_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17419_ _04672_ _04673_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__or2_1
XFILLER_18_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18399_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[31\]
+ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20430_ systolic_inst.B_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[5\]
+ systolic_inst.A_outs\[5\]\[6\] VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__and4_1
XFILLER_105_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload220 clknet_leaf_53_clk VGND VGND VPWR VPWR clkload220/Y sky130_fd_sc_hd__clkinv_4
X_20361_ _07297_ _07298_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__and2b_1
XFILLER_88_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload231 clknet_leaf_78_clk VGND VGND VPWR VPWR clkload231/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
Xclkload242 clknet_leaf_79_clk VGND VGND VPWR VPWR clkload242/Y sky130_fd_sc_hd__clkinv_4
XFILLER_88_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22100_ net109 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _08851_ sky130_fd_sc_hd__and2_1
Xclkload253 clknet_leaf_92_clk VGND VGND VPWR VPWR clkload253/Y sky130_fd_sc_hd__inv_6
Xclkbuf_5_15__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_15__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xclkload264 clknet_leaf_107_clk VGND VGND VPWR VPWR clkload264/Y sky130_fd_sc_hd__clkinv_4
X_23080_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[1\]\[0\]
+ _09745_ _09743_ VGND VGND VPWR VPWR _09751_ sky130_fd_sc_hd__a31o_1
XFILLER_179_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload275 clknet_leaf_143_clk VGND VGND VPWR VPWR clkload275/Y sky130_fd_sc_hd__clkinv_2
X_20292_ _07228_ _07231_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__xor2_1
Xclkload286 clknet_leaf_190_clk VGND VGND VPWR VPWR clkload286/Y sky130_fd_sc_hd__inv_6
Xclkload297 clknet_leaf_177_clk VGND VGND VPWR VPWR clkload297/Y sky130_fd_sc_hd__clkinv_8
X_22031_ _08806_ _08807_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__or2_1
XFILLER_114_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26770_ clknet_leaf_95_clk _00572_ net5 VGND VGND VPWR VPWR B_in\[42\] sky130_fd_sc_hd__dfrtp_1
X_23982_ _10516_ systolic_inst.B_shift\[8\]\[2\] net72 VGND VGND VPWR VPWR _02012_
+ sky130_fd_sc_hd__mux2_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25721_ systolic_inst.acc_wires\[6\]\[5\] C_out\[197\] net11 VGND VGND VPWR VPWR
+ _03023_ sky130_fd_sc_hd__mux2_1
XFILLER_112_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22933_ _09554_ _09610_ VGND VGND VPWR VPWR _09612_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28440_ clknet_leaf_35_clk _02238_ VGND VGND VPWR VPWR systolic_inst.A_shift\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_216_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25652_ systolic_inst.acc_wires\[4\]\[0\] C_out\[128\] net28 VGND VGND VPWR VPWR
+ _02954_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_216_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22864_ _09503_ _09505_ VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__nor2_1
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24603_ C_out\[128\] net103 net75 ser_C.shift_reg\[128\] _10771_ VGND VGND VPWR VPWR
+ _02378_ sky130_fd_sc_hd__a221o_1
X_21815_ _08590_ _08617_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__xnor2_1
X_28371_ clknet_leaf_5_clk _02169_ VGND VGND VPWR VPWR systolic_inst.A_shift\[20\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25583_ systolic_inst.acc_wires\[1\]\[27\] C_out\[59\] net52 VGND VGND VPWR VPWR
+ _02885_ sky130_fd_sc_hd__mux2_1
XFILLER_197_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22795_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[6\] _09477_ net122
+ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__mux2_1
XFILLER_52_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27322_ clknet_leaf_329_clk _01120_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24534_ net114 ser_C.shift_reg\[95\] VGND VGND VPWR VPWR _10737_ sky130_fd_sc_hd__and2_1
X_21746_ _08443_ _08550_ VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__nand2_1
XFILLER_169_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27253_ clknet_leaf_281_clk _01051_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24465_ C_out\[59\] net100 net82 ser_C.shift_reg\[59\] _10702_ VGND VGND VPWR VPWR
+ _02309_ sky130_fd_sc_hd__a221o_1
XFILLER_185_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21677_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[7\] VGND VGND VPWR
+ VPWR _08485_ sky130_fd_sc_hd__nand2_4
XFILLER_8_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26204_ clknet_leaf_14_A_in_serial_clk _00012_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_23416_ _10040_ _10041_ VGND VGND VPWR VPWR _10042_ sky130_fd_sc_hd__nor2_1
X_20628_ net63 _07554_ _07555_ systolic_inst.acc_wires\[5\]\[1\] net109 VGND VGND
+ VPWR VPWR _01619_ sky130_fd_sc_hd__a32o_1
X_27184_ clknet_leaf_261_clk _00982_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24396_ net7 ser_C.shift_reg\[26\] VGND VGND VPWR VPWR _10668_ sky130_fd_sc_hd__and2_1
XFILLER_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26135_ deser_B.serial_word\[90\] deser_B.shift_reg\[90\] net56 VGND VGND VPWR VPWR
+ _03437_ sky130_fd_sc_hd__mux2_1
X_20559_ _07489_ _07490_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__and2_1
X_23347_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[3\]
+ systolic_inst.A_outs\[0\]\[4\] VGND VGND VPWR VPWR _09975_ sky130_fd_sc_hd__and4_1
XFILLER_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14080_ deser_B.shift_reg\[114\] deser_B.shift_reg\[115\] deser_B.receiving VGND
+ VGND VPWR VPWR _00906_ sky130_fd_sc_hd__mux2_1
X_26066_ deser_B.serial_word\[21\] deser_B.shift_reg\[21\] net55 VGND VGND VPWR VPWR
+ _03368_ sky130_fd_sc_hd__mux2_1
X_23278_ systolic_inst.A_outs\[0\]\[1\] systolic_inst.A_shift\[0\]\[1\] net121 VGND
+ VGND VPWR VPWR _01907_ sky130_fd_sc_hd__mux2_1
XFILLER_106_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25017_ C_out\[335\] net97 net80 ser_C.shift_reg\[335\] _10978_ VGND VGND VPWR VPWR
+ _02585_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_56_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22229_ _08946_ _08974_ VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_56_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_205_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_205_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_205_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17770_ _04983_ _04986_ _04985_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__o21a_1
XFILLER_232_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14982_ _12061_ _12067_ _12101_ net107 VGND VGND VPWR VPWR _12103_ sky130_fd_sc_hd__a31o_1
X_26968_ clknet_leaf_24_A_in_serial_clk _00766_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_201_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_197_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16721_ _04026_ _04042_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__xnor2_1
X_28707_ clknet_leaf_190_clk _02505_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[255\]
+ sky130_fd_sc_hd__dfrtp_1
X_25919_ systolic_inst.acc_wires\[12\]\[11\] C_out\[395\] net18 VGND VGND VPWR VPWR
+ _03221_ sky130_fd_sc_hd__mux2_1
XFILLER_43_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13933_ deser_A.serial_word\[94\] deser_A.shift_reg\[94\] net57 VGND VGND VPWR VPWR
+ _00759_ sky130_fd_sc_hd__mux2_1
XFILLER_93_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29687_ clknet_leaf_105_clk _03482_ net151 VGND VGND VPWR VPWR ser_C.bit_idx\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_26899_ clknet_leaf_12_A_in_serial_clk _00697_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19440_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[7\]\[6\]
+ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_193_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28638_ clknet_leaf_179_clk _02436_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[186\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16652_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[5\] _03973_ _03974_
+ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_234_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_193_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13864_ deser_A.serial_word\[25\] deser_A.shift_reg\[25\] net58 VGND VGND VPWR VPWR
+ _00690_ sky130_fd_sc_hd__mux2_1
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15603_ _12650_ _12658_ VGND VGND VPWR VPWR _12659_ sky130_fd_sc_hd__nand2_1
XFILLER_90_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19371_ systolic_inst.B_outs\[7\]\[5\] systolic_inst.A_outs\[7\]\[7\] _06408_ _06407_
+ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__a31o_1
XFILLER_234_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28569_ clknet_leaf_175_clk _02367_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16583_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[6\]\[0\] net120 VGND
+ VGND VPWR VPWR _01210_ sky130_fd_sc_hd__mux2_1
X_13795_ B_in\[102\] deser_B.word_buffer\[102\] _00005_ VGND VGND VPWR VPWR _00632_
+ sky130_fd_sc_hd__mux2_1
XFILLER_222_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18322_ _05480_ _05484_ _05486_ net60 VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__a31o_1
XFILLER_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15534_ systolic_inst.A_outs\[13\]\[2\] systolic_inst.B_outs\[13\]\[5\] _12555_ _12554_
+ VGND VGND VPWR VPWR _12592_ sky130_fd_sc_hd__a31o_1
XFILLER_163_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18253_ net66 _05427_ _05428_ systolic_inst.acc_wires\[9\]\[9\] net107 VGND VGND
+ VPWR VPWR _01371_ sky130_fd_sc_hd__a32o_1
XFILLER_15_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15465_ _12494_ _12523_ _12524_ VGND VGND VPWR VPWR _12525_ sky130_fd_sc_hd__and3_1
X_17204_ _04464_ _04465_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__a21o_1
X_14416_ _11561_ _11563_ _11562_ VGND VGND VPWR VPWR _11599_ sky130_fd_sc_hd__o21ba_1
XFILLER_175_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18184_ _05149_ _05288_ _05361_ _05359_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__a31o_1
X_15396_ _12452_ _12457_ VGND VGND VPWR VPWR _12459_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17135_ _04418_ _04420_ _04423_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__a21oi_2
X_14347_ _11529_ _11530_ VGND VGND VPWR VPWR _11532_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17066_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[11\]\[13\]
+ _04359_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__a21oi_1
X_14278_ _11421_ _11423_ VGND VGND VPWR VPWR _11465_ sky130_fd_sc_hd__and2b_1
XFILLER_171_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16017_ _12994_ _13013_ VGND VGND VPWR VPWR _13015_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13229_ deser_A.word_buffer\[67\] deser_A.serial_word\[67\] net127 VGND VGND VPWR
+ VPWR _00077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_260_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_260_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_135_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17968_ systolic_inst.A_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[2\] systolic_inst.B_outs\[9\]\[6\]
+ systolic_inst.B_outs\[9\]\[7\] VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_105_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19707_ _06708_ _06709_ net120 VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__o21a_1
XFILLER_22_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16919_ _04232_ _04233_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__xnor2_1
X_17899_ _05059_ _05093_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__nor2_1
XFILLER_225_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19638_ _06644_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__inv_2
XFILLER_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19569_ _06596_ _06598_ _06601_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__a21oi_2
XFILLER_41_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21600_ _08404_ _08408_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__and2_1
XFILLER_146_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22580_ _09298_ _09299_ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_1085 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21531_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[4\] _08343_
+ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__a21bo_1
XFILLER_181_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21462_ _08289_ _08293_ _08294_ _11713_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__a31o_1
X_24250_ systolic_inst.A_shift\[17\]\[1\] net70 net83 systolic_inst.A_shift\[18\]\[1\]
+ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__a22o_1
XFILLER_147_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23201_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[20\]
+ VGND VGND VPWR VPWR _09854_ sky130_fd_sc_hd__nand2_1
XFILLER_222_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20413_ _07319_ _07349_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_96_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21393_ _08233_ _08236_ _08237_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__or3_1
X_24181_ systolic_inst.A_shift\[25\]\[4\] net70 _10505_ systolic_inst.A_shift\[26\]\[4\]
+ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23132_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[1\]\[10\]
+ VGND VGND VPWR VPWR _09795_ sky130_fd_sc_hd__or2_1
XFILLER_162_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20344_ _07281_ _07282_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_92_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27940_ clknet_leaf_170_clk _01738_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_23063_ _09653_ _09717_ VGND VGND VPWR VPWR _09737_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20275_ systolic_inst.A_outs\[5\]\[4\] _07215_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_241_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_241_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22014_ _08793_ _08792_ systolic_inst.acc_wires\[3\]\[21\] net106 VGND VGND VPWR
+ VPWR _01767_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_153_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27871_ clknet_leaf_309_clk _01669_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26822_ clknet_leaf_70_clk _00624_ net135 VGND VGND VPWR VPWR B_in\[94\] sky130_fd_sc_hd__dfrtp_1
X_29610_ clknet_leaf_28_B_in_serial_clk _03405_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_251_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_251_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_102_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29541_ clknet_leaf_105_clk _00009_ net152 VGND VGND VPWR VPWR systolic_inst.ce_local
+ sky130_fd_sc_hd__dfrtp_4
X_26753_ clknet_leaf_57_clk _00555_ net137 VGND VGND VPWR VPWR B_in\[25\] sky130_fd_sc_hd__dfrtp_1
X_23965_ systolic_inst.B_shift\[13\]\[2\] B_in\[42\] _00008_ VGND VGND VPWR VPWR _10508_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25704_ systolic_inst.acc_wires\[5\]\[20\] C_out\[180\] net45 VGND VGND VPWR VPWR
+ _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_1_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22916_ systolic_inst.A_outs\[1\]\[4\] systolic_inst.B_outs\[1\]\[6\] _11277_ systolic_inst.A_outs\[1\]\[3\]
+ VGND VGND VPWR VPWR _09595_ sky130_fd_sc_hd__o2bb2a_1
X_29472_ clknet_leaf_284_clk _03270_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[444\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26684_ clknet_leaf_28_B_in_serial_clk _00487_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23896_ systolic_inst.B_shift\[17\]\[0\] B_in\[72\] _00008_ VGND VGND VPWR VPWR _10481_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28423_ clknet_leaf_22_clk _02221_ VGND VGND VPWR VPWR systolic_inst.A_shift\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25635_ systolic_inst.acc_wires\[3\]\[15\] C_out\[111\] net51 VGND VGND VPWR VPWR
+ _02937_ sky130_fd_sc_hd__mux2_1
XFILLER_216_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22847_ systolic_inst.A_outs\[1\]\[2\] systolic_inst.B_outs\[1\]\[6\] _09526_ VGND
+ VGND VPWR VPWR _09528_ sky130_fd_sc_hd__and3_1
XFILLER_186_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28354_ clknet_leaf_342_clk _02152_ VGND VGND VPWR VPWR systolic_inst.A_shift\[24\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25566_ systolic_inst.acc_wires\[1\]\[10\] C_out\[42\] net36 VGND VGND VPWR VPWR
+ _02868_ sky130_fd_sc_hd__mux2_1
X_13580_ deser_B.word_buffer\[16\] deser_B.serial_word\[16\] net124 VGND VGND VPWR
+ VPWR _00417_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22778_ systolic_inst.A_outs\[1\]\[1\] systolic_inst.B_outs\[1\]\[6\] VGND VGND VPWR
+ VPWR _09461_ sky130_fd_sc_hd__nand2_1
XFILLER_231_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27305_ clknet_leaf_329_clk _01103_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_24517_ C_out\[85\] net100 net82 ser_C.shift_reg\[85\] _10728_ VGND VGND VPWR VPWR
+ _02335_ sky130_fd_sc_hd__a221o_1
XFILLER_212_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21729_ _08517_ _08535_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__xor2_1
X_28285_ clknet_leaf_57_clk _02083_ VGND VGND VPWR VPWR systolic_inst.B_shift\[19\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25497_ systolic_inst.cycle_cnt\[22\] systolic_inst.cycle_cnt\[21\] _11225_ VGND
+ VGND VPWR VPWR _11228_ sky130_fd_sc_hd__and3_1
XFILLER_157_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15250_ _12347_ _12348_ _12341_ _12345_ VGND VGND VPWR VPWR _12349_ sky130_fd_sc_hd__o211ai_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27236_ clknet_leaf_278_clk _01034_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24448_ net114 ser_C.shift_reg\[52\] VGND VGND VPWR VPWR _10694_ sky130_fd_sc_hd__and2_1
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14201_ _11387_ _11388_ _11389_ VGND VGND VPWR VPWR _11390_ sky130_fd_sc_hd__or3_1
XFILLER_240_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27167_ clknet_leaf_253_clk _00965_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15181_ _12280_ _12284_ _12287_ _12288_ VGND VGND VPWR VPWR _12290_ sky130_fd_sc_hd__o211a_1
X_24379_ C_out\[16\] net104 _10643_ ser_C.shift_reg\[16\] _10659_ VGND VGND VPWR VPWR
+ _02266_ sky130_fd_sc_hd__a221o_1
XFILLER_201_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26118_ deser_B.serial_word\[73\] deser_B.shift_reg\[73\] _00001_ VGND VGND VPWR
+ VPWR _03420_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14132_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[10\]\[0\] net120 VGND
+ VGND VPWR VPWR _00954_ sky130_fd_sc_hd__mux2_1
XFILLER_181_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27098_ clknet_leaf_7_B_in_serial_clk _00896_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_207_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26049_ deser_B.serial_word\[4\] deser_B.shift_reg\[4\] net55 VGND VGND VPWR VPWR
+ _03351_ sky130_fd_sc_hd__mux2_1
X_14063_ deser_B.shift_reg\[97\] deser_B.shift_reg\[98\] net126 VGND VGND VPWR VPWR
+ _00889_ sky130_fd_sc_hd__mux2_1
X_18940_ _06037_ _06039_ _06040_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_176_Left_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18871_ _05973_ _05976_ _05979_ net61 VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__a31o_1
XFILLER_80_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_242_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_242_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_141_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17822_ systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[3\]
+ systolic_inst.B_outs\[9\]\[0\] VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_141_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14965_ _12085_ _12084_ VGND VGND VPWR VPWR _12086_ sky130_fd_sc_hd__nand2b_1
XFILLER_94_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17753_ _04967_ _04969_ _04975_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__a21o_1
XFILLER_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13916_ deser_A.serial_word\[77\] deser_A.shift_reg\[77\] net57 VGND VGND VPWR VPWR
+ _00742_ sky130_fd_sc_hd__mux2_1
XFILLER_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16704_ _03990_ _04025_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17684_ _04901_ _04908_ _04914_ _04907_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__a211o_1
X_14896_ _12018_ _12017_ VGND VGND VPWR VPWR _12019_ sky130_fd_sc_hd__nand2b_1
X_19423_ _06467_ _06471_ _06474_ _06475_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__o211a_1
X_16635_ _03958_ _03959_ _03942_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__a21oi_1
X_13847_ deser_A.serial_word\[8\] deser_A.shift_reg\[8\] net58 VGND VGND VPWR VPWR
+ _00673_ sky130_fd_sc_hd__mux2_1
XFILLER_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_185_Left_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19354_ _06348_ _06412_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_139_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16566_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[30\]
+ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__nand2_1
X_13778_ B_in\[85\] deser_B.word_buffer\[85\] net85 VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__mux2_1
XFILLER_210_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18305_ _05469_ _05472_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__nor2_1
XFILLER_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15517_ _12547_ _12549_ _12548_ VGND VGND VPWR VPWR _12575_ sky130_fd_sc_hd__o21bai_1
XFILLER_231_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19285_ _06310_ _06346_ systolic_inst.A_outs\[7\]\[7\] VGND VGND VPWR VPWR _06347_
+ sky130_fd_sc_hd__and3b_1
X_16497_ _03852_ _03853_ _03854_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_171_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18236_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[9\]\[7\]
+ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_171_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15448_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[3\] _12491_ _12489_
+ VGND VGND VPWR VPWR _12508_ sky130_fd_sc_hd__a31o_1
XFILLER_90_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18167_ _05327_ _05329_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_1392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15379_ systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[2\]
+ systolic_inst.B_outs\[13\]\[0\] VGND VGND VPWR VPWR _12443_ sky130_fd_sc_hd__a22oi_1
XFILLER_172_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap101 net103 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_12
XFILLER_209_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17118_ systolic_inst.acc_wires\[11\]\[20\] systolic_inst.acc_wires\[11\]\[21\] systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__o21a_1
Xmax_cap123 deser_B.serial_word_ready VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_12
XFILLER_7_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18098_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[11\] _05287_ net116
+ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__mux2_1
Xmax_cap134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_194_Left_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17049_ _04335_ _04341_ _04343_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__o21a_1
XFILLER_239_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20060_ _07039_ _07040_ _07038_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_233_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_233_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_135_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23750_ _10353_ _10355_ VGND VGND VPWR VPWR _10358_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ _07810_ _07813_ _07811_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_124_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22701_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.B_outs\[1\]\[2\] _09387_ VGND
+ VGND VPWR VPWR _09388_ sky130_fd_sc_hd__nand3_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23681_ _10250_ _10278_ _10279_ VGND VGND VPWR VPWR _10300_ sky130_fd_sc_hd__a21bo_1
XFILLER_80_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20893_ _07738_ _07769_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__xnor2_1
X_25420_ _11179_ systolic_inst.A_shift\[0\]\[1\] net71 VGND VGND VPWR VPWR _02787_
+ sky130_fd_sc_hd__mux2_1
X_22632_ _09344_ _09343_ systolic_inst.acc_wires\[2\]\[24\] net109 VGND VGND VPWR
+ VPWR _01834_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_213_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25351_ ser_C.parallel_data\[502\] net98 net78 ser_C.shift_reg\[502\] _11145_ VGND
+ VGND VPWR VPWR _02752_ sky130_fd_sc_hd__a221o_1
X_22563_ _09284_ _09285_ VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__and2_1
XFILLER_142_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_230_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_230_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24302_ _10624_ systolic_inst.A_shift\[11\]\[6\] net71 VGND VGND VPWR VPWR _02224_
+ sky130_fd_sc_hd__mux2_1
XFILLER_210_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28070_ clknet_leaf_119_clk _01868_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_21514_ _08325_ _08326_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__nand2_1
XFILLER_167_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25282_ net111 ser_C.shift_reg\[469\] VGND VGND VPWR VPWR _11111_ sky130_fd_sc_hd__and2_1
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22494_ _09220_ _09221_ _09219_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27021_ clknet_leaf_23_B_in_serial_clk _00819_ net137 VGND VGND VPWR VPWR deser_B.shift_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24233_ systolic_inst.A_shift\[19\]\[0\] A_in\[64\] net59 VGND VGND VPWR VPWR _10602_
+ sky130_fd_sc_hd__mux2_1
X_21445_ _08278_ _08281_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__xor2_1
XFILLER_182_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21376_ _08221_ _08222_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__nand2_1
X_24164_ _10583_ systolic_inst.A_shift\[27\]\[5\] net70 VGND VGND VPWR VPWR _02127_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23115_ _09774_ _09775_ _09773_ VGND VGND VPWR VPWR _09781_ sky130_fd_sc_hd__a21bo_1
X_20327_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[4\] _07263_ _07264_
+ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__a22o_1
XFILLER_134_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24095_ systolic_inst.B_shift\[23\]\[3\] B_in\[59\] net59 VGND VGND VPWR VPWR _10557_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28972_ clknet_leaf_64_clk _02770_ VGND VGND VPWR VPWR systolic_inst.A_shift\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_181_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23046_ _09691_ _09694_ _09719_ VGND VGND VPWR VPWR _09721_ sky130_fd_sc_hd__and3_1
X_27923_ clknet_leaf_145_clk _01721_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_20258_ systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[3\]
+ systolic_inst.B_outs\[5\]\[0\] VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__a22o_1
XFILLER_103_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_224_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_224_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_49_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27854_ clknet_leaf_35_clk _01652_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_20189_ _07154_ _07155_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__nand2_1
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26805_ clknet_leaf_82_clk _00607_ net153 VGND VGND VPWR VPWR B_in\[77\] sky130_fd_sc_hd__dfrtp_1
XFILLER_114_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27785_ clknet_leaf_182_clk _01583_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24997_ C_out\[325\] net97 net80 ser_C.shift_reg\[325\] _10968_ VGND VGND VPWR VPWR
+ _02575_ sky130_fd_sc_hd__a221o_1
XFILLER_85_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26736_ clknet_leaf_99_clk _00538_ net152 VGND VGND VPWR VPWR B_in\[8\] sky130_fd_sc_hd__dfrtp_1
X_29524_ clknet_leaf_260_clk _03322_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[496\]
+ sky130_fd_sc_hd__dfrtp_1
X_14750_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.B_outs\[9\]\[2\] net115 VGND
+ VGND VPWR VPWR _01020_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23948_ systolic_inst.B_shift\[14\]\[6\] B_in\[22\] net59 VGND VGND VPWR VPWR _10503_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13701_ B_in\[8\] deser_B.word_buffer\[8\] net84 VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__mux2_1
X_29455_ clknet_leaf_288_clk _03253_ net136 VGND VGND VPWR VPWR C_out\[427\] sky130_fd_sc_hd__dfrtp_1
X_26667_ clknet_leaf_6_B_in_serial_clk _00470_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14681_ _11833_ _11834_ _11835_ VGND VGND VPWR VPWR _11837_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_47_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23879_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[29\]
+ VGND VGND VPWR VPWR _10467_ sky130_fd_sc_hd__xor2_1
XFILLER_60_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16420_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[12\]\[9\]
+ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__nor2_1
XFILLER_60_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25618_ systolic_inst.acc_wires\[2\]\[30\] C_out\[94\] net50 VGND VGND VPWR VPWR
+ _02920_ sky130_fd_sc_hd__mux2_1
X_28406_ clknet_leaf_88_clk _02204_ VGND VGND VPWR VPWR systolic_inst.B_shift\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13632_ deser_B.word_buffer\[68\] deser_B.serial_word\[68\] net123 VGND VGND VPWR
+ VPWR _00469_ sky130_fd_sc_hd__mux2_1
XFILLER_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29386_ clknet_leaf_245_clk _03184_ net145 VGND VGND VPWR VPWR C_out\[358\] sky130_fd_sc_hd__dfrtp_1
X_26598_ clknet_leaf_3_B_in_serial_clk _00401_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16351_ _03729_ _03728_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__and2b_1
X_28337_ clknet_leaf_2_clk _02135_ VGND VGND VPWR VPWR systolic_inst.A_shift\[26\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_25549_ systolic_inst.acc_wires\[0\]\[25\] C_out\[25\] net53 VGND VGND VPWR VPWR
+ _02851_ sky130_fd_sc_hd__mux2_1
XFILLER_213_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13563_ deser_A.shift_reg\[127\] net2 net130 VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15302_ _12392_ VGND VGND VPWR VPWR _12393_ sky130_fd_sc_hd__inv_2
XFILLER_199_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19070_ _06117_ _06120_ _06137_ _06138_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_188_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28268_ clknet_leaf_47_clk _02066_ VGND VGND VPWR VPWR systolic_inst.B_shift\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_16282_ _03661_ _03662_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_217_Right_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13494_ deser_A.shift_reg\[58\] deser_A.shift_reg\[59\] net130 VGND VGND VPWR VPWR
+ _00331_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18021_ _05175_ _05177_ _05212_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__a21o_1
XFILLER_199_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15233_ net107 systolic_inst.acc_wires\[14\]\[12\] _12332_ _12334_ VGND VGND VPWR
+ VPWR _01054_ sky130_fd_sc_hd__a22o_1
X_27219_ clknet_leaf_291_clk _01017_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_28199_ clknet_leaf_53_clk _01997_ VGND VGND VPWR VPWR systolic_inst.B_shift\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15164_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[14\]\[3\]
+ VGND VGND VPWR VPWR _12275_ sky130_fd_sc_hd__nand2_1
XFILLER_197_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14115_ systolic_inst.B_shift\[12\]\[7\] net72 _11333_ B_in\[103\] VGND VGND VPWR
+ VPWR _00937_ sky130_fd_sc_hd__a22o_1
XFILLER_126_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19972_ _06967_ _06966_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__and2b_1
X_15095_ _12179_ _12182_ _12210_ VGND VGND VPWR VPWR _12212_ sky130_fd_sc_hd__or3_1
XFILLER_153_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14046_ deser_B.shift_reg\[80\] deser_B.shift_reg\[81\] deser_B.receiving VGND VGND
+ VPWR VPWR _00872_ sky130_fd_sc_hd__mux2_1
X_18923_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[18\]
+ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_215_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_215_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_136_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18854_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[8\]\[9\]
+ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__nor2_1
XFILLER_171_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17805_ systolic_inst.A_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[1\]
+ systolic_inst.B_outs\[9\]\[0\] VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__a22o_1
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15997_ _12983_ _12994_ _12995_ VGND VGND VPWR VPWR _12996_ sky130_fd_sc_hd__nand3_1
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18785_ _05834_ _05882_ _05881_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__o21ba_1
XFILLER_212_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17736_ _04917_ _04918_ _04940_ _04960_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__a211o_1
X_14948_ net118 _12067_ _12068_ _12069_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__a31o_1
XFILLER_82_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14879_ systolic_inst.B_outs\[14\]\[3\] systolic_inst.A_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\]
+ systolic_inst.A_outs\[14\]\[4\] VGND VGND VPWR VPWR _12002_ sky130_fd_sc_hd__and4_1
X_17667_ net60 _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__nor2_1
XFILLER_208_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19406_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[7\]\[1\]
+ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_173_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16618_ _03943_ _03942_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[3\]
+ net105 VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_196_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17598_ _11712_ _04841_ _04843_ systolic_inst.acc_wires\[10\]\[3\] net107 VGND VGND
+ VPWR VPWR _01301_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19337_ _06396_ _06397_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__or2_1
X_16549_ _03894_ _03896_ _03892_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__o21a_1
XFILLER_91_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19268_ _06274_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_132_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18219_ _05390_ _05394_ _05397_ _05398_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__o211a_1
XFILLER_176_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19199_ _06261_ _06262_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__xor2_1
XFILLER_117_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21230_ _08074_ _08096_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__or2_1
XFILLER_163_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21161_ _08028_ _08029_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_113_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20112_ _07087_ _07090_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__nand2_1
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21092_ systolic_inst.A_outs\[4\]\[4\] systolic_inst.B_outs\[4\]\[6\] VGND VGND VPWR
+ VPWR _07963_ sky130_fd_sc_hd__nand2_1
XFILLER_113_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_206_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_206_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20043_ net68 _07029_ _07031_ systolic_inst.acc_wires\[6\]\[4\] net106 VGND VGND
+ VPWR VPWR _01558_ sky130_fd_sc_hd__a32o_1
X_24920_ net110 ser_C.shift_reg\[288\] VGND VGND VPWR VPWR _10930_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_126_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24851_ C_out\[252\] net98 net78 ser_C.shift_reg\[252\] _10895_ VGND VGND VPWR VPWR
+ _02502_ sky130_fd_sc_hd__a221o_1
XFILLER_150_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23802_ _10401_ _10402_ VGND VGND VPWR VPWR _10403_ sky130_fd_sc_hd__nand2_1
XFILLER_6_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27570_ clknet_leaf_298_clk _01368_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24782_ net113 ser_C.shift_reg\[219\] VGND VGND VPWR VPWR _10861_ sky130_fd_sc_hd__and2_1
XFILLER_113_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_236_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ _08775_ _08776_ _08774_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__a21o_1
XFILLER_39_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_236_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26521_ clknet_leaf_4_A_in_serial_clk _00324_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_187_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23733_ _10340_ _10341_ _10342_ VGND VGND VPWR VPWR _10344_ sky130_fd_sc_hd__and3_1
XFILLER_148_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20945_ _07784_ _07819_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__or2_1
XFILLER_226_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_232_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29240_ clknet_leaf_176_clk _03038_ net148 VGND VGND VPWR VPWR C_out\[212\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_232_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26452_ clknet_leaf_9_clk _00259_ net132 VGND VGND VPWR VPWR A_in\[120\] sky130_fd_sc_hd__dfrtp_1
XFILLER_187_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23664_ _10154_ _10195_ _10222_ VGND VGND VPWR VPWR _10283_ sky130_fd_sc_hd__o21bai_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20876_ _07750_ _07752_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__or2_1
XFILLER_230_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25403_ systolic_inst.A_shift\[2\]\[1\] A_in\[9\] net59 VGND VGND VPWR VPWR _11171_
+ sky130_fd_sc_hd__mux2_1
X_22615_ _09328_ _09329_ _09327_ VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__o21ai_1
XFILLER_186_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29171_ clknet_leaf_43_clk _02969_ net142 VGND VGND VPWR VPWR C_out\[143\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26383_ clknet_leaf_14_clk _00190_ net133 VGND VGND VPWR VPWR A_in\[51\] sky130_fd_sc_hd__dfrtp_1
XFILLER_224_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23595_ _10216_ VGND VGND VPWR VPWR _10217_ sky130_fd_sc_hd__inv_2
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28122_ clknet_leaf_125_clk _01920_ net144 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25334_ net112 ser_C.shift_reg\[495\] VGND VGND VPWR VPWR _11137_ sky130_fd_sc_hd__and2_1
X_22546_ _09254_ _09270_ VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__nor2_1
XFILLER_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28053_ clknet_leaf_51_clk _01851_ net144 VGND VGND VPWR VPWR systolic_inst.B_outs\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_195_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25265_ ser_C.parallel_data\[459\] net102 net74 ser_C.shift_reg\[459\] _11102_ VGND
+ VGND VPWR VPWR _02709_ sky130_fd_sc_hd__a221o_1
X_22477_ net65 _09211_ _09212_ systolic_inst.acc_wires\[2\]\[1\] net109 VGND VGND
+ VPWR VPWR _01811_ sky130_fd_sc_hd__a32o_1
XFILLER_194_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27004_ clknet_leaf_15_B_in_serial_clk _00802_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_183_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24216_ _10593_ systolic_inst.A_shift\[20\]\[7\] net71 VGND VGND VPWR VPWR _02169_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21428_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[26\]
+ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__or2_1
XFILLER_135_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25196_ net111 ser_C.shift_reg\[426\] VGND VGND VPWR VPWR _11068_ sky130_fd_sc_hd__and2_1
XFILLER_205_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24147_ systolic_inst.A_shift\[29\]\[5\] A_in\[109\] net59 VGND VGND VPWR VPWR _10575_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21359_ _08204_ _08205_ _08199_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__or3b_1
XFILLER_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24078_ systolic_inst.B_shift\[3\]\[5\] _11332_ net83 systolic_inst.B_shift\[7\]\[5\]
+ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__a22o_1
X_28955_ clknet_leaf_259_clk _02753_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23029_ _09654_ _09704_ VGND VGND VPWR VPWR _09705_ sky130_fd_sc_hd__xnor2_1
X_27906_ clknet_leaf_136_clk _01704_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_15920_ _12940_ _12942_ _12944_ VGND VGND VPWR VPWR _12945_ sky130_fd_sc_hd__or3_1
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28886_ clknet_leaf_331_clk _02684_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[434\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15851_ net67 _12885_ _12886_ systolic_inst.acc_wires\[13\]\[14\] net108 VGND VGND
+ VPWR VPWR _01120_ sky130_fd_sc_hd__a32o_1
X_27837_ clknet_leaf_207_clk _01635_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_177_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _11927_ VGND VGND VPWR VPWR _11928_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_177_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15782_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[13\]\[5\]
+ VGND VGND VPWR VPWR _12827_ sky130_fd_sc_hd__or2_1
X_18570_ _05692_ _05698_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27768_ clknet_leaf_204_clk _01566_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29507_ clknet_leaf_272_clk _03305_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[479\]
+ sky130_fd_sc_hd__dfrtp_1
X_14733_ _11877_ _11880_ VGND VGND VPWR VPWR _11881_ sky130_fd_sc_hd__nand2_1
X_17521_ _04771_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__xnor2_1
X_26719_ clknet_leaf_31_B_in_serial_clk _00522_ net134 VGND VGND VPWR VPWR deser_B.word_buffer\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_27699_ clknet_leaf_197_clk _01497_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17452_ net105 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[10\] _04706_
+ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__a21bo_1
XFILLER_229_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _11802_ _11807_ _11812_ _11816_ VGND VGND VPWR VPWR _11822_ sky130_fd_sc_hd__or4_1
X_29438_ clknet_leaf_332_clk _03236_ net131 VGND VGND VPWR VPWR C_out\[410\] sky130_fd_sc_hd__dfrtp_1
XFILLER_232_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16403_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[12\]\[6\]
+ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__nand2_1
X_13615_ deser_B.word_buffer\[51\] deser_B.serial_word\[51\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__mux2_1
X_17383_ _04608_ _04610_ _04607_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__o21ba_1
XFILLER_242_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29369_ clknet_leaf_232_clk _03167_ net147 VGND VGND VPWR VPWR C_out\[341\] sky130_fd_sc_hd__dfrtp_1
X_14595_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[15\]\[9\]
+ _11758_ VGND VGND VPWR VPWR _11763_ sky130_fd_sc_hd__a21oi_1
XFILLER_198_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19122_ _06186_ _06187_ _06175_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__o21bai_1
X_16334_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[13\] _03713_ net115
+ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__mux2_1
X_13546_ deser_A.shift_reg\[110\] deser_A.shift_reg\[111\] net129 VGND VGND VPWR VPWR
+ _00383_ sky130_fd_sc_hd__mux2_1
XFILLER_201_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19053_ _06108_ _06110_ _06121_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__a21oi_1
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16265_ _03592_ _03610_ _03609_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__o21a_1
X_13477_ deser_A.shift_reg\[41\] deser_A.shift_reg\[42\] net130 VGND VGND VPWR VPWR
+ _00314_ sky130_fd_sc_hd__mux2_1
X_15216_ net107 systolic_inst.acc_wires\[14\]\[10\] _11712_ _12319_ VGND VGND VPWR
+ VPWR _01052_ sky130_fd_sc_hd__a22o_1
X_18004_ systolic_inst.A_outs\[9\]\[4\] systolic_inst.B_outs\[9\]\[5\] VGND VGND VPWR
+ VPWR _05196_ sky130_fd_sc_hd__nand2_1
XFILLER_173_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16196_ _03577_ _03578_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15147_ net118 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[14\]\[0\]
+ VGND VGND VPWR VPWR _12261_ sky130_fd_sc_hd__a21oi_1
XFILLER_236_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19955_ systolic_inst.B_outs\[6\]\[6\] systolic_inst.A_outs\[6\]\[7\] VGND VGND VPWR
+ VPWR _06951_ sky130_fd_sc_hd__nand2_1
X_15078_ _12141_ _12195_ VGND VGND VPWR VPWR _12196_ sky130_fd_sc_hd__and2b_1
XFILLER_141_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14029_ deser_B.shift_reg\[63\] deser_B.shift_reg\[64\] net126 VGND VGND VPWR VPWR
+ _00855_ sky130_fd_sc_hd__mux2_1
XFILLER_141_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18906_ _06007_ _06008_ _06002_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__or3b_1
X_19886_ _06816_ _06847_ _06848_ _06815_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__nor4b_1
XFILLER_68_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18837_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[8\]\[6\]
+ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__nand2_1
XFILLER_3_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18768_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[13\] _05891_
+ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__a21o_1
XFILLER_236_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17719_ _04938_ _04944_ _04945_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18699_ _05787_ _05789_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__nand3_1
XFILLER_224_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20730_ _07641_ _07642_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__nand2_1
XFILLER_24_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20661_ _07580_ _07581_ _07582_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__and3_1
XFILLER_149_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22400_ _09093_ _09109_ _09107_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_119_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20592_ systolic_inst.A_outs\[5\]\[6\] _11276_ _07494_ _07497_ _07522_ VGND VGND
+ VPWR VPWR _07523_ sky130_fd_sc_hd__o311a_1
X_23380_ _10005_ _10006_ VGND VGND VPWR VPWR _10007_ sky130_fd_sc_hd__and2_1
XFILLER_31_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22331_ _09029_ _09037_ _09036_ VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__a21bo_1
XFILLER_178_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25050_ net112 ser_C.shift_reg\[353\] VGND VGND VPWR VPWR _10995_ sky130_fd_sc_hd__and2_1
X_22262_ _08989_ _09006_ VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24001_ systolic_inst.B_shift\[9\]\[4\] B_in\[12\] _00008_ VGND VGND VPWR VPWR _10526_
+ sky130_fd_sc_hd__mux2_1
XFILLER_145_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21213_ _08028_ _08080_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_225_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22193_ _08937_ _08938_ _08915_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21144_ _08011_ _08012_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_221_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25952_ systolic_inst.acc_wires\[13\]\[12\] C_out\[428\] net19 VGND VGND VPWR VPWR
+ _03254_ sky130_fd_sc_hd__mux2_1
XFILLER_59_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28740_ clknet_leaf_296_clk _02538_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[288\]
+ sky130_fd_sc_hd__dfrtp_1
X_21075_ _07903_ _07905_ _07945_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__and3_1
XFILLER_24_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_238_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20026_ _07014_ _07015_ _07016_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_31_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24903_ C_out\[278\] net103 net75 ser_C.shift_reg\[278\] _10921_ VGND VGND VPWR VPWR
+ _02528_ sky130_fd_sc_hd__a221o_1
X_28671_ clknet_leaf_185_clk _02469_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[219\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25883_ systolic_inst.acc_wires\[11\]\[7\] C_out\[359\] net39 VGND VGND VPWR VPWR
+ _03185_ sky130_fd_sc_hd__mux2_1
XFILLER_219_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24834_ net113 ser_C.shift_reg\[245\] VGND VGND VPWR VPWR _10887_ sky130_fd_sc_hd__and2_1
X_27622_ clknet_leaf_317_clk _01420_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_206_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27553_ clknet_leaf_298_clk _01351_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24765_ C_out\[209\] net99 net79 ser_C.shift_reg\[209\] _10852_ VGND VGND VPWR VPWR
+ _02459_ sky130_fd_sc_hd__a221o_1
XFILLER_61_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21977_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[15\]
+ _08757_ _08760_ _08761_ VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__a221oi_2
XFILLER_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26504_ clknet_leaf_16_A_in_serial_clk _00307_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_23716_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[0\]\[4\]
+ VGND VGND VPWR VPWR _10329_ sky130_fd_sc_hd__or2_1
XFILLER_226_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27484_ clknet_leaf_296_clk _01282_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_20928_ systolic_inst.A_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\]
+ systolic_inst.A_outs\[4\]\[2\] VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__a22oi_1
XFILLER_109_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24696_ net112 ser_C.shift_reg\[176\] VGND VGND VPWR VPWR _10818_ sky130_fd_sc_hd__and2_1
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29223_ clknet_leaf_211_clk _03021_ net147 VGND VGND VPWR VPWR C_out\[195\] sky130_fd_sc_hd__dfrtp_1
X_26435_ clknet_leaf_1_clk _00242_ net131 VGND VGND VPWR VPWR A_in\[103\] sky130_fd_sc_hd__dfrtp_1
XFILLER_202_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23647_ _10256_ _10265_ VGND VGND VPWR VPWR _10267_ sky130_fd_sc_hd__xnor2_1
XFILLER_230_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20859_ systolic_inst.A_outs\[4\]\[0\] systolic_inst.B_outs\[4\]\[3\] _07729_ VGND
+ VGND VPWR VPWR _07737_ sky130_fd_sc_hd__a21o_1
XFILLER_35_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13400_ A_in\[109\] deser_A.word_buffer\[109\] net96 VGND VGND VPWR VPWR _00248_
+ sky130_fd_sc_hd__mux2_1
X_29154_ clknet_leaf_169_clk _02952_ net148 VGND VGND VPWR VPWR C_out\[126\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14380_ _11562_ _11563_ VGND VGND VPWR VPWR _11564_ sky130_fd_sc_hd__nor2_1
X_26366_ clknet_leaf_25_clk _00173_ net137 VGND VGND VPWR VPWR A_in\[34\] sky130_fd_sc_hd__dfrtp_1
X_23578_ _10119_ _10159_ _10080_ VGND VGND VPWR VPWR _10200_ sky130_fd_sc_hd__o21bai_1
XFILLER_126_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28105_ clknet_leaf_156_clk _01903_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25317_ ser_C.parallel_data\[485\] net97 net77 ser_C.shift_reg\[485\] _11128_ VGND
+ VGND VPWR VPWR _02735_ sky130_fd_sc_hd__a221o_1
X_13331_ A_in\[40\] deser_A.word_buffer\[40\] net93 VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__mux2_1
X_29085_ clknet_leaf_111_clk _02883_ net151 VGND VGND VPWR VPWR C_out\[57\] sky130_fd_sc_hd__dfrtp_1
X_22529_ net60 _09256_ VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__nor2_1
X_26297_ clknet_leaf_25_A_in_serial_clk _00105_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_210_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28036_ clknet_leaf_159_clk _01834_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_202_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16050_ _13016_ _13046_ VGND VGND VPWR VPWR _13047_ sky130_fd_sc_hd__nand2_1
X_25248_ net111 ser_C.shift_reg\[452\] VGND VGND VPWR VPWR _11094_ sky130_fd_sc_hd__and2_1
X_13262_ deser_A.word_buffer\[100\] deser_A.serial_word\[100\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__mux2_1
XFILLER_108_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15001_ _12111_ _12119_ VGND VGND VPWR VPWR _12121_ sky130_fd_sc_hd__or2_1
XFILLER_237_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25179_ C_out\[416\] net103 net75 ser_C.shift_reg\[416\] _11059_ VGND VGND VPWR VPWR
+ _02666_ sky130_fd_sc_hd__a221o_1
X_13193_ deser_A.word_buffer\[31\] deser_A.serial_word\[31\] net128 VGND VGND VPWR
+ VPWR _00041_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19740_ _06712_ _06715_ _06717_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_8_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28938_ clknet_leaf_259_clk _02736_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[486\]
+ sky130_fd_sc_hd__dfrtp_1
X_16952_ _04265_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__nor2_1
XFILLER_238_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15903_ net67 _12929_ _12930_ systolic_inst.acc_wires\[13\]\[22\] net108 VGND VGND
+ VPWR VPWR _01128_ sky130_fd_sc_hd__a32o_1
X_19671_ _06668_ _06674_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__and2_1
XFILLER_38_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28869_ clknet_leaf_300_clk _02667_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[417\]
+ sky130_fd_sc_hd__dfrtp_1
X_16883_ _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__inv_2
XFILLER_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18622_ _05748_ _05749_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__and2b_1
XFILLER_237_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15834_ _12870_ _12871_ VGND VGND VPWR VPWR _12872_ sky130_fd_sc_hd__nor2_1
XFILLER_46_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18553_ _05682_ _05681_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__nand2b_1
X_15765_ _12812_ VGND VGND VPWR VPWR _12813_ sky130_fd_sc_hd__inv_2
XFILLER_205_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17504_ _04711_ _04727_ _04725_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__o21a_1
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14716_ _11850_ _11852_ _11864_ _11865_ _11858_ VGND VGND VPWR VPWR _11866_ sky130_fd_sc_hd__a311oi_4
X_15696_ _12720_ _12748_ VGND VGND VPWR VPWR _12749_ sky130_fd_sc_hd__nand2b_1
X_18484_ _05606_ _05614_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_159_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14647_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[16\]
+ _11804_ VGND VGND VPWR VPWR _11808_ sky130_fd_sc_hd__a21oi_1
X_17435_ _04647_ _04655_ _04654_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_155_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ _11745_ _11746_ _11747_ VGND VGND VPWR VPWR _11749_ sky130_fd_sc_hd__nand3_1
XANTENNA_29 net142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17366_ _04621_ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19105_ _06170_ _06171_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__or2_1
XFILLER_14_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16317_ _03632_ _03696_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__nand2_1
X_13529_ deser_A.shift_reg\[93\] deser_A.shift_reg\[94\] net129 VGND VGND VPWR VPWR
+ _00366_ sky130_fd_sc_hd__mux2_1
XFILLER_186_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17297_ _04523_ _04525_ _04554_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_168_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19036_ _06105_ _06106_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__or2_1
X_16248_ systolic_inst.B_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\] VGND VGND
+ VPWR VPWR _03630_ sky130_fd_sc_hd__or2_1
XFILLER_51_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16179_ _03561_ _03562_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_110_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19938_ _06902_ _06904_ _06933_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__nand3_1
XFILLER_60_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19869_ _06865_ _06866_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_108_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21900_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[3\]\[5\]
+ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22880_ _09558_ _09559_ VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__nor2_1
XFILLER_3_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21831_ _08602_ _08604_ _08634_ VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_69_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24550_ net113 ser_C.shift_reg\[103\] VGND VGND VPWR VPWR _10745_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21762_ _08528_ _08530_ _08566_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__nand3_1
XFILLER_169_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23501_ _10123_ _10124_ VGND VGND VPWR VPWR _10125_ sky130_fd_sc_hd__or2_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20713_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[5\]\[14\]
+ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__nand2_1
X_24481_ C_out\[67\] _11302_ net81 ser_C.shift_reg\[67\] _10710_ VGND VGND VPWR VPWR
+ _02317_ sky130_fd_sc_hd__a221o_1
XFILLER_211_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21693_ _08499_ _08500_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__nand2_1
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26220_ clknet_leaf_8_A_in_serial_clk _00028_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23432_ _10015_ _10017_ _10056_ _10057_ VGND VGND VPWR VPWR _10058_ sky130_fd_sc_hd__a211oi_1
XFILLER_71_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20644_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[5\]\[4\]
+ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26151_ deser_B.serial_word\[106\] deser_B.shift_reg\[106\] _00001_ VGND VGND VPWR
+ VPWR _03453_ sky130_fd_sc_hd__mux2_1
XFILLER_32_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23363_ systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[6\]
+ systolic_inst.B_outs\[0\]\[0\] VGND VGND VPWR VPWR _09990_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_227_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20575_ _07504_ _07505_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__xor2_1
XFILLER_20_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_227_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25102_ net113 ser_C.shift_reg\[379\] VGND VGND VPWR VPWR _11021_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22314_ _08985_ _09055_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__and2_1
XFILLER_165_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26082_ deser_B.serial_word\[37\] deser_B.shift_reg\[37\] net55 VGND VGND VPWR VPWR
+ _03384_ sky130_fd_sc_hd__mux2_1
X_23294_ _09924_ VGND VGND VPWR VPWR _09925_ sky130_fd_sc_hd__inv_2
XFILLER_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25033_ C_out\[343\] net97 net77 ser_C.shift_reg\[343\] _10986_ VGND VGND VPWR VPWR
+ _02593_ sky130_fd_sc_hd__a221o_1
X_22245_ systolic_inst.B_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\] systolic_inst.A_outs\[2\]\[4\]
+ systolic_inst.A_outs\[2\]\[5\] VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__and4_1
XFILLER_156_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22176_ systolic_inst.A_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[3\] systolic_inst.A_outs\[2\]\[3\]
+ systolic_inst.B_outs\[2\]\[4\] VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__nand4_2
XFILLER_133_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21127_ _07995_ _07996_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__nand2_1
XFILLER_120_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26984_ clknet_leaf_0_A_in_serial_clk _00782_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28723_ clknet_leaf_312_clk _02521_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[271\]
+ sky130_fd_sc_hd__dfrtp_1
X_21058_ systolic_inst.A_outs\[4\]\[2\] _07852_ _07928_ VGND VGND VPWR VPWR _07930_
+ sky130_fd_sc_hd__o21a_1
XFILLER_28_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25935_ systolic_inst.acc_wires\[12\]\[27\] C_out\[411\] net21 VGND VGND VPWR VPWR
+ _03237_ sky130_fd_sc_hd__mux2_1
XFILLER_87_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_203_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20009_ _07001_ _07002_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__xnor2_1
X_28654_ clknet_leaf_203_clk _02452_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[202\]
+ sky130_fd_sc_hd__dfrtp_1
X_13880_ deser_A.serial_word\[41\] deser_A.shift_reg\[41\] net58 VGND VGND VPWR VPWR
+ _00706_ sky130_fd_sc_hd__mux2_1
X_25866_ systolic_inst.acc_wires\[10\]\[22\] C_out\[342\] net11 VGND VGND VPWR VPWR
+ _03168_ sky130_fd_sc_hd__mux2_1
XFILLER_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27605_ clknet_leaf_203_clk _01403_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_24817_ C_out\[235\] net99 net79 ser_C.shift_reg\[235\] _10878_ VGND VGND VPWR VPWR
+ _02485_ sky130_fd_sc_hd__a221o_1
XFILLER_41_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25797_ systolic_inst.acc_wires\[8\]\[17\] C_out\[273\] net28 VGND VGND VPWR VPWR
+ _03099_ sky130_fd_sc_hd__mux2_1
X_28585_ clknet_leaf_309_clk _02383_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15550_ _12607_ _12606_ VGND VGND VPWR VPWR _12608_ sky130_fd_sc_hd__and2b_1
X_24748_ net112 ser_C.shift_reg\[202\] VGND VGND VPWR VPWR _10844_ sky130_fd_sc_hd__and2_1
XFILLER_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27536_ clknet_leaf_310_clk _01334_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_43_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14501_ _11593_ _11679_ VGND VGND VPWR VPWR _11681_ sky130_fd_sc_hd__nand2_1
XFILLER_188_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27467_ clknet_leaf_236_clk _01265_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_15481_ systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[6\] systolic_inst.A_outs\[13\]\[7\]
+ systolic_inst.B_outs\[13\]\[0\] VGND VGND VPWR VPWR _12540_ sky130_fd_sc_hd__a22o_1
XFILLER_203_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24679_ C_out\[166\] net103 net76 ser_C.shift_reg\[166\] _10809_ VGND VGND VPWR VPWR
+ _02416_ sky130_fd_sc_hd__a221o_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29206_ clknet_leaf_204_clk _03004_ net146 VGND VGND VPWR VPWR C_out\[178\] sky130_fd_sc_hd__dfrtp_1
X_14432_ _11614_ VGND VGND VPWR VPWR _11615_ sky130_fd_sc_hd__inv_2
X_17220_ _04473_ _04475_ _04479_ _04480_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__o22a_1
X_26418_ clknet_leaf_7_clk _00225_ net134 VGND VGND VPWR VPWR A_in\[86\] sky130_fd_sc_hd__dfrtp_1
X_27398_ clknet_leaf_332_clk _01196_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17151_ _04435_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__xnor2_1
X_29137_ clknet_leaf_168_clk _02935_ net148 VGND VGND VPWR VPWR C_out\[109\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26349_ clknet_leaf_63_clk _00156_ net135 VGND VGND VPWR VPWR A_in\[17\] sky130_fd_sc_hd__dfrtp_1
X_14363_ _11503_ _11505_ _11545_ VGND VGND VPWR VPWR _11548_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_150_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16102_ systolic_inst.A_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[4\]
+ systolic_inst.B_outs\[12\]\[3\] VGND VGND VPWR VPWR _13097_ sky130_fd_sc_hd__a22oi_1
XFILLER_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13314_ A_in\[23\] deser_A.word_buffer\[23\] net91 VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__mux2_1
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29068_ clknet_leaf_116_clk _02866_ net152 VGND VGND VPWR VPWR C_out\[40\] sky130_fd_sc_hd__dfrtp_1
XFILLER_116_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17082_ _04376_ _04377_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__nor2_1
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14294_ _11477_ _11479_ VGND VGND VPWR VPWR _11480_ sky130_fd_sc_hd__nand2_1
XFILLER_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16033_ _13028_ _13029_ VGND VGND VPWR VPWR _13030_ sky130_fd_sc_hd__or2_1
X_28019_ clknet_leaf_154_clk _01817_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13245_ deser_A.word_buffer\[83\] deser_A.serial_word\[83\] net127 VGND VGND VPWR
+ VPWR _00093_ sky130_fd_sc_hd__mux2_1
XFILLER_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13176_ deser_A.word_buffer\[14\] deser_A.serial_word\[14\] net127 VGND VGND VPWR
+ VPWR _00024_ sky130_fd_sc_hd__mux2_1
XFILLER_97_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17984_ _05176_ _05146_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__nand2b_1
XFILLER_96_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19723_ systolic_inst.A_outs\[6\]\[1\] systolic_inst.B_outs\[6\]\[6\] VGND VGND VPWR
+ VPWR _06726_ sky130_fd_sc_hd__nand2_1
XFILLER_172_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16935_ _04224_ _04225_ _04221_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__a21bo_1
XFILLER_238_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19654_ _06638_ _06645_ _06647_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__a21bo_1
XFILLER_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16866_ _04130_ _04147_ _04145_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_0_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18605_ _05695_ _05731_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__and2_1
XFILLER_203_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15817_ _12850_ _12856_ VGND VGND VPWR VPWR _12857_ sky130_fd_sc_hd__nand2_1
X_19585_ _06613_ _06614_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_103_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16797_ _04061_ _04078_ _04077_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__o21ba_1
XFILLER_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18536_ systolic_inst.B_outs\[8\]\[3\] systolic_inst.A_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\]
+ systolic_inst.A_outs\[8\]\[4\] VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__and4_1
XFILLER_94_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15748_ net115 _12788_ _12798_ VGND VGND VPWR VPWR _12799_ sky130_fd_sc_hd__and3_1
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18467_ net108 _05598_ _05599_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__or3_1
XFILLER_179_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15679_ _12730_ _12731_ VGND VGND VPWR VPWR _12733_ sky130_fd_sc_hd__and2b_1
XFILLER_209_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17418_ _04602_ _04671_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18398_ net66 _05551_ _05552_ systolic_inst.acc_wires\[9\]\[30\] net105 VGND VGND
+ VPWR VPWR _01392_ sky130_fd_sc_hd__a32o_1
XFILLER_140_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17349_ _04599_ _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload210 clknet_leaf_43_clk VGND VGND VPWR VPWR clkload210/Y sky130_fd_sc_hd__bufinv_16
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20360_ systolic_inst.A_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\] systolic_inst.B_outs\[5\]\[5\]
+ systolic_inst.A_outs\[5\]\[2\] VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__a22o_1
Xclkload221 clknet_leaf_56_clk VGND VGND VPWR VPWR clkload221/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_105_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload232 clknet_leaf_83_clk VGND VGND VPWR VPWR clkload232/Y sky130_fd_sc_hd__clkinv_2
XFILLER_228_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload243 clknet_leaf_96_clk VGND VGND VPWR VPWR clkload243/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload254 clknet_leaf_93_clk VGND VGND VPWR VPWR clkload254/Y sky130_fd_sc_hd__bufinv_16
X_19019_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[2\]\[0\] net119 VGND
+ VGND VPWR VPWR _01466_ sky130_fd_sc_hd__mux2_1
X_20291_ _07229_ _07230_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__nor2_1
Xclkload265 clknet_leaf_40_clk VGND VGND VPWR VPWR clkload265/X sky130_fd_sc_hd__clkbuf_4
Xclkload276 clknet_leaf_144_clk VGND VGND VPWR VPWR clkload276/Y sky130_fd_sc_hd__clkinv_4
Xclkload287 clknet_leaf_191_clk VGND VGND VPWR VPWR clkload287/Y sky130_fd_sc_hd__clkinv_8
X_22030_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[24\]
+ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__and2_1
Xclkload298 clknet_leaf_178_clk VGND VGND VPWR VPWR clkload298/Y sky130_fd_sc_hd__clkinv_8
XFILLER_216_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23981_ systolic_inst.B_shift\[12\]\[2\] B_in\[66\] _00008_ VGND VGND VPWR VPWR _10516_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25720_ systolic_inst.acc_wires\[6\]\[4\] C_out\[196\] net47 VGND VGND VPWR VPWR
+ _03022_ sky130_fd_sc_hd__mux2_1
XFILLER_116_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22932_ _09554_ _09610_ VGND VGND VPWR VPWR _09611_ sky130_fd_sc_hd__nand2_1
XFILLER_228_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25651_ systolic_inst.acc_wires\[3\]\[31\] C_out\[127\] net49 VGND VGND VPWR VPWR
+ _02953_ sky130_fd_sc_hd__mux2_1
XFILLER_228_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22863_ _09512_ _09542_ VGND VGND VPWR VPWR _09544_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_216_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_216_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24602_ net110 ser_C.shift_reg\[129\] VGND VGND VPWR VPWR _10771_ sky130_fd_sc_hd__and2_1
X_21814_ _08590_ _08617_ VGND VGND VPWR VPWR _08618_ sky130_fd_sc_hd__nand2b_1
X_28370_ clknet_leaf_4_clk _02168_ VGND VGND VPWR VPWR systolic_inst.A_shift\[20\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xwire51 net52 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_8
X_25582_ systolic_inst.acc_wires\[1\]\[26\] C_out\[58\] net52 VGND VGND VPWR VPWR
+ _02884_ sky130_fd_sc_hd__mux2_1
X_22794_ _09446_ _09476_ VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__xnor2_1
XFILLER_227_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27321_ clknet_leaf_329_clk _01119_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_24533_ C_out\[93\] net100 net82 ser_C.shift_reg\[93\] _10736_ VGND VGND VPWR VPWR
+ _02343_ sky130_fd_sc_hd__a221o_1
XFILLER_52_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21745_ _08443_ _08550_ VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__or2_1
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27252_ clknet_leaf_271_clk _01050_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24464_ net114 ser_C.shift_reg\[60\] VGND VGND VPWR VPWR _10702_ sky130_fd_sc_hd__and2_1
XFILLER_185_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21676_ _08482_ _08483_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__or2_1
XFILLER_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26203_ clknet_leaf_14_A_in_serial_clk _00011_ net143 VGND VGND VPWR VPWR deser_A.word_buffer\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_1253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23415_ systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[5\] systolic_inst.A_outs\[0\]\[6\]
+ systolic_inst.B_outs\[0\]\[1\] VGND VGND VPWR VPWR _10041_ sky130_fd_sc_hd__a22oi_1
X_20627_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[5\]\[0\]
+ _07551_ _07552_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__a22o_1
X_27183_ clknet_leaf_264_clk _00981_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24395_ C_out\[24\] net104 _10643_ ser_C.shift_reg\[24\] _10667_ VGND VGND VPWR VPWR
+ _02274_ sky130_fd_sc_hd__a221o_1
XFILLER_137_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26134_ deser_B.serial_word\[89\] deser_B.shift_reg\[89\] net56 VGND VGND VPWR VPWR
+ _03436_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23346_ systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[3\] systolic_inst.A_outs\[0\]\[4\]
+ systolic_inst.B_outs\[0\]\[1\] VGND VGND VPWR VPWR _09974_ sky130_fd_sc_hd__a22oi_1
XFILLER_138_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20558_ _07422_ _07427_ _07457_ _07489_ _07456_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__a311oi_2
XFILLER_138_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_89_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26065_ deser_B.serial_word\[20\] deser_B.shift_reg\[20\] net55 VGND VGND VPWR VPWR
+ _03367_ sky130_fd_sc_hd__mux2_1
XFILLER_152_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23277_ systolic_inst.A_outs\[0\]\[0\] systolic_inst.A_shift\[0\]\[0\] net121 VGND
+ VGND VPWR VPWR _01906_ sky130_fd_sc_hd__mux2_1
XFILLER_180_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20489_ _07422_ _07423_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__nand2_1
X_25016_ net111 ser_C.shift_reg\[336\] VGND VGND VPWR VPWR _10978_ sky130_fd_sc_hd__and2_1
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22228_ _08971_ _08972_ VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_205_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22159_ _08897_ _08905_ VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__xor2_1
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_205_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14981_ _12061_ _12067_ _12101_ VGND VGND VPWR VPWR _12102_ sky130_fd_sc_hd__a21oi_1
X_26967_ clknet_leaf_24_A_in_serial_clk _00765_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28706_ clknet_leaf_184_clk _02504_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[254\]
+ sky130_fd_sc_hd__dfrtp_1
X_16720_ _04003_ _04039_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_197_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25918_ systolic_inst.acc_wires\[12\]\[10\] C_out\[394\] net18 VGND VGND VPWR VPWR
+ _03220_ sky130_fd_sc_hd__mux2_1
X_13932_ deser_A.serial_word\[93\] deser_A.shift_reg\[93\] net57 VGND VGND VPWR VPWR
+ _00758_ sky130_fd_sc_hd__mux2_1
X_29686_ clknet_leaf_105_clk _03481_ net152 VGND VGND VPWR VPWR ser_C.bit_idx\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26898_ clknet_leaf_10_A_in_serial_clk _00696_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28637_ clknet_leaf_182_clk _02435_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[185\]
+ sky130_fd_sc_hd__dfrtp_1
X_13863_ deser_A.serial_word\[24\] deser_A.shift_reg\[24\] net58 VGND VGND VPWR VPWR
+ _00689_ sky130_fd_sc_hd__mux2_1
XFILLER_78_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16651_ _03973_ _03974_ systolic_inst.A_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[5\]
+ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_193_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25849_ systolic_inst.acc_wires\[10\]\[5\] C_out\[325\] net12 VGND VGND VPWR VPWR
+ _03151_ sky130_fd_sc_hd__mux2_1
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15602_ _12655_ _12656_ VGND VGND VPWR VPWR _12658_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19370_ net105 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[13\] _06428_
+ _06429_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__a22o_1
X_28568_ clknet_leaf_165_clk _02366_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_13794_ B_in\[101\] deser_B.word_buffer\[101\] _00005_ VGND VGND VPWR VPWR _00631_
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16582_ systolic_inst.A_outs\[11\]\[7\] systolic_inst.A_outs\[10\]\[7\] net118 VGND
+ VGND VPWR VPWR _01209_ sky130_fd_sc_hd__mux2_1
XFILLER_234_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18321_ _05480_ _05484_ _05486_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_5_21__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_21__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_27519_ clknet_leaf_232_clk _01317_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15533_ _12587_ _12590_ VGND VGND VPWR VPWR _12591_ sky130_fd_sc_hd__xnor2_1
X_28499_ clknet_leaf_112_clk _02297_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15464_ _12517_ _12518_ _12522_ VGND VGND VPWR VPWR _12524_ sky130_fd_sc_hd__a21o_1
X_18252_ _05419_ _05422_ _05425_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__a21bo_1
XFILLER_188_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14415_ _11594_ _11597_ VGND VGND VPWR VPWR _11598_ sky130_fd_sc_hd__xor2_1
X_17203_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[1\]
+ systolic_inst.A_outs\[10\]\[2\] VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__and4_1
X_15395_ _12452_ _12457_ VGND VGND VPWR VPWR _12458_ sky130_fd_sc_hd__nand2_1
X_18183_ net116 _05368_ _05369_ _05346_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__a31o_1
XFILLER_156_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17134_ _04421_ _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__or2_1
XFILLER_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14346_ systolic_inst.A_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[6\] _11529_ VGND
+ VGND VPWR VPWR _11531_ sky130_fd_sc_hd__and3_1
XFILLER_156_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17065_ _04361_ _04362_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__nand2_1
XFILLER_170_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14277_ _11446_ _11463_ VGND VGND VPWR VPWR _11464_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16016_ _12994_ _13013_ VGND VGND VPWR VPWR _13014_ sky130_fd_sc_hd__nor2_1
XFILLER_48_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13228_ deser_A.word_buffer\[66\] deser_A.serial_word\[66\] net127 VGND VGND VPWR
+ VPWR _00076_ sky130_fd_sc_hd__mux2_1
XFILLER_174_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13159_ B_in_valid A_in_valid net6 systolic_inst.ce_local VGND VGND VPWR VPWR _11306_
+ sky130_fd_sc_hd__a31o_4
XFILLER_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17967_ systolic_inst.A_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[5\] VGND VGND VPWR
+ VPWR _05160_ sky130_fd_sc_hd__nand2_1
X_19706_ _06708_ _06709_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16918_ _04233_ _04232_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__nand2b_1
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17898_ systolic_inst.A_outs\[9\]\[1\] systolic_inst.B_outs\[9\]\[6\] VGND VGND VPWR
+ VPWR _05093_ sky130_fd_sc_hd__nand2_1
X_19637_ _06641_ _06642_ _06643_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__a21o_1
X_16849_ systolic_inst.B_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\] VGND VGND
+ VPWR VPWR _04167_ sky130_fd_sc_hd__or2_1
XFILLER_26_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19568_ _06599_ _06600_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18519_ _05647_ _05648_ _05625_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19499_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[7\]\[13\]
+ _06537_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21530_ net106 _08341_ _08342_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__or3_1
XFILLER_209_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21461_ _08289_ _08293_ _08294_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__a21oi_1
XFILLER_222_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23200_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[20\]
+ VGND VGND VPWR VPWR _09853_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20412_ _07346_ _07347_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__xnor2_1
X_24180_ systolic_inst.A_shift\[25\]\[3\] net70 _10505_ systolic_inst.A_shift\[26\]\[3\]
+ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__a22o_1
XFILLER_105_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21392_ systolic_inst.acc_wires\[4\]\[16\] systolic_inst.acc_wires\[4\]\[17\] systolic_inst.acc_wires\[4\]\[18\]
+ systolic_inst.acc_wires\[4\]\[19\] systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_96_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23131_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[1\]\[10\]
+ VGND VGND VPWR VPWR _09794_ sky130_fd_sc_hd__nand2_1
XFILLER_134_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20343_ _07279_ _07280_ _07246_ _07248_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__a211o_1
XFILLER_162_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23062_ _09656_ _09722_ _09720_ VGND VGND VPWR VPWR _09736_ sky130_fd_sc_hd__a21oi_1
X_20274_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[3\]
+ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_241_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22013_ _08783_ _08789_ _08790_ net60 VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__a31o_1
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_241_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27870_ clknet_leaf_310_clk _01668_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_192_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26821_ clknet_leaf_70_clk _00623_ net135 VGND VGND VPWR VPWR B_in\[93\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29540_ clknet_leaf_34_clk net59 net136 VGND VGND VPWR VPWR systolic_inst.load_acc
+ sky130_fd_sc_hd__dfrtp_4
X_23964_ _10507_ systolic_inst.B_shift\[9\]\[1\] net72 VGND VGND VPWR VPWR _02003_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26752_ clknet_leaf_57_clk _00554_ net137 VGND VGND VPWR VPWR B_in\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_99_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22915_ systolic_inst.A_outs\[1\]\[3\] systolic_inst.A_outs\[1\]\[4\] systolic_inst.B_outs\[1\]\[6\]
+ systolic_inst.B_outs\[1\]\[7\] VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__and4b_1
X_25703_ systolic_inst.acc_wires\[5\]\[19\] C_out\[179\] net45 VGND VGND VPWR VPWR
+ _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_216_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26683_ clknet_leaf_24_B_in_serial_clk _00486_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[85\]
+ sky130_fd_sc_hd__dfrtp_1
X_29471_ clknet_leaf_285_clk _03269_ net136 VGND VGND VPWR VPWR ser_C.parallel_data\[443\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23895_ _10480_ _10479_ systolic_inst.acc_wires\[0\]\[31\] _11258_ VGND VGND VPWR
+ VPWR _01961_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28422_ clknet_leaf_23_clk _02220_ VGND VGND VPWR VPWR systolic_inst.A_shift\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25634_ systolic_inst.acc_wires\[3\]\[14\] C_out\[110\] net51 VGND VGND VPWR VPWR
+ _02936_ sky130_fd_sc_hd__mux2_1
X_22846_ systolic_inst.A_outs\[1\]\[2\] systolic_inst.B_outs\[1\]\[6\] VGND VGND VPWR
+ VPWR _09527_ sky130_fd_sc_hd__nand2_1
XFILLER_204_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25565_ systolic_inst.acc_wires\[1\]\[9\] C_out\[41\] net36 VGND VGND VPWR VPWR _02867_
+ sky130_fd_sc_hd__mux2_1
X_28353_ clknet_leaf_343_clk _02151_ VGND VGND VPWR VPWR systolic_inst.A_shift\[24\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22777_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[4\] _09457_ _09458_
+ VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__a22o_1
XFILLER_73_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24516_ net114 ser_C.shift_reg\[86\] VGND VGND VPWR VPWR _10728_ sky130_fd_sc_hd__and2_1
XFILLER_227_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27304_ clknet_leaf_288_clk _01102_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_197_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21728_ _08532_ _08533_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_45_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25496_ _11225_ _11227_ systolic_inst.cycle_cnt\[21\] VGND VGND VPWR VPWR _02815_
+ sky130_fd_sc_hd__mux2_1
X_28284_ clknet_leaf_61_clk _02082_ VGND VGND VPWR VPWR systolic_inst.B_shift\[19\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24447_ C_out\[50\] _11302_ net81 ser_C.shift_reg\[50\] _10693_ VGND VGND VPWR VPWR
+ _02300_ sky130_fd_sc_hd__a221o_1
X_27235_ clknet_leaf_275_clk _01033_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_21659_ _08467_ _08466_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__nand2b_1
XFILLER_240_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14200_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\]
+ systolic_inst.A_outs\[15\]\[1\] VGND VGND VPWR VPWR _11389_ sky130_fd_sc_hd__a22oi_2
XFILLER_201_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27166_ clknet_leaf_273_clk _00964_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_15180_ _12287_ _12288_ _12280_ _12284_ VGND VGND VPWR VPWR _12289_ sky130_fd_sc_hd__a211o_1
X_24378_ net7 ser_C.shift_reg\[17\] VGND VGND VPWR VPWR _10659_ sky130_fd_sc_hd__and2_1
XFILLER_240_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26117_ deser_B.serial_word\[72\] deser_B.shift_reg\[72\] _00001_ VGND VGND VPWR
+ VPWR _03419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14131_ systolic_inst.A_outs\[15\]\[7\] systolic_inst.A_outs\[14\]\[7\] net120 VGND
+ VGND VPWR VPWR _00953_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23329_ _09955_ _09956_ _09944_ VGND VGND VPWR VPWR _09958_ sky130_fd_sc_hd__o21ai_1
X_27097_ clknet_leaf_7_B_in_serial_clk _00895_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26048_ deser_B.serial_word\[3\] deser_B.shift_reg\[3\] net55 VGND VGND VPWR VPWR
+ _03350_ sky130_fd_sc_hd__mux2_1
X_14062_ deser_B.shift_reg\[96\] deser_B.shift_reg\[97\] net126 VGND VGND VPWR VPWR
+ _00888_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18870_ _05973_ _05976_ _05979_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__a21oi_1
X_17821_ _05008_ _05018_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__or2_1
XFILLER_239_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27999_ clknet_leaf_152_clk _01797_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17752_ systolic_inst.acc_wires\[10\]\[24\] systolic_inst.acc_wires\[10\]\[25\] systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__o21a_1
X_14964_ _12041_ _12043_ _12042_ VGND VGND VPWR VPWR _12085_ sky130_fd_sc_hd__o21ba_1
XFILLER_235_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16703_ _04019_ _04023_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__xnor2_1
X_13915_ deser_A.serial_word\[76\] deser_A.shift_reg\[76\] net57 VGND VGND VPWR VPWR
+ _00741_ sky130_fd_sc_hd__mux2_1
X_29669_ clknet_leaf_27_B_in_serial_clk _03464_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[117\]
+ sky130_fd_sc_hd__dfrtp_1
X_17683_ _04916_ _04915_ systolic_inst.acc_wires\[10\]\[15\] net105 VGND VGND VPWR
+ VPWR _01313_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14895_ _11966_ _11967_ _11980_ _11979_ _11948_ VGND VGND VPWR VPWR _12018_ sky130_fd_sc_hd__o32a_1
XFILLER_208_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19422_ _06474_ _06475_ _06467_ _06471_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__a211o_1
XFILLER_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16634_ _03956_ _03957_ _03937_ _03940_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__o211ai_2
XFILLER_90_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13846_ deser_A.serial_word\[7\] deser_A.shift_reg\[7\] net58 VGND VGND VPWR VPWR
+ _00672_ sky130_fd_sc_hd__mux2_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19353_ _06348_ _06412_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_139_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13777_ B_in\[84\] deser_B.word_buffer\[84\] net85 VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__mux2_1
XFILLER_16_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16565_ _03906_ _03908_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__a21o_1
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18304_ _05469_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__nand2_1
XFILLER_43_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15516_ systolic_inst.B_outs\[13\]\[7\] _12540_ _12541_ VGND VGND VPWR VPWR _12574_
+ sky130_fd_sc_hd__a21bo_1
X_19284_ systolic_inst.B_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\] VGND VGND VPWR
+ VPWR _06346_ sky130_fd_sc_hd__or2_1
X_16496_ _03853_ _03854_ _03852_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__a21o_1
XFILLER_231_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18235_ net66 _05411_ _05413_ systolic_inst.acc_wires\[9\]\[6\] net107 VGND VGND
+ VPWR VPWR _01368_ sky130_fd_sc_hd__a32o_1
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15447_ _12506_ VGND VGND VPWR VPWR _12507_ sky130_fd_sc_hd__inv_2
XFILLER_54_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18166_ _05351_ _05352_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__nand2_1
X_15378_ net107 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _12442_ sky130_fd_sc_hd__and2_1
XFILLER_15_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17117_ _04406_ _04407_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__and2_1
Xmax_cap102 net103 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_12
Xmax_cap113 net114 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_12
X_14329_ _11476_ _11477_ _11479_ _11481_ _11475_ VGND VGND VPWR VPWR _11514_ sky130_fd_sc_hd__a32o_1
XFILLER_176_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap124 deser_B.serial_word_ready VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_130_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18097_ _05285_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__xnor2_1
Xmax_cap135 net153 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_130_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17048_ _04325_ _04348_ _04338_ _04347_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18999_ systolic_inst.acc_wires\[8\]\[28\] systolic_inst.acc_wires\[8\]\[29\] systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20961_ _07775_ _07808_ _07807_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__a21oi_1
XFILLER_241_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22700_ _09379_ _09385_ VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__xnor2_1
XFILLER_242_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23680_ _10297_ _10298_ VGND VGND VPWR VPWR _10299_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20892_ _07767_ _07768_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_85_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22631_ _09337_ _09339_ _09342_ net60 VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_234_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_2_1__leaf_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
X_25350_ net112 ser_C.shift_reg\[503\] VGND VGND VPWR VPWR _11145_ sky130_fd_sc_hd__and2_1
XFILLER_55_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22562_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[2\]\[14\]
+ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__nand2_1
XFILLER_194_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_230_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24301_ systolic_inst.A_shift\[12\]\[6\] A_in\[54\] net59 VGND VGND VPWR VPWR _10624_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_230_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21513_ systolic_inst.A_outs\[3\]\[1\] systolic_inst.B_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\]
+ systolic_inst.A_outs\[3\]\[0\] VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_230_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25281_ ser_C.parallel_data\[467\] net102 net74 ser_C.shift_reg\[467\] _11110_ VGND
+ VGND VPWR VPWR _02717_ sky130_fd_sc_hd__a221o_1
XFILLER_72_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22493_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[2\]\[4\]
+ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__or2_1
XFILLER_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27020_ clknet_leaf_23_B_in_serial_clk _00818_ net137 VGND VGND VPWR VPWR deser_B.shift_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24232_ _10601_ systolic_inst.A_shift\[19\]\[7\] net70 VGND VGND VPWR VPWR _02177_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21444_ _08279_ _08280_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__nand2_1
XFILLER_194_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24163_ systolic_inst.A_shift\[28\]\[5\] A_in\[101\] net59 VGND VGND VPWR VPWR _10583_
+ sky130_fd_sc_hd__mux2_1
X_21375_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[18\]
+ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__nand2_1
XFILLER_79_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23114_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[1\]\[7\]
+ VGND VGND VPWR VPWR _09780_ sky130_fd_sc_hd__or2_1
XFILLER_150_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20326_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[4\] _07263_ _07264_
+ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__nand4_2
XFILLER_150_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28971_ clknet_leaf_55_clk _02769_ VGND VGND VPWR VPWR systolic_inst.B_shift\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_24094_ _10556_ systolic_inst.B_shift\[19\]\[2\] net71 VGND VGND VPWR VPWR _02084_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_181_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27922_ clknet_leaf_145_clk _01720_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_23045_ _09691_ _09694_ _09719_ VGND VGND VPWR VPWR _09720_ sky130_fd_sc_hd__a21oi_1
X_20257_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[2\]
+ systolic_inst.A_outs\[5\]\[3\] VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__nand4_2
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27853_ clknet_leaf_36_clk _01651_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_88_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20188_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[26\]
+ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__nand2_1
XFILLER_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26804_ clknet_leaf_82_clk _00606_ net5 VGND VGND VPWR VPWR B_in\[76\] sky130_fd_sc_hd__dfrtp_1
XFILLER_48_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27784_ clknet_leaf_185_clk _01582_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_218_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24996_ net111 ser_C.shift_reg\[326\] VGND VGND VPWR VPWR _10968_ sky130_fd_sc_hd__and2_1
XFILLER_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29523_ clknet_leaf_260_clk _03321_ net140 VGND VGND VPWR VPWR ser_C.parallel_data\[495\]
+ sky130_fd_sc_hd__dfrtp_1
X_26735_ clknet_leaf_96_clk _00537_ net5 VGND VGND VPWR VPWR B_in\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23947_ _10502_ systolic_inst.B_shift\[10\]\[5\] _11332_ VGND VGND VPWR VPWR _01991_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13700_ B_in\[7\] deser_B.word_buffer\[7\] net84 VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__mux2_1
XFILLER_84_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29454_ clknet_leaf_289_clk _03252_ net136 VGND VGND VPWR VPWR C_out\[426\] sky130_fd_sc_hd__dfrtp_1
X_14680_ _11834_ _11835_ _11833_ VGND VGND VPWR VPWR _11836_ sky130_fd_sc_hd__o21ai_1
X_23878_ _11258_ systolic_inst.acc_wires\[0\]\[28\] net64 _10466_ VGND VGND VPWR VPWR
+ _01958_ sky130_fd_sc_hd__a22o_1
X_26666_ clknet_leaf_4_B_in_serial_clk _00469_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28405_ clknet_leaf_89_clk _02203_ VGND VGND VPWR VPWR systolic_inst.B_shift\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13631_ deser_B.word_buffer\[67\] deser_B.serial_word\[67\] net123 VGND VGND VPWR
+ VPWR _00468_ sky130_fd_sc_hd__mux2_1
XFILLER_32_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25617_ systolic_inst.acc_wires\[2\]\[29\] C_out\[93\] net50 VGND VGND VPWR VPWR
+ _02919_ sky130_fd_sc_hd__mux2_1
X_22829_ _09509_ _09510_ VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29385_ clknet_leaf_245_clk _03183_ net145 VGND VGND VPWR VPWR C_out\[357\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26597_ clknet_leaf_1_A_in_serial_clk _00400_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_213_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16350_ _03659_ _03706_ _03705_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__o21ba_1
X_28336_ clknet_leaf_343_clk _02134_ VGND VGND VPWR VPWR systolic_inst.A_shift\[26\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13562_ deser_A.shift_reg\[126\] deser_A.shift_reg\[127\] net130 VGND VGND VPWR VPWR
+ _00399_ sky130_fd_sc_hd__mux2_1
X_25548_ systolic_inst.acc_wires\[0\]\[24\] C_out\[24\] net53 VGND VGND VPWR VPWR
+ _02850_ sky130_fd_sc_hd__mux2_1
XFILLER_198_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_188_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_181_Right_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15301_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[23\]
+ VGND VGND VPWR VPWR _12392_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_188_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16281_ systolic_inst.A_outs\[12\]\[5\] systolic_inst.B_outs\[12\]\[6\] systolic_inst.A_outs\[12\]\[6\]
+ systolic_inst.B_outs\[12\]\[7\] VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__and4b_1
X_25479_ systolic_inst.ce_local _11215_ VGND VGND VPWR VPWR _11217_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_188_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28267_ clknet_leaf_78_clk _02065_ VGND VGND VPWR VPWR systolic_inst.B_shift\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13493_ deser_A.shift_reg\[57\] deser_A.shift_reg\[58\] net130 VGND VGND VPWR VPWR
+ _00330_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_160_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_160_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_199_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18020_ _05186_ _05211_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15232_ net61 _12333_ VGND VGND VPWR VPWR _12334_ sky130_fd_sc_hd__nor2_1
X_27218_ clknet_leaf_292_clk _01016_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_60_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28198_ clknet_leaf_48_clk _01996_ VGND VGND VPWR VPWR systolic_inst.B_shift\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15163_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[14\]\[3\]
+ VGND VGND VPWR VPWR _12274_ sky130_fd_sc_hd__and2_1
XFILLER_153_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27149_ clknet_leaf_276_clk _00947_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_197_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14114_ systolic_inst.B_shift\[12\]\[6\] net72 _11333_ B_in\[102\] VGND VGND VPWR
+ VPWR _00936_ sky130_fd_sc_hd__a22o_1
XFILLER_4_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19971_ _06923_ _06936_ _06934_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__o21a_1
X_15094_ _12179_ _12182_ _12210_ VGND VGND VPWR VPWR _12211_ sky130_fd_sc_hd__o21ai_1
XFILLER_180_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14045_ deser_B.shift_reg\[79\] deser_B.shift_reg\[80\] deser_B.receiving VGND VGND
+ VPWR VPWR _00871_ sky130_fd_sc_hd__mux2_1
XFILLER_180_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18922_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[18\]
+ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__or2_1
XFILLER_171_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18853_ net63 _05964_ _05965_ systolic_inst.acc_wires\[8\]\[8\] net108 VGND VGND
+ VPWR VPWR _01434_ sky130_fd_sc_hd__a32o_1
XFILLER_171_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17804_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__inv_2
XFILLER_212_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18784_ _05834_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15996_ systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[3\]
+ systolic_inst.B_outs\[12\]\[0\] VGND VGND VPWR VPWR _12995_ sky130_fd_sc_hd__a22o_1
XFILLER_208_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17735_ _04939_ _04946_ _04951_ _04956_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__nand4_1
XFILLER_212_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14947_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[8\] VGND
+ VGND VPWR VPWR _12069_ sky130_fd_sc_hd__and2_1
XFILLER_76_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17666_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[10\]\[12\]
+ _04898_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__and3_1
X_14878_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[5\] VGND VGND
+ VPWR VPWR _12001_ sky130_fd_sc_hd__nand2_1
XFILLER_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19405_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[7\]\[1\]
+ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__and2_1
XFILLER_224_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16617_ _03928_ _03930_ _03941_ net105 VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_173_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13829_ _11323_ _11324_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__nor2_1
XFILLER_63_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17597_ _04842_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_35_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19336_ _06394_ _06395_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__and2_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16548_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[27\]
+ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19267_ _06327_ _06328_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_151_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_151_clk
+ sky130_fd_sc_hd__clkbuf_8
X_16479_ _03839_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__inv_2
XFILLER_206_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18218_ _05397_ _05398_ _05390_ _05394_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__a211o_1
XFILLER_178_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19198_ _06262_ _06261_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__nand2b_1
XFILLER_129_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18149_ _05336_ _05335_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__and2b_1
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21160_ _07992_ _08027_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_44_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20111_ _07082_ _07089_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__nand2_1
X_21091_ _07923_ _07961_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__xor2_1
XFILLER_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20042_ _07030_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__inv_2
XFILLER_113_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24850_ net113 ser_C.shift_reg\[253\] VGND VGND VPWR VPWR _10895_ sky130_fd_sc_hd__and2_1
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23801_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[16\]
+ VGND VGND VPWR VPWR _10402_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24781_ C_out\[217\] net98 net78 ser_C.shift_reg\[217\] _10860_ VGND VGND VPWR VPWR
+ _02467_ sky130_fd_sc_hd__a221o_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_236_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21993_ _08766_ _08768_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__nand2_1
XFILLER_27_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_236_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_236_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23732_ _10340_ _10341_ _10342_ VGND VGND VPWR VPWR _10343_ sky130_fd_sc_hd__a21o_1
X_26520_ clknet_leaf_10_A_in_serial_clk _00323_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20944_ _07814_ _07818_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__xnor2_1
XFILLER_214_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_232_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_232_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[13\] _10282_ net122
+ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__mux2_1
X_26451_ clknet_leaf_10_clk _00258_ net132 VGND VGND VPWR VPWR A_in\[119\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_232_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20875_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\]
+ systolic_inst.A_outs\[4\]\[0\] VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__a22oi_1
X_22614_ _09321_ _09322_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__and2b_1
X_25402_ _11170_ systolic_inst.A_shift\[1\]\[0\] net71 VGND VGND VPWR VPWR _02778_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29170_ clknet_leaf_43_clk _02968_ net137 VGND VGND VPWR VPWR C_out\[142\] sky130_fd_sc_hd__dfrtp_1
X_26382_ clknet_leaf_19_clk _00189_ net133 VGND VGND VPWR VPWR A_in\[50\] sky130_fd_sc_hd__dfrtp_1
X_23594_ _10213_ _10214_ _10173_ _10176_ VGND VGND VPWR VPWR _10216_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_42_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28121_ clknet_leaf_125_clk _01919_ net144 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_25333_ ser_C.parallel_data\[493\] net97 net77 ser_C.shift_reg\[493\] _11136_ VGND
+ VGND VPWR VPWR _02743_ sky130_fd_sc_hd__a221o_1
X_22545_ _09260_ _09265_ _09266_ VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__nand3_1
XFILLER_194_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_142_clk clknet_5_25__leaf_clk VGND VGND VPWR VPWR clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28052_ clknet_leaf_51_clk _01850_ net143 VGND VGND VPWR VPWR systolic_inst.B_outs\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_25264_ net111 ser_C.shift_reg\[460\] VGND VGND VPWR VPWR _11102_ sky130_fd_sc_hd__and2_1
X_22476_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[2\]\[0\]
+ _09208_ _09209_ VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__a22o_1
XFILLER_154_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27003_ clknet_leaf_15_B_in_serial_clk _00801_ net152 VGND VGND VPWR VPWR deser_B.shift_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24215_ systolic_inst.A_shift\[21\]\[7\] A_in\[87\] net59 VGND VGND VPWR VPWR _10593_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21427_ net63 _08265_ _08266_ systolic_inst.acc_wires\[4\]\[25\] _11258_ VGND VGND
+ VPWR VPWR _01707_ sky130_fd_sc_hd__a32o_1
XFILLER_108_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25195_ C_out\[424\] net102 net74 ser_C.shift_reg\[424\] _11067_ VGND VGND VPWR VPWR
+ _02674_ sky130_fd_sc_hd__a221o_1
XFILLER_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24146_ _10574_ systolic_inst.A_shift\[28\]\[4\] net70 VGND VGND VPWR VPWR _02118_
+ sky130_fd_sc_hd__mux2_1
X_21358_ net63 _08206_ _08207_ systolic_inst.acc_wires\[4\]\[15\] _11258_ VGND VGND
+ VPWR VPWR _01697_ sky130_fd_sc_hd__a32o_1
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20309_ _07217_ _07220_ _07247_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__nor3_1
X_24077_ systolic_inst.B_shift\[3\]\[4\] _11332_ net83 systolic_inst.B_shift\[7\]\[4\]
+ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__a22o_1
X_28954_ clknet_leaf_262_clk _02752_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[502\]
+ sky130_fd_sc_hd__dfrtp_1
X_21289_ net63 _08146_ _08148_ systolic_inst.acc_wires\[4\]\[5\] net108 VGND VGND
+ VPWR VPWR _01687_ sky130_fd_sc_hd__a32o_1
XFILLER_81_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23028_ _09702_ _09703_ VGND VGND VPWR VPWR _09704_ sky130_fd_sc_hd__nor2_1
X_27905_ clknet_leaf_138_clk _01703_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28885_ clknet_leaf_331_clk _02683_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[433\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27836_ clknet_leaf_206_clk _01634_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15850_ _12881_ _12884_ VGND VGND VPWR VPWR _12886_ sky130_fd_sc_hd__or2_1
XFILLER_130_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _11905_ _11908_ _11926_ VGND VGND VPWR VPWR _11927_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_177_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27767_ clknet_leaf_208_clk _01565_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15781_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[13\]\[5\]
+ VGND VGND VPWR VPWR _12826_ sky130_fd_sc_hd__nand2_1
X_24979_ C_out\[316\] net97 net80 ser_C.shift_reg\[316\] _10959_ VGND VGND VPWR VPWR
+ _02566_ sky130_fd_sc_hd__a221o_1
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29506_ clknet_leaf_265_clk _03304_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17520_ systolic_inst.A_outs\[10\]\[6\] _11275_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__nor2_1
X_26718_ clknet_leaf_29_B_in_serial_clk _00521_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_14732_ _11878_ _11879_ VGND VGND VPWR VPWR _11880_ sky130_fd_sc_hd__nand2_1
XFILLER_233_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27698_ clknet_leaf_197_clk _01496_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29437_ clknet_leaf_335_clk _03235_ net131 VGND VGND VPWR VPWR C_out\[409\] sky130_fd_sc_hd__dfrtp_1
X_17451_ net105 _04704_ _04705_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__or3_1
XFILLER_166_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26649_ clknet_leaf_20_B_in_serial_clk _00452_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ _11819_ _11820_ VGND VGND VPWR VPWR _11821_ sky130_fd_sc_hd__and2_1
XFILLER_33_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16402_ net67 _03771_ _03773_ systolic_inst.acc_wires\[12\]\[5\] net108 VGND VGND
+ VPWR VPWR _01175_ sky130_fd_sc_hd__a32o_1
X_13614_ deser_B.word_buffer\[50\] deser_B.serial_word\[50\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__mux2_1
X_29368_ clknet_leaf_232_clk _03166_ net147 VGND VGND VPWR VPWR C_out\[340\] sky130_fd_sc_hd__dfrtp_1
X_17382_ _04599_ _04605_ _04604_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__a21o_1
XFILLER_207_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14594_ _11760_ _11761_ VGND VGND VPWR VPWR _11762_ sky130_fd_sc_hd__and2_1
XFILLER_242_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19121_ _06186_ _06187_ _06175_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__or3b_1
X_16333_ _03711_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__xnor2_1
X_28319_ clknet_leaf_0_clk _02117_ VGND VGND VPWR VPWR systolic_inst.A_shift\[28\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13545_ deser_A.shift_reg\[109\] deser_A.shift_reg\[110\] net129 VGND VGND VPWR VPWR
+ _00382_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_133_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_9_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29299_ clknet_leaf_312_clk _03097_ net141 VGND VGND VPWR VPWR C_out\[271\] sky130_fd_sc_hd__dfrtp_1
XFILLER_125_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19052_ _06108_ _06110_ _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__and3_1
XFILLER_51_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16264_ _03629_ _03645_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__xor2_1
X_13476_ deser_A.shift_reg\[40\] deser_A.shift_reg\[41\] net130 VGND VGND VPWR VPWR
+ _00313_ sky130_fd_sc_hd__mux2_1
XFILLER_9_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18003_ _05191_ _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__xnor2_1
X_15215_ _12316_ _12318_ VGND VGND VPWR VPWR _12319_ sky130_fd_sc_hd__xor2_1
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16195_ _03578_ _03577_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_11_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15146_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[14\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _12260_ sky130_fd_sc_hd__a21o_1
XFILLER_154_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19954_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[12\] _06950_ net119
+ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__mux2_1
X_15077_ _12193_ _12194_ VGND VGND VPWR VPWR _12195_ sky130_fd_sc_hd__nor2_1
XFILLER_142_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14028_ deser_B.shift_reg\[62\] deser_B.shift_reg\[63\] net126 VGND VGND VPWR VPWR
+ _00854_ sky130_fd_sc_hd__mux2_1
X_18905_ net63 _06009_ _06010_ systolic_inst.acc_wires\[8\]\[15\] net108 VGND VGND
+ VPWR VPWR _01441_ sky130_fd_sc_hd__a32o_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19885_ _06881_ _06882_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__xor2_1
XFILLER_136_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18836_ net63 _05949_ _05951_ systolic_inst.acc_wires\[8\]\[5\] net108 VGND VGND
+ VPWR VPWR _01431_ sky130_fd_sc_hd__a32o_1
XFILLER_67_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18767_ net117 _05889_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_121_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15979_ net115 _12979_ VGND VGND VPWR VPWR _12980_ sky130_fd_sc_hd__nand2_1
XFILLER_76_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17718_ _04945_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18698_ _05764_ _05823_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17649_ _04876_ _04881_ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__a21oi_1
XFILLER_224_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20660_ _07580_ _07581_ _07582_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__a21o_1
XFILLER_211_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19319_ systolic_inst.B_outs\[7\]\[5\] systolic_inst.A_outs\[7\]\[7\] VGND VGND VPWR
+ VPWR _06380_ sky130_fd_sc_hd__nand2_1
XFILLER_143_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_124_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20591_ _11276_ systolic_inst.A_outs\[5\]\[7\] _07469_ _07494_ VGND VGND VPWR VPWR
+ _07522_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_119_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22330_ _09071_ _09072_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__nand2_1
XFILLER_108_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22261_ _09004_ _09005_ VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_22_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24000_ _10525_ systolic_inst.B_shift\[5\]\[3\] _11332_ VGND VGND VPWR VPWR _02021_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21212_ _08077_ _08078_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22192_ _08915_ _08937_ _08938_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__and3_1
XFILLER_191_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_225_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21143_ _08011_ _08012_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__and2b_1
XFILLER_219_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25951_ systolic_inst.acc_wires\[13\]\[11\] C_out\[427\] net19 VGND VGND VPWR VPWR
+ _03253_ sky130_fd_sc_hd__mux2_1
X_21074_ _07903_ _07905_ _07945_ VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_238_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20025_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[6\]\[0\]
+ _07010_ _07008_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__a31o_1
XFILLER_24_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24902_ net110 ser_C.shift_reg\[279\] VGND VGND VPWR VPWR _10921_ sky130_fd_sc_hd__and2_1
X_28670_ clknet_leaf_187_clk _02468_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[218\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25882_ systolic_inst.acc_wires\[11\]\[6\] C_out\[358\] net38 VGND VGND VPWR VPWR
+ _03184_ sky130_fd_sc_hd__mux2_1
XFILLER_101_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27621_ clknet_leaf_315_clk _01419_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24833_ C_out\[243\] net98 net78 ser_C.shift_reg\[243\] _10886_ VGND VGND VPWR VPWR
+ _02493_ sky130_fd_sc_hd__a221o_1
XFILLER_115_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_61_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27552_ clknet_leaf_299_clk _01350_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_21976_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[3\]\[14\]
+ _08752_ VGND VGND VPWR VPWR _08761_ sky130_fd_sc_hd__and3_1
X_24764_ net113 ser_C.shift_reg\[210\] VGND VGND VPWR VPWR _10852_ sky130_fd_sc_hd__and2_1
Xclkbuf_5_2__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26503_ clknet_leaf_15_A_in_serial_clk _00306_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_23715_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[0\]\[4\]
+ VGND VGND VPWR VPWR _10328_ sky130_fd_sc_hd__nand2_1
X_20927_ _07780_ _07782_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__nand2_1
X_24695_ C_out\[174\] net104 net76 ser_C.shift_reg\[174\] _10817_ VGND VGND VPWR VPWR
+ _02424_ sky130_fd_sc_hd__a221o_1
X_27483_ clknet_leaf_41_clk _01281_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_70_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29222_ clknet_leaf_210_clk _03020_ net147 VGND VGND VPWR VPWR C_out\[194\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26434_ clknet_leaf_1_clk _00241_ net131 VGND VGND VPWR VPWR A_in\[102\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23646_ _10256_ _10265_ VGND VGND VPWR VPWR _10266_ sky130_fd_sc_hd__nor2_1
XFILLER_70_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20858_ net108 systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[2\] _07734_
+ _07736_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__a22o_1
XFILLER_109_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_999 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29153_ clknet_leaf_172_clk _02951_ net148 VGND VGND VPWR VPWR C_out\[125\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_115_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
X_23577_ _10197_ _10198_ VGND VGND VPWR VPWR _10199_ sky130_fd_sc_hd__nor2_1
X_26365_ clknet_leaf_25_clk _00172_ net137 VGND VGND VPWR VPWR A_in\[33\] sky130_fd_sc_hd__dfrtp_1
XFILLER_195_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20789_ _07687_ _07689_ _07691_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__o21ai_1
XFILLER_161_1254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28104_ clknet_leaf_156_clk _01902_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13330_ A_in\[39\] deser_A.word_buffer\[39\] net93 VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__mux2_1
X_22528_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[2\]\[8\]
+ _09252_ VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__and3_1
XFILLER_195_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25316_ net112 ser_C.shift_reg\[486\] VGND VGND VPWR VPWR _11128_ sky130_fd_sc_hd__and2_1
X_29084_ clknet_leaf_111_clk _02882_ net151 VGND VGND VPWR VPWR C_out\[56\] sky130_fd_sc_hd__dfrtp_1
XFILLER_194_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26296_ clknet_leaf_27_A_in_serial_clk _00104_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_70_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_210_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28035_ clknet_leaf_158_clk _01833_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_210_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ deser_A.word_buffer\[99\] deser_A.serial_word\[99\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__mux2_1
X_22459_ _09196_ _09197_ VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__xor2_1
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25247_ ser_C.parallel_data\[450\] net102 net74 ser_C.shift_reg\[450\] _11093_ VGND
+ VGND VPWR VPWR _02700_ sky130_fd_sc_hd__a221o_1
XFILLER_202_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15000_ _12111_ _12119_ VGND VGND VPWR VPWR _12120_ sky130_fd_sc_hd__nand2_1
XFILLER_108_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25178_ net110 ser_C.shift_reg\[417\] VGND VGND VPWR VPWR _11059_ sky130_fd_sc_hd__and2_1
X_13192_ deser_A.word_buffer\[30\] deser_A.serial_word\[30\] net128 VGND VGND VPWR
+ VPWR _00040_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24129_ systolic_inst.A_shift\[30\]\[4\] A_in\[116\] net59 VGND VGND VPWR VPWR _10566_
+ sky130_fd_sc_hd__mux2_1
XFILLER_237_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28937_ clknet_leaf_260_clk _02735_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[485\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16951_ _04263_ _04264_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__and2b_1
XFILLER_173_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15902_ _12926_ _12927_ _12928_ VGND VGND VPWR VPWR _12930_ sky130_fd_sc_hd__or3_1
XFILLER_133_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19670_ _06668_ _06674_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__nor2_1
XFILLER_77_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28868_ clknet_leaf_300_clk _02666_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[416\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16882_ _04197_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__nand2_1
XFILLER_237_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18621_ _05704_ _05712_ _05711_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__a21o_1
X_27819_ clknet_leaf_144_clk _01617_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_15833_ _12867_ _12868_ _12869_ VGND VGND VPWR VPWR _12871_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28799_ clknet_leaf_235_clk _02597_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18552_ _05643_ _05645_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__and2b_1
XFILLER_92_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15764_ _12808_ _12809_ _12810_ VGND VGND VPWR VPWR _12812_ sky130_fd_sc_hd__and3_1
XFILLER_92_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17503_ _04742_ _04755_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__xnor2_1
X_14715_ systolic_inst.acc_wires\[15\]\[26\] systolic_inst.acc_wires\[15\]\[27\] systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _11865_ sky130_fd_sc_hd__o21a_1
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18483_ _05606_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_159_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15695_ _12746_ _12747_ VGND VGND VPWR VPWR _12748_ sky130_fd_sc_hd__xnor2_1
X_17434_ _04687_ _04688_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__nand2_1
X_14646_ _11806_ VGND VGND VPWR VPWR _11807_ sky130_fd_sc_hd__inv_2
XFILLER_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_106_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_19 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17365_ _04544_ _04581_ _04583_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__a21oi_1
XFILLER_207_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14577_ _11745_ _11746_ _11747_ VGND VGND VPWR VPWR _11748_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_109_Left_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19104_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[5\]
+ systolic_inst.A_outs\[7\]\[6\] VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__and4_1
X_16316_ _03694_ _03695_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__and2_1
XFILLER_201_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13528_ deser_A.shift_reg\[92\] deser_A.shift_reg\[93\] net129 VGND VGND VPWR VPWR
+ _00365_ sky130_fd_sc_hd__mux2_1
XFILLER_173_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17296_ _04552_ _04553_ _04530_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19035_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[1\]
+ systolic_inst.A_outs\[7\]\[2\] VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__and4_1
XFILLER_185_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16247_ _03627_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__nand2_1
XFILLER_220_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13459_ deser_A.shift_reg\[23\] deser_A.shift_reg\[24\] deser_A.receiving VGND VGND
+ VPWR VPWR _00296_ sky130_fd_sc_hd__mux2_1
XFILLER_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16178_ systolic_inst.B_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[5\]
+ systolic_inst.A_outs\[12\]\[6\] VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__and4_1
XFILLER_86_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15129_ _12243_ _12244_ VGND VGND VPWR VPWR _12245_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19937_ _06902_ _06904_ _06933_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__a21o_1
XFILLER_151_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Left_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19868_ _06866_ _06865_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__nand2b_1
XFILLER_29_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18819_ _05935_ _05936_ _05928_ _05932_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__a211o_1
X_19799_ _06797_ _06798_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_108_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21830_ _08584_ _08633_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_69_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21761_ _08528_ _08530_ _08566_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_218_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_345_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_345_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20712_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[5\]\[14\]
+ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__or2_1
X_23500_ systolic_inst.A_outs\[0\]\[6\] _10080_ _10079_ _10078_ VGND VGND VPWR VPWR
+ _10124_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24480_ net112 ser_C.shift_reg\[68\] VGND VGND VPWR VPWR _10710_ sky130_fd_sc_hd__and2_1
XFILLER_169_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21692_ _08459_ _08461_ _08498_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__nand3_1
XFILLER_145_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_127_Left_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23431_ _10054_ _10055_ _09993_ _09996_ VGND VGND VPWR VPWR _10057_ sky130_fd_sc_hd__o211a_1
X_20643_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[5\]\[4\]
+ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__nand2_1
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26150_ deser_B.serial_word\[105\] deser_B.shift_reg\[105\] _00001_ VGND VGND VPWR
+ VPWR _03452_ sky130_fd_sc_hd__mux2_1
XFILLER_177_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23362_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[5\] _09989_ net121
+ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__mux2_1
XFILLER_149_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20574_ _07504_ _07505_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_227_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22313_ _08985_ _09055_ VGND VGND VPWR VPWR _09056_ sky130_fd_sc_hd__nor2_1
X_25101_ C_out\[377\] net98 net78 ser_C.shift_reg\[377\] _11020_ VGND VGND VPWR VPWR
+ _02627_ sky130_fd_sc_hd__a221o_1
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26081_ deser_B.serial_word\[36\] deser_B.shift_reg\[36\] net55 VGND VGND VPWR VPWR
+ _03383_ sky130_fd_sc_hd__mux2_1
X_23293_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[2\] _09922_ _09923_
+ VGND VGND VPWR VPWR _09924_ sky130_fd_sc_hd__and4_1
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25032_ net112 ser_C.shift_reg\[344\] VGND VGND VPWR VPWR _10986_ sky130_fd_sc_hd__and2_1
X_22244_ _08982_ _08988_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22175_ _08894_ _08921_ VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__xor2_1
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21126_ _07955_ _07994_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__nand2_1
XFILLER_105_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26983_ clknet_leaf_29_A_in_serial_clk _00781_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28722_ clknet_leaf_311_clk _02520_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[270\]
+ sky130_fd_sc_hd__dfrtp_1
X_21057_ systolic_inst.A_outs\[4\]\[2\] _07852_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__nor2_1
X_25934_ systolic_inst.acc_wires\[12\]\[26\] C_out\[410\] net21 VGND VGND VPWR VPWR
+ _03236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20008_ _06921_ _06981_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_203_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28653_ clknet_leaf_203_clk _02451_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[201\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25865_ systolic_inst.acc_wires\[10\]\[21\] C_out\[341\] net11 VGND VGND VPWR VPWR
+ _03167_ sky130_fd_sc_hd__mux2_1
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27604_ clknet_leaf_202_clk _01402_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_24816_ net113 ser_C.shift_reg\[236\] VGND VGND VPWR VPWR _10878_ sky130_fd_sc_hd__and2_1
X_28584_ clknet_leaf_309_clk _02382_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25796_ systolic_inst.acc_wires\[8\]\[16\] C_out\[272\] net28 VGND VGND VPWR VPWR
+ _03098_ sky130_fd_sc_hd__mux2_1
XFILLER_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27535_ clknet_leaf_316_clk _01333_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_24747_ C_out\[200\] net97 net80 ser_C.shift_reg\[200\] _10843_ VGND VGND VPWR VPWR
+ _02450_ sky130_fd_sc_hd__a221o_1
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21959_ net68 _08745_ _08746_ systolic_inst.acc_wires\[3\]\[13\] net106 VGND VGND
+ VPWR VPWR _01759_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_336_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_336_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14500_ _11593_ _11679_ VGND VGND VPWR VPWR _11680_ sky130_fd_sc_hd__or2_1
XFILLER_226_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27466_ clknet_leaf_236_clk _01264_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_15480_ _12515_ _12517_ VGND VGND VPWR VPWR _12539_ sky130_fd_sc_hd__nand2_1
XFILLER_242_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24678_ net111 ser_C.shift_reg\[167\] VGND VGND VPWR VPWR _10809_ sky130_fd_sc_hd__and2_1
XFILLER_15_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29205_ clknet_leaf_207_clk _03003_ net147 VGND VGND VPWR VPWR C_out\[177\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_212_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14431_ _11575_ _11578_ _11612_ VGND VGND VPWR VPWR _11614_ sky130_fd_sc_hd__and3_1
X_26417_ clknet_leaf_7_clk _00224_ net133 VGND VGND VPWR VPWR A_in\[85\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_212_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ _10246_ _10247_ _10249_ VGND VGND VPWR VPWR _10250_ sky130_fd_sc_hd__and3_1
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27397_ clknet_leaf_335_clk _01195_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29136_ clknet_leaf_168_clk _02934_ net148 VGND VGND VPWR VPWR C_out\[108\] sky130_fd_sc_hd__dfrtp_1
X_17150_ _04429_ _04433_ _04430_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26348_ clknet_leaf_63_clk _00155_ net135 VGND VGND VPWR VPWR A_in\[16\] sky130_fd_sc_hd__dfrtp_1
X_14362_ _11545_ _11513_ VGND VGND VPWR VPWR _11547_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_150_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16101_ systolic_inst.B_outs\[12\]\[3\] systolic_inst.A_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\]
+ systolic_inst.A_outs\[12\]\[4\] VGND VGND VPWR VPWR _13096_ sky130_fd_sc_hd__and4_1
X_13313_ A_in\[22\] deser_A.word_buffer\[22\] net91 VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__mux2_1
X_29067_ clknet_leaf_115_clk _02865_ net149 VGND VGND VPWR VPWR C_out\[39\] sky130_fd_sc_hd__dfrtp_1
X_14293_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[6\]
+ systolic_inst.A_outs\[15\]\[7\] VGND VGND VPWR VPWR _11479_ sky130_fd_sc_hd__nand4_1
X_17081_ _04376_ _04377_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__nand2_1
XFILLER_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26279_ clknet_leaf_20_A_in_serial_clk _00087_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_100_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28018_ clknet_leaf_154_clk _01816_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16032_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[4\]
+ systolic_inst.A_outs\[12\]\[5\] VGND VGND VPWR VPWR _13029_ sky130_fd_sc_hd__and4_1
X_13244_ deser_A.word_buffer\[82\] deser_A.serial_word\[82\] net127 VGND VGND VPWR
+ VPWR _00092_ sky130_fd_sc_hd__mux2_1
XFILLER_155_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13175_ deser_A.word_buffer\[13\] deser_A.serial_word\[13\] net127 VGND VGND VPWR
+ VPWR _00023_ sky130_fd_sc_hd__mux2_1
XFILLER_108_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17983_ _05173_ _05174_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__xor2_1
XFILLER_111_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19722_ systolic_inst.A_outs\[6\]\[1\] systolic_inst.B_outs\[6\]\[5\] systolic_inst.B_outs\[6\]\[6\]
+ systolic_inst.A_outs\[6\]\[0\] VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__a22oi_1
X_16934_ _04248_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__and2b_1
XFILLER_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19653_ _06652_ _06658_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16865_ _04166_ _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__xor2_1
XFILLER_238_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18604_ _05695_ _05731_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__nor2_1
X_15816_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[13\]\[9\]
+ _12851_ VGND VGND VPWR VPWR _12856_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19584_ _06607_ _06611_ _06608_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__a21bo_1
X_16796_ _04096_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__xor2_1
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18535_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[5\] VGND VGND VPWR
+ VPWR _05665_ sky130_fd_sc_hd__nand2_1
XFILLER_209_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _12794_ _12797_ VGND VGND VPWR VPWR _12798_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_327_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_327_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18466_ _05579_ _05596_ _05597_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__and3_1
XFILLER_233_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15678_ _12731_ _12730_ VGND VGND VPWR VPWR _12732_ sky130_fd_sc_hd__and2b_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17417_ _04602_ _04671_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__nor2_1
XFILLER_178_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14629_ _11788_ _11791_ VGND VGND VPWR VPWR _11793_ sky130_fd_sc_hd__or2_1
XFILLER_53_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18397_ _05547_ _05550_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17348_ _04600_ _04603_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload200 clknet_leaf_68_clk VGND VGND VPWR VPWR clkload200/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload211 clknet_leaf_45_clk VGND VGND VPWR VPWR clkload211/Y sky130_fd_sc_hd__clkinv_2
XFILLER_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17279_ systolic_inst.A_outs\[10\]\[2\] systolic_inst.B_outs\[10\]\[3\] systolic_inst.A_outs\[10\]\[3\]
+ systolic_inst.B_outs\[10\]\[4\] VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__nand4_2
XFILLER_174_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload222 clknet_leaf_128_clk VGND VGND VPWR VPWR clkload222/Y sky130_fd_sc_hd__bufinv_16
Xclkload233 clknet_leaf_84_clk VGND VGND VPWR VPWR clkload233/Y sky130_fd_sc_hd__clkinv_4
XFILLER_220_1181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19018_ systolic_inst.A_outs\[7\]\[7\] systolic_inst.A_outs\[6\]\[7\] net119 VGND
+ VGND VPWR VPWR _01465_ sky130_fd_sc_hd__mux2_1
Xclkload244 clknet_leaf_97_clk VGND VGND VPWR VPWR clkload244/X sky130_fd_sc_hd__clkbuf_8
XFILLER_228_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload255 clknet_leaf_94_clk VGND VGND VPWR VPWR clkload255/Y sky130_fd_sc_hd__clkinv_4
X_20290_ systolic_inst.B_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[4\]
+ systolic_inst.A_outs\[5\]\[5\] VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__and4_1
Xclkload266 clknet_leaf_133_clk VGND VGND VPWR VPWR clkload266/Y sky130_fd_sc_hd__inv_6
XFILLER_173_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload277 clknet_leaf_146_clk VGND VGND VPWR VPWR clkload277/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload288 clknet_leaf_192_clk VGND VGND VPWR VPWR clkload288/Y sky130_fd_sc_hd__clkinv_4
Xclkload299 clknet_leaf_179_clk VGND VGND VPWR VPWR clkload299/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_142_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23980_ _10515_ systolic_inst.B_shift\[8\]\[1\] net72 VGND VGND VPWR VPWR _02011_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22931_ _09607_ _09608_ VGND VGND VPWR VPWR _09610_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25650_ systolic_inst.acc_wires\[3\]\[30\] C_out\[126\] net49 VGND VGND VPWR VPWR
+ _02952_ sky130_fd_sc_hd__mux2_1
X_22862_ _09512_ _09542_ VGND VGND VPWR VPWR _09543_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_216_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24601_ C_out\[127\] net99 net80 ser_C.shift_reg\[127\] _10770_ VGND VGND VPWR VPWR
+ _02377_ sky130_fd_sc_hd__a221o_1
X_21813_ _08615_ _08616_ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__xnor2_1
X_25581_ systolic_inst.acc_wires\[1\]\[25\] C_out\[57\] net52 VGND VGND VPWR VPWR
+ _02883_ sky130_fd_sc_hd__mux2_1
XFILLER_227_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22793_ _09474_ _09475_ VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_318_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_318_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_145_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27320_ clknet_leaf_289_clk _01118_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24532_ net114 ser_C.shift_reg\[94\] VGND VGND VPWR VPWR _10736_ sky130_fd_sc_hd__and2_1
X_21744_ systolic_inst.A_outs\[3\]\[6\] _08519_ _08520_ _08485_ VGND VGND VPWR VPWR
+ _08550_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_227_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27251_ clknet_leaf_275_clk _01049_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24463_ C_out\[58\] net100 net82 ser_C.shift_reg\[58\] _10701_ VGND VGND VPWR VPWR
+ _02308_ sky130_fd_sc_hd__a221o_1
X_21675_ _08443_ _08481_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__and2_1
XFILLER_169_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26202_ clknet_leaf_15_A_in_serial_clk _00010_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23414_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[5\]
+ systolic_inst.A_outs\[0\]\[6\] VGND VGND VPWR VPWR _10040_ sky130_fd_sc_hd__and4_1
X_20626_ _07553_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__inv_2
X_24394_ net7 ser_C.shift_reg\[25\] VGND VGND VPWR VPWR _10667_ sky130_fd_sc_hd__and2_1
X_27182_ clknet_leaf_265_clk _00980_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23345_ _09946_ _09971_ _09972_ VGND VGND VPWR VPWR _09973_ sky130_fd_sc_hd__a21o_1
X_26133_ deser_B.serial_word\[88\] deser_B.shift_reg\[88\] net56 VGND VGND VPWR VPWR
+ _03435_ sky130_fd_sc_hd__mux2_1
X_20557_ _07422_ _07427_ _07457_ _07456_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__a31o_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23276_ _09917_ _09916_ systolic_inst.acc_wires\[1\]\[31\] net109 VGND VGND VPWR
+ VPWR _01905_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_180_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26064_ deser_B.serial_word\[19\] deser_B.shift_reg\[19\] net55 VGND VGND VPWR VPWR
+ _03366_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20488_ _07420_ _07421_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__nand2_1
XFILLER_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22227_ _08972_ _08971_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__nand2b_1
XFILLER_180_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25015_ C_out\[334\] net97 net80 ser_C.shift_reg\[334\] _10977_ VGND VGND VPWR VPWR
+ _02584_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_56_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22158_ _08897_ _08905_ VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__nor2_1
XFILLER_152_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_205_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21109_ _07952_ _07978_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__xnor2_1
X_22089_ systolic_inst.B_outs\[1\]\[3\] systolic_inst.B_shift\[1\]\[3\] net122 VGND
+ VGND VPWR VPWR _01789_ sky130_fd_sc_hd__mux2_1
X_14980_ _12098_ _12099_ VGND VGND VPWR VPWR _12101_ sky130_fd_sc_hd__nand2_1
X_26966_ clknet_leaf_23_A_in_serial_clk _00764_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28705_ clknet_leaf_185_clk _02503_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[253\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_197_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25917_ systolic_inst.acc_wires\[12\]\[9\] C_out\[393\] net17 VGND VGND VPWR VPWR
+ _03219_ sky130_fd_sc_hd__mux2_1
X_13931_ deser_A.serial_word\[92\] deser_A.shift_reg\[92\] net57 VGND VGND VPWR VPWR
+ _00757_ sky130_fd_sc_hd__mux2_1
X_29685_ clknet_leaf_105_clk _03480_ net152 VGND VGND VPWR VPWR ser_C.bit_idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_197_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26897_ clknet_leaf_6_A_in_serial_clk _00695_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28636_ clknet_leaf_181_clk _02434_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[184\]
+ sky130_fd_sc_hd__dfrtp_1
X_16650_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[3\] _03970_ _03971_
+ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__o2bb2a_1
X_13862_ deser_A.serial_word\[23\] deser_A.shift_reg\[23\] net58 VGND VGND VPWR VPWR
+ _00688_ sky130_fd_sc_hd__mux2_1
X_25848_ systolic_inst.acc_wires\[10\]\[4\] C_out\[324\] net14 VGND VGND VPWR VPWR
+ _03150_ sky130_fd_sc_hd__mux2_1
XFILLER_16_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15601_ _12656_ _12655_ VGND VGND VPWR VPWR _12657_ sky130_fd_sc_hd__nand2b_1
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28567_ clknet_leaf_165_clk _02365_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[115\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_309_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_309_clk
+ sky130_fd_sc_hd__clkbuf_8
X_16581_ systolic_inst.A_outs\[11\]\[6\] systolic_inst.A_outs\[10\]\[6\] net118 VGND
+ VGND VPWR VPWR _01208_ sky130_fd_sc_hd__mux2_1
X_13793_ B_in\[100\] deser_B.word_buffer\[100\] _00005_ VGND VGND VPWR VPWR _00630_
+ sky130_fd_sc_hd__mux2_1
X_25779_ systolic_inst.acc_wires\[7\]\[31\] C_out\[255\] net43 VGND VGND VPWR VPWR
+ _03081_ sky130_fd_sc_hd__mux2_1
XFILLER_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18320_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[19\]
+ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27518_ clknet_leaf_201_clk _01316_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_15532_ _12588_ _12589_ VGND VGND VPWR VPWR _12590_ sky130_fd_sc_hd__and2b_1
XFILLER_215_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28498_ clknet_leaf_117_clk _02296_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18251_ _05425_ _05426_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__or2_1
XFILLER_31_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15463_ _12517_ _12518_ _12522_ VGND VGND VPWR VPWR _12523_ sky130_fd_sc_hd__nand3_2
X_27449_ clknet_leaf_235_clk _01247_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_231_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17202_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.A_outs\[10\]\[2\] VGND VGND
+ VPWR VPWR _04465_ sky130_fd_sc_hd__nand2_1
X_14414_ _11595_ _11596_ VGND VGND VPWR VPWR _11597_ sky130_fd_sc_hd__or2_1
XFILLER_129_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18182_ _05342_ _05366_ _05367_ _05365_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__o31ai_1
X_15394_ _12455_ _12456_ VGND VGND VPWR VPWR _12457_ sky130_fd_sc_hd__and2_1
XFILLER_204_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29119_ clknet_leaf_163_clk _02917_ net151 VGND VGND VPWR VPWR C_out\[91\] sky130_fd_sc_hd__dfrtp_1
X_17133_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[24\]
+ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__and2_1
XFILLER_156_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14345_ systolic_inst.A_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[6\] VGND VGND
+ VPWR VPWR _11530_ sky130_fd_sc_hd__nand2_1
XFILLER_11_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17064_ _04361_ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__and2_1
XFILLER_170_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14276_ _11419_ _11460_ VGND VGND VPWR VPWR _11463_ sky130_fd_sc_hd__xor2_1
XFILLER_143_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16015_ _12991_ _13012_ VGND VGND VPWR VPWR _13013_ sky130_fd_sc_hd__xnor2_1
X_13227_ deser_A.word_buffer\[65\] deser_A.serial_word\[65\] net127 VGND VGND VPWR
+ VPWR _00075_ sky130_fd_sc_hd__mux2_1
XFILLER_170_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13158_ deser_B.serial_toggle_sync2 deser_B.serial_toggle_sync1 VGND VGND VPWR VPWR
+ _00005_ sky130_fd_sc_hd__xor2_4
XFILLER_151_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17966_ _05157_ _05158_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19705_ _06661_ _06680_ _06679_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__a21bo_1
X_16917_ _04201_ _04204_ _04202_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_105_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17897_ systolic_inst.A_outs\[9\]\[1\] systolic_inst.B_outs\[9\]\[5\] systolic_inst.B_outs\[9\]\[6\]
+ systolic_inst.A_outs\[9\]\[0\] VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__a22oi_1
XFILLER_211_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19636_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[1\]
+ systolic_inst.A_outs\[6\]\[2\] VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__and4_1
X_16848_ _04164_ _04165_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__nand2_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_195_Right_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19567_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[24\]
+ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__and2_1
XFILLER_241_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16779_ systolic_inst.B_outs\[11\]\[3\] systolic_inst.B_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[5\]
+ systolic_inst.A_outs\[11\]\[6\] VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__and4_1
XFILLER_179_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18518_ _05625_ _05647_ _05648_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_17_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19498_ _06539_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__and2_1
XFILLER_179_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18449_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.A_outs\[8\]\[1\] systolic_inst.B_outs\[8\]\[3\]
+ systolic_inst.B_outs\[8\]\[4\] VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__nand4_1
X_21460_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[31\]
+ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_135_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20411_ _07346_ _07347_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_135_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21391_ _08211_ _08235_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__nor2_1
XFILLER_119_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23130_ _09789_ _09791_ _09793_ systolic_inst.acc_wires\[1\]\[9\] net109 VGND VGND
+ VPWR VPWR _01883_ sky130_fd_sc_hd__a32o_1
XFILLER_190_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20342_ _07246_ _07248_ _07279_ _07280_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__o211a_1
XFILLER_88_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23061_ _09516_ _09652_ _09727_ _09725_ VGND VGND VPWR VPWR _09735_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_92_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20273_ systolic_inst.B_outs\[5\]\[1\] systolic_inst.A_outs\[5\]\[3\] systolic_inst.A_outs\[5\]\[4\]
+ systolic_inst.B_outs\[5\]\[0\] VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22012_ _08783_ _08789_ _08790_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_241_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_241_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26820_ clknet_leaf_69_clk _00622_ net135 VGND VGND VPWR VPWR B_in\[92\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26751_ clknet_leaf_56_clk _00553_ net137 VGND VGND VPWR VPWR B_in\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_112_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23963_ systolic_inst.B_shift\[13\]\[1\] B_in\[41\] _00008_ VGND VGND VPWR VPWR _10507_
+ sky130_fd_sc_hd__mux2_1
XFILLER_217_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_95_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_151_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25702_ systolic_inst.acc_wires\[5\]\[18\] C_out\[178\] net45 VGND VGND VPWR VPWR
+ _03004_ sky130_fd_sc_hd__mux2_1
X_22914_ systolic_inst.B_outs\[1\]\[5\] systolic_inst.A_outs\[1\]\[5\] VGND VGND VPWR
+ VPWR _09593_ sky130_fd_sc_hd__nand2_1
X_29470_ clknet_leaf_286_clk _03268_ net136 VGND VGND VPWR VPWR ser_C.parallel_data\[442\]
+ sky130_fd_sc_hd__dfrtp_1
X_26682_ clknet_leaf_25_B_in_serial_clk _00485_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_23894_ _10473_ _10477_ _10478_ _11713_ VGND VGND VPWR VPWR _10480_ sky130_fd_sc_hd__a31o_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28421_ clknet_leaf_20_clk _02219_ VGND VGND VPWR VPWR systolic_inst.A_shift\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25633_ systolic_inst.acc_wires\[3\]\[13\] C_out\[109\] net49 VGND VGND VPWR VPWR
+ _02935_ sky130_fd_sc_hd__mux2_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22845_ systolic_inst.A_outs\[1\]\[1\] systolic_inst.B_outs\[1\]\[7\] VGND VGND VPWR
+ VPWR _09526_ sky130_fd_sc_hd__and2b_1
XFILLER_77_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28352_ clknet_leaf_343_clk _02150_ VGND VGND VPWR VPWR systolic_inst.A_shift\[24\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25564_ systolic_inst.acc_wires\[1\]\[8\] C_out\[40\] net36 VGND VGND VPWR VPWR _02866_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_A_in_serial_clk clknet_2_3__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_17_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_22776_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[4\] _09457_ _09458_
+ VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__nand4_2
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27303_ clknet_leaf_288_clk _01101_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_24515_ C_out\[84\] net100 net82 ser_C.shift_reg\[84\] _10727_ VGND VGND VPWR VPWR
+ _02334_ sky130_fd_sc_hd__a221o_1
XFILLER_223_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21727_ _08532_ _08533_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__nand2b_1
X_28283_ clknet_leaf_48_clk _02081_ VGND VGND VPWR VPWR systolic_inst.B_shift\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25495_ _00008_ _11225_ VGND VGND VPWR VPWR _11227_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27234_ clknet_leaf_275_clk _01032_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24446_ net114 ser_C.shift_reg\[51\] VGND VGND VPWR VPWR _10693_ sky130_fd_sc_hd__and2_1
XFILLER_197_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21658_ _08412_ _08427_ _08426_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__o21a_1
XFILLER_40_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20609_ _07514_ _07518_ _07519_ _07538_ VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__a31o_1
X_27165_ clknet_leaf_273_clk _00963_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24377_ C_out\[15\] net104 _10643_ ser_C.shift_reg\[15\] _10658_ VGND VGND VPWR VPWR
+ _02265_ sky130_fd_sc_hd__a221o_1
X_21589_ _08372_ _08397_ _08398_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__nor3_1
X_26116_ deser_B.serial_word\[71\] deser_B.shift_reg\[71\] _00001_ VGND VGND VPWR
+ VPWR _03418_ sky130_fd_sc_hd__mux2_1
XFILLER_193_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_186_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14130_ systolic_inst.A_outs\[15\]\[6\] systolic_inst.A_outs\[14\]\[6\] net118 VGND
+ VGND VPWR VPWR _00952_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23328_ _09944_ _09955_ _09956_ VGND VGND VPWR VPWR _09957_ sky130_fd_sc_hd__or3_1
X_27096_ clknet_leaf_7_B_in_serial_clk _00894_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_186_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_207_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26047_ deser_B.serial_word\[2\] deser_B.shift_reg\[2\] net55 VGND VGND VPWR VPWR
+ _03349_ sky130_fd_sc_hd__mux2_1
X_14061_ deser_B.shift_reg\[95\] deser_B.shift_reg\[96\] net126 VGND VGND VPWR VPWR
+ _00887_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23259_ net109 systolic_inst.acc_wires\[1\]\[28\] net65 _09903_ VGND VGND VPWR VPWR
+ _01902_ sky130_fd_sc_hd__a22o_1
XFILLER_152_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_199_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17820_ systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[3\] VGND VGND VPWR
+ VPWR _05018_ sky130_fd_sc_hd__nand2_1
XFILLER_239_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27998_ clknet_leaf_152_clk _01796_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17751_ _04972_ _04973_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__nand2_1
XFILLER_43_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14963_ _12080_ _12083_ VGND VGND VPWR VPWR _12084_ sky130_fd_sc_hd__xnor2_1
X_26949_ clknet_leaf_3_A_in_serial_clk _00747_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[82\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_86_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_48_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16702_ _04023_ _04019_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__nand2b_1
XFILLER_207_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13914_ deser_A.serial_word\[75\] deser_A.shift_reg\[75\] net57 VGND VGND VPWR VPWR
+ _00740_ sky130_fd_sc_hd__mux2_1
X_29668_ clknet_leaf_27_B_in_serial_clk _03463_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_17682_ _04905_ _04910_ _04914_ net60 VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__a31o_1
XFILLER_48_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14894_ _12000_ _12016_ VGND VGND VPWR VPWR _12017_ sky130_fd_sc_hd__xnor2_1
X_19421_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[7\]\[3\]
+ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__or2_1
X_28619_ clknet_leaf_215_clk _02417_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16633_ _03937_ _03940_ _03956_ _03957_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__a211o_1
X_13845_ deser_A.serial_word\[6\] deser_A.shift_reg\[6\] net58 VGND VGND VPWR VPWR
+ _00671_ sky130_fd_sc_hd__mux2_1
X_29599_ clknet_leaf_18_B_in_serial_clk _03394_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19352_ _06409_ _06410_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__xnor2_1
X_16564_ systolic_inst.acc_wires\[12\]\[28\] systolic_inst.acc_wires\[12\]\[29\] systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__o21a_1
X_13776_ B_in\[83\] deser_B.word_buffer\[83\] net85 VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18303_ _05470_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__nand2_1
XFILLER_31_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15515_ _12510_ _12545_ _12544_ VGND VGND VPWR VPWR _12573_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_175_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19283_ _06343_ _06344_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__nand2_1
XFILLER_128_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16495_ _03845_ _03847_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__nand2_1
XFILLER_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18234_ _05412_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__inv_2
X_15446_ systolic_inst.A_outs\[13\]\[4\] _12469_ _12487_ _12486_ _12483_ VGND VGND
+ VPWR VPWR _12506_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_171_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18165_ _05262_ _05350_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__nand2_1
X_15377_ _12441_ _12439_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[1\]
+ net107 VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_17116_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[22\]
+ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__nand2_1
Xmax_cap103 net104 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_12
XFILLER_117_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14328_ _11503_ _11505_ VGND VGND VPWR VPWR _11513_ sky130_fd_sc_hd__nand2_1
Xmax_cap114 net7 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_12
XFILLER_209_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18096_ _05249_ _05252_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__nor2_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap125 deser_B.receiving VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_12
Xmax_cap147 net149 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_16
XFILLER_144_668 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17047_ _04331_ _04347_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__nor2_1
XFILLER_171_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14259_ _11406_ _11445_ VGND VGND VPWR VPWR _11446_ sky130_fd_sc_hd__xnor2_1
XFILLER_217_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18998_ net108 systolic_inst.acc_wires\[8\]\[29\] net66 _06089_ VGND VGND VPWR VPWR
+ _01455_ sky130_fd_sc_hd__a22o_1
XFILLER_79_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17949_ _05103_ _05106_ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__nor3_1
XFILLER_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_77_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_113_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20960_ _07822_ _07823_ _07825_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19619_ systolic_inst.A_outs\[6\]\[7\] systolic_inst.A_outs\[5\]\[7\] net120 VGND
+ VGND VPWR VPWR _01529_ sky130_fd_sc_hd__mux2_1
X_20891_ _07765_ _07766_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__and2b_1
XFILLER_242_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22630_ _09337_ _09339_ _09342_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__a21oi_2
XFILLER_241_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_234_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_234_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22561_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[2\]\[14\]
+ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__or2_1
XFILLER_107_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_230_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21512_ systolic_inst.A_outs\[3\]\[0\] systolic_inst.A_outs\[3\]\[1\] systolic_inst.B_outs\[3\]\[3\]
+ systolic_inst.B_outs\[3\]\[4\] VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__nand4_1
X_24300_ _10623_ systolic_inst.A_shift\[11\]\[5\] net71 VGND VGND VPWR VPWR _02223_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_230_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_230_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22492_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[2\]\[4\]
+ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__nand2_1
X_25280_ net111 ser_C.shift_reg\[468\] VGND VGND VPWR VPWR _11110_ sky130_fd_sc_hd__and2_1
XFILLER_221_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21443_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[28\]
+ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24231_ systolic_inst.A_shift\[20\]\[7\] A_in\[79\] net59 VGND VGND VPWR VPWR _10601_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24162_ _10582_ systolic_inst.A_shift\[27\]\[4\] net70 VGND VGND VPWR VPWR _02126_
+ sky130_fd_sc_hd__mux2_1
X_21374_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[18\]
+ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__or2_1
XFILLER_174_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23113_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[1\]\[7\]
+ VGND VGND VPWR VPWR _09779_ sky130_fd_sc_hd__nand2_1
X_20325_ systolic_inst.B_outs\[5\]\[3\] systolic_inst.A_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\]
+ systolic_inst.A_outs\[5\]\[2\] VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__a22o_1
X_28970_ clknet_leaf_56_clk _02768_ VGND VGND VPWR VPWR systolic_inst.B_shift\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24093_ systolic_inst.B_shift\[23\]\[2\] B_in\[58\] net59 VGND VGND VPWR VPWR _10556_
+ sky130_fd_sc_hd__mux2_1
XFILLER_235_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_181_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27921_ clknet_leaf_145_clk _01719_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_23044_ _09717_ _09718_ VGND VGND VPWR VPWR _09719_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_231_Right_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20256_ _07196_ _07197_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27852_ clknet_leaf_36_clk _01650_ net137 VGND VGND VPWR VPWR systolic_inst.A_outs\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_38_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20187_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[26\]
+ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__or2_1
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26803_ clknet_leaf_91_clk _00605_ net5 VGND VGND VPWR VPWR B_in\[75\] sky130_fd_sc_hd__dfrtp_1
XFILLER_118_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27783_ clknet_leaf_185_clk _01581_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_218_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24995_ C_out\[324\] net97 net80 ser_C.shift_reg\[324\] _10967_ VGND VGND VPWR VPWR
+ _02574_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_68_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
X_29522_ clknet_leaf_258_clk _03320_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[494\]
+ sky130_fd_sc_hd__dfrtp_1
X_26734_ clknet_leaf_96_clk _00536_ net153 VGND VGND VPWR VPWR B_in\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_91_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23946_ systolic_inst.B_shift\[14\]\[5\] B_in\[21\] net59 VGND VGND VPWR VPWR _10502_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29453_ clknet_leaf_289_clk _03251_ net136 VGND VGND VPWR VPWR C_out\[425\] sky130_fd_sc_hd__dfrtp_1
X_26665_ clknet_leaf_4_B_in_serial_clk _00468_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23877_ _10462_ _10465_ VGND VGND VPWR VPWR _10466_ sky130_fd_sc_hd__xor2_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28404_ clknet_leaf_88_clk _02202_ VGND VGND VPWR VPWR systolic_inst.B_shift\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25616_ systolic_inst.acc_wires\[2\]\[28\] C_out\[92\] net50 VGND VGND VPWR VPWR
+ _02918_ sky130_fd_sc_hd__mux2_1
XFILLER_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13630_ deser_B.word_buffer\[66\] deser_B.serial_word\[66\] net123 VGND VGND VPWR
+ VPWR _00467_ sky130_fd_sc_hd__mux2_1
X_22828_ _09444_ _09445_ _09475_ _09474_ VGND VGND VPWR VPWR _09510_ sky130_fd_sc_hd__a31o_1
X_29384_ clknet_leaf_245_clk _03182_ net145 VGND VGND VPWR VPWR C_out\[356\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26596_ clknet_leaf_0_A_in_serial_clk _00399_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28335_ clknet_leaf_343_clk _02133_ VGND VGND VPWR VPWR systolic_inst.A_shift\[26\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25547_ systolic_inst.acc_wires\[0\]\[23\] C_out\[23\] net53 VGND VGND VPWR VPWR
+ _02849_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13561_ deser_A.shift_reg\[125\] deser_A.shift_reg\[126\] net130 VGND VGND VPWR VPWR
+ _00398_ sky130_fd_sc_hd__mux2_1
X_22759_ _09411_ _09414_ _09441_ VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__nor3_1
XFILLER_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15300_ _11712_ _12390_ _12391_ systolic_inst.acc_wires\[14\]\[22\] net107 VGND VGND
+ VPWR VPWR _01064_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_188_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28266_ clknet_leaf_76_clk _02064_ VGND VGND VPWR VPWR systolic_inst.B_shift\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16280_ systolic_inst.B_outs\[12\]\[6\] systolic_inst.A_outs\[12\]\[6\] _11260_ systolic_inst.A_outs\[12\]\[5\]
+ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__o2bb2a_1
X_25478_ systolic_inst.ce_local _11215_ VGND VGND VPWR VPWR _11216_ sky130_fd_sc_hd__and2_1
XFILLER_212_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_188_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13492_ deser_A.shift_reg\[56\] deser_A.shift_reg\[57\] net130 VGND VGND VPWR VPWR
+ _00329_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15231_ _12329_ _12330_ VGND VGND VPWR VPWR _12333_ sky130_fd_sc_hd__nor2_1
X_27217_ clknet_leaf_292_clk _01015_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_24429_ C_out\[41\] _11302_ net81 ser_C.shift_reg\[41\] _10684_ VGND VGND VPWR VPWR
+ _02291_ sky130_fd_sc_hd__a221o_1
XFILLER_240_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28197_ clknet_leaf_48_clk _01995_ VGND VGND VPWR VPWR systolic_inst.B_shift\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15162_ _11712_ _12271_ _12273_ systolic_inst.acc_wires\[14\]\[2\] net107 VGND VGND
+ VPWR VPWR _01044_ sky130_fd_sc_hd__a32o_1
X_27148_ clknet_leaf_252_clk _00946_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14113_ systolic_inst.B_shift\[12\]\[5\] net72 _11333_ B_in\[101\] VGND VGND VPWR
+ VPWR _00935_ sky130_fd_sc_hd__a22o_1
XFILLER_125_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19970_ _06924_ _06965_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__xnor2_1
X_27079_ clknet_leaf_28_B_in_serial_clk _00877_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15093_ _12181_ _12209_ VGND VGND VPWR VPWR _12210_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14044_ deser_B.shift_reg\[78\] deser_B.shift_reg\[79\] deser_B.receiving VGND VGND
+ VPWR VPWR _00870_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18921_ net108 systolic_inst.acc_wires\[8\]\[17\] net66 _06024_ VGND VGND VPWR VPWR
+ _01443_ sky130_fd_sc_hd__a22o_1
XFILLER_141_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18852_ _05956_ _05960_ _05963_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__nand3_1
XFILLER_84_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17803_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.A_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\]
+ systolic_inst.A_outs\[9\]\[1\] VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__and4_1
X_18783_ _05904_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__nor2_1
X_15995_ _12982_ _12993_ VGND VGND VPWR VPWR _12994_ sky130_fd_sc_hd__or2_1
XFILLER_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_59_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_83_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17734_ _11712_ _04958_ _04959_ systolic_inst.acc_wires\[10\]\[23\] net105 VGND VGND
+ VPWR VPWR _01321_ sky130_fd_sc_hd__a32o_1
X_14946_ _12064_ _12065_ VGND VGND VPWR VPWR _12068_ sky130_fd_sc_hd__nand2b_1
XFILLER_48_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17665_ _04892_ _04893_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__a21o_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14877_ _11963_ _11999_ VGND VGND VPWR VPWR _12000_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19404_ net119 _06459_ _06460_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__a21oi_1
X_16616_ _03928_ _03930_ _03941_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__a21oi_1
X_13828_ deser_B.bit_idx\[2\] _11320_ _11321_ VGND VGND VPWR VPWR _11324_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17596_ _04838_ _04839_ _04840_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__and3_1
XFILLER_63_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19335_ _06394_ _06395_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__nor2_1
X_16547_ net108 systolic_inst.acc_wires\[12\]\[26\] net67 _03897_ VGND VGND VPWR VPWR
+ _01196_ sky130_fd_sc_hd__a22o_1
XFILLER_210_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13759_ B_in\[66\] deser_B.word_buffer\[66\] net87 VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19266_ _06328_ _06327_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__nand2b_1
X_16478_ _03825_ _03829_ _03835_ _03838_ _03830_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__o221a_1
XFILLER_148_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18217_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[9\]\[4\]
+ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__or2_1
X_15429_ systolic_inst.A_outs\[13\]\[2\] systolic_inst.B_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\]
+ systolic_inst.A_outs\[13\]\[1\] VGND VGND VPWR VPWR _12490_ sky130_fd_sc_hd__a22oi_1
XFILLER_191_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19197_ _06207_ _06222_ _06221_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__o21a_1
XFILLER_223_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18148_ _05291_ _05304_ _05302_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__o21a_1
XFILLER_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18079_ _05268_ _05267_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__nand2b_1
XFILLER_85_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20110_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[6\]\[13\]
+ _07083_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__a21oi_1
XFILLER_160_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21090_ systolic_inst.A_outs\[4\]\[5\] _07884_ _07960_ VGND VGND VPWR VPWR _07961_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_154_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20041_ _07026_ _07027_ _07028_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__and3_1
XFILLER_63_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23800_ _10399_ _10400_ VGND VGND VPWR VPWR _10401_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24780_ net113 ser_C.shift_reg\[218\] VGND VGND VPWR VPWR _10860_ sky130_fd_sc_hd__and2_1
XFILLER_27_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21992_ systolic_inst.acc_wires\[3\]\[16\] systolic_inst.acc_wires\[3\]\[17\] systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__o21ai_1
XFILLER_22_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_236_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_236_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_236_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23731_ _10335_ _10336_ _10334_ VGND VGND VPWR VPWR _10342_ sky130_fd_sc_hd__a21bo_1
X_20943_ _07816_ _07817_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__nor2_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_232_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26450_ clknet_leaf_10_clk _00257_ net132 VGND VGND VPWR VPWR A_in\[118\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_232_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _10280_ _10281_ VGND VGND VPWR VPWR _10282_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20874_ _07750_ VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__inv_2
XFILLER_109_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25401_ systolic_inst.A_shift\[2\]\[0\] A_in\[8\] net59 VGND VGND VPWR VPWR _11170_
+ sky130_fd_sc_hd__mux2_1
X_22613_ systolic_inst.acc_wires\[2\]\[20\] systolic_inst.acc_wires\[2\]\[21\] systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__o21a_1
X_26381_ clknet_leaf_20_clk _00188_ net133 VGND VGND VPWR VPWR A_in\[49\] sky130_fd_sc_hd__dfrtp_1
XFILLER_197_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23593_ _10173_ _10176_ _10213_ _10214_ VGND VGND VPWR VPWR _10215_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_42_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28120_ clknet_leaf_126_clk _01918_ net142 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_25332_ net112 ser_C.shift_reg\[494\] VGND VGND VPWR VPWR _11136_ sky130_fd_sc_hd__and2_1
X_22544_ net109 systolic_inst.acc_wires\[2\]\[11\] net65 _09269_ VGND VGND VPWR VPWR
+ _01821_ sky130_fd_sc_hd__a22o_1
XFILLER_167_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28051_ clknet_leaf_129_clk _01849_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_25263_ ser_C.parallel_data\[458\] net102 net74 ser_C.shift_reg\[458\] _11101_ VGND
+ VGND VPWR VPWR _02708_ sky130_fd_sc_hd__a221o_1
X_22475_ _09210_ VGND VGND VPWR VPWR _09211_ sky130_fd_sc_hd__inv_2
XFILLER_194_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27002_ clknet_leaf_15_B_in_serial_clk _00800_ net152 VGND VGND VPWR VPWR deser_B.shift_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24214_ _10592_ systolic_inst.A_shift\[20\]\[6\] net71 VGND VGND VPWR VPWR _02168_
+ sky130_fd_sc_hd__mux2_1
X_21426_ _08260_ _08262_ _08264_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25194_ net111 ser_C.shift_reg\[425\] VGND VGND VPWR VPWR _11067_ sky130_fd_sc_hd__and2_1
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21357_ _08204_ _08205_ _08198_ _08202_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__o211ai_1
X_24145_ systolic_inst.A_shift\[29\]\[4\] A_in\[108\] net59 VGND VGND VPWR VPWR _10574_
+ sky130_fd_sc_hd__mux2_1
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20308_ _07217_ _07220_ _07247_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__o21a_1
XFILLER_190_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24076_ systolic_inst.B_shift\[3\]\[3\] _11332_ net83 systolic_inst.B_shift\[7\]\[3\]
+ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__a22o_1
X_28953_ clknet_leaf_263_clk _02751_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[501\]
+ sky130_fd_sc_hd__dfrtp_1
X_21288_ _08147_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__inv_2
XFILLER_235_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23027_ _09700_ _09701_ VGND VGND VPWR VPWR _09703_ sky130_fd_sc_hd__and2b_1
X_27904_ clknet_leaf_43_clk _01702_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_20239_ net116 systolic_inst.B_outs\[5\]\[0\] systolic_inst.A_outs\[5\]\[0\] VGND
+ VGND VPWR VPWR _07184_ sky130_fd_sc_hd__and3_1
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28884_ clknet_leaf_328_clk _02682_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[432\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27835_ clknet_leaf_145_clk _01633_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14800_ _11918_ _11924_ VGND VGND VPWR VPWR _11926_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_177_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27766_ clknet_leaf_210_clk _01564_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_15780_ net66 _12823_ _12825_ systolic_inst.acc_wires\[13\]\[4\] net107 VGND VGND
+ VPWR VPWR _01110_ sky130_fd_sc_hd__a32o_1
XFILLER_218_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24978_ net111 ser_C.shift_reg\[317\] VGND VGND VPWR VPWR _10959_ sky130_fd_sc_hd__and2_1
XFILLER_188_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26717_ clknet_leaf_29_B_in_serial_clk _00520_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29505_ clknet_leaf_266_clk _03303_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[477\]
+ sky130_fd_sc_hd__dfrtp_1
X_14731_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[30\]
+ VGND VGND VPWR VPWR _11879_ sky130_fd_sc_hd__or2_1
XFILLER_218_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23929_ systolic_inst.A_shift\[3\]\[1\] net71 _11333_ A_in\[25\] VGND VGND VPWR VPWR
+ _01979_ sky130_fd_sc_hd__a22o_1
XFILLER_57_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27697_ clknet_leaf_196_clk _01495_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29436_ clknet_leaf_335_clk _03234_ net131 VGND VGND VPWR VPWR C_out\[408\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17450_ _04665_ _04703_ _04702_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__a21oi_2
X_26648_ clknet_leaf_20_B_in_serial_clk _00451_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_14662_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[20\]
+ VGND VGND VPWR VPWR _11820_ sky130_fd_sc_hd__nand2_1
XFILLER_232_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16401_ _03772_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__inv_2
X_13613_ deser_B.word_buffer\[49\] deser_B.serial_word\[49\] net124 VGND VGND VPWR
+ VPWR _00450_ sky130_fd_sc_hd__mux2_1
XFILLER_232_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29367_ clknet_leaf_201_clk _03165_ net147 VGND VGND VPWR VPWR C_out\[339\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17381_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[8\] _04637_ net118
+ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__mux2_1
XFILLER_214_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26579_ clknet_leaf_28_A_in_serial_clk _00382_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_14593_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[15\]\[10\]
+ VGND VGND VPWR VPWR _11761_ sky130_fd_sc_hd__or2_1
X_19120_ _06184_ _06185_ _06156_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16332_ _03681_ _03686_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__nor2_1
X_28318_ clknet_leaf_2_clk _02116_ VGND VGND VPWR VPWR systolic_inst.A_shift\[28\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13544_ deser_A.shift_reg\[108\] deser_A.shift_reg\[109\] net129 VGND VGND VPWR VPWR
+ _00381_ sky130_fd_sc_hd__mux2_1
XFILLER_242_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29298_ clknet_leaf_311_clk _03096_ net141 VGND VGND VPWR VPWR C_out\[270\] sky130_fd_sc_hd__dfrtp_1
XFILLER_203_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19051_ _06114_ _06119_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__xnor2_1
X_28249_ clknet_leaf_80_clk _02047_ VGND VGND VPWR VPWR systolic_inst.B_shift\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16263_ _03643_ _03644_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__nand2_1
XFILLER_125_1088 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13475_ deser_A.shift_reg\[39\] deser_A.shift_reg\[40\] net129 VGND VGND VPWR VPWR
+ _00312_ sky130_fd_sc_hd__mux2_1
XFILLER_201_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18002_ _05192_ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__nor2_1
X_15214_ _12311_ _12317_ VGND VGND VPWR VPWR _12318_ sky130_fd_sc_hd__nand2_1
XFILLER_195_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16194_ _03536_ _03537_ _03539_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__o21a_1
XFILLER_51_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_19_B_in_serial_clk clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_19_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_15145_ _12259_ _12252_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ net107 VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_142_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19953_ _06946_ _06948_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_112_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15076_ _12191_ _12192_ VGND VGND VPWR VPWR _12194_ sky130_fd_sc_hd__and2b_1
X_14027_ deser_B.shift_reg\[61\] deser_B.shift_reg\[62\] net126 VGND VGND VPWR VPWR
+ _00853_ sky130_fd_sc_hd__mux2_1
X_18904_ _06007_ _06008_ _06001_ _06005_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__o211ai_1
XFILLER_84_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19884_ _06881_ _06882_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__or2_1
XFILLER_67_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18835_ _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__inv_2
XFILLER_132_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15978_ systolic_inst.A_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[1\]
+ systolic_inst.B_outs\[12\]\[0\] VGND VGND VPWR VPWR _12979_ sky130_fd_sc_hd__a22o_1
X_18766_ _05856_ _05861_ _05888_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_121_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17717_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[21\]
+ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__xnor2_2
XFILLER_48_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14929_ _11976_ _12010_ _12012_ VGND VGND VPWR VPWR _12051_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18697_ _05820_ _05821_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_82_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17648_ _04884_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__nand2_1
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17579_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[10\]\[1\]
+ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__nand2_1
XFILLER_225_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19318_ _06377_ _06378_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__nor2_1
XFILLER_182_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20590_ net109 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[14\] VGND
+ VGND VPWR VPWR _07521_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_119_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19249_ _06277_ _06311_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__xor2_1
XFILLER_143_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22260_ _08929_ _08964_ _08966_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__a21oi_2
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21211_ _08077_ _08078_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_22_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22191_ _08935_ _08936_ _08906_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_225_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21142_ _07962_ _07970_ _07969_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__a21o_1
XFILLER_133_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25950_ systolic_inst.acc_wires\[13\]\[10\] C_out\[426\] net19 VGND VGND VPWR VPWR
+ _03252_ sky130_fd_sc_hd__mux2_1
X_21073_ _07913_ _07944_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20024_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[6\]\[2\]
+ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__or2_1
X_24901_ C_out\[277\] net103 net75 ser_C.shift_reg\[277\] _10920_ VGND VGND VPWR VPWR
+ _02527_ sky130_fd_sc_hd__a221o_1
XFILLER_28_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_238_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25881_ systolic_inst.acc_wires\[11\]\[5\] C_out\[357\] net38 VGND VGND VPWR VPWR
+ _03183_ sky130_fd_sc_hd__mux2_1
XFILLER_100_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27620_ clknet_leaf_318_clk _01418_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24832_ net113 ser_C.shift_reg\[244\] VGND VGND VPWR VPWR _10886_ sky130_fd_sc_hd__and2_1
XFILLER_58_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27551_ clknet_leaf_299_clk _01349_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_24763_ C_out\[208\] net99 net79 ser_C.shift_reg\[208\] _10851_ VGND VGND VPWR VPWR
+ _02458_ sky130_fd_sc_hd__a221o_1
X_21975_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[3\]\[12\]
+ _08741_ _08743_ VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__a31o_1
XFILLER_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26502_ clknet_leaf_15_A_in_serial_clk _00305_ net137 VGND VGND VPWR VPWR deser_A.shift_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_23714_ net63 _10325_ _10327_ systolic_inst.acc_wires\[0\]\[3\] _11258_ VGND VGND
+ VPWR VPWR _01933_ sky130_fd_sc_hd__a32o_1
X_27482_ clknet_leaf_41_clk _01280_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_20926_ _07759_ _07776_ _07778_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__o21a_1
X_24694_ net112 ser_C.shift_reg\[175\] VGND VGND VPWR VPWR _10817_ sky130_fd_sc_hd__and2_1
XFILLER_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29221_ clknet_leaf_208_clk _03019_ net147 VGND VGND VPWR VPWR C_out\[193\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26433_ clknet_leaf_0_clk _00240_ net134 VGND VGND VPWR VPWR A_in\[101\] sky130_fd_sc_hd__dfrtp_1
X_23645_ _10262_ _10264_ VGND VGND VPWR VPWR _10265_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20857_ net108 _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__nor2_1
XFILLER_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29152_ clknet_leaf_172_clk _02950_ net148 VGND VGND VPWR VPWR C_out\[124\] sky130_fd_sc_hd__dfrtp_1
X_26364_ clknet_leaf_24_clk _00171_ net135 VGND VGND VPWR VPWR A_in\[32\] sky130_fd_sc_hd__dfrtp_1
XFILLER_161_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23576_ _11267_ systolic_inst.B_outs\[0\]\[7\] _10120_ VGND VGND VPWR VPWR _10198_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_214_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20788_ _07687_ _07689_ _07691_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__or3_1
XFILLER_167_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28103_ clknet_leaf_111_clk _01901_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25315_ ser_C.parallel_data\[484\] net97 net77 ser_C.shift_reg\[484\] _11127_ VGND
+ VGND VPWR VPWR _02734_ sky130_fd_sc_hd__a221o_1
X_29083_ clknet_leaf_110_clk _02881_ net151 VGND VGND VPWR VPWR C_out\[55\] sky130_fd_sc_hd__dfrtp_1
X_22527_ _09250_ _09252_ VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__nand2_1
XFILLER_211_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26295_ clknet_leaf_27_A_in_serial_clk _00103_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28034_ clknet_leaf_158_clk _01832_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_210_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25246_ net111 ser_C.shift_reg\[451\] VGND VGND VPWR VPWR _11093_ sky130_fd_sc_hd__and2_1
X_13260_ deser_A.word_buffer\[98\] deser_A.serial_word\[98\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22458_ _09148_ _09152_ _09174_ _09175_ VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__o31a_1
XFILLER_196_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21409_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[23\]
+ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__xor2_1
XFILLER_124_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13191_ deser_A.word_buffer\[29\] deser_A.serial_word\[29\] net128 VGND VGND VPWR
+ VPWR _00039_ sky130_fd_sc_hd__mux2_1
X_25177_ C_out\[415\] net101 net73 ser_C.shift_reg\[415\] _11058_ VGND VGND VPWR VPWR
+ _02665_ sky130_fd_sc_hd__a221o_1
X_22389_ systolic_inst.B_outs\[2\]\[5\] systolic_inst.A_outs\[2\]\[7\] VGND VGND VPWR
+ VPWR _09130_ sky130_fd_sc_hd__nand2_1
XFILLER_159_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24128_ _10565_ systolic_inst.A_shift\[29\]\[3\] net71 VGND VGND VPWR VPWR _02109_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24059_ systolic_inst.B_shift\[19\]\[1\] B_in\[25\] net59 VGND VGND VPWR VPWR _10547_
+ sky130_fd_sc_hd__mux2_1
X_28936_ clknet_leaf_260_clk _02734_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[484\]
+ sky130_fd_sc_hd__dfrtp_1
X_16950_ _04264_ _04263_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__and2b_1
XFILLER_238_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15901_ _12927_ _12928_ _12926_ VGND VGND VPWR VPWR _12929_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16881_ _04056_ _04196_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__nand2_2
X_28867_ clknet_leaf_333_clk _02665_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[415\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15832_ _12867_ _12868_ _12869_ VGND VGND VPWR VPWR _12870_ sky130_fd_sc_hd__and3_1
X_18620_ _05739_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__xnor2_1
X_27818_ clknet_leaf_143_clk _01616_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_28798_ clknet_leaf_236_clk _02596_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[346\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_204_Left_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15763_ _12808_ _12809_ _12810_ VGND VGND VPWR VPWR _12811_ sky130_fd_sc_hd__a21o_1
X_18551_ _05664_ _05680_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27749_ clknet_leaf_209_clk _01547_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14714_ _11857_ _11861_ VGND VGND VPWR VPWR _11864_ sky130_fd_sc_hd__nor2_1
X_17502_ _04753_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__nand2_1
X_18482_ _05612_ _05613_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__or2_1
XFILLER_73_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ systolic_inst.A_outs\[13\]\[6\] _11272_ VGND VGND VPWR VPWR _12747_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_159_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _04678_ _04686_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__or2_1
X_14645_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[17\]
+ VGND VGND VPWR VPWR _11806_ sky130_fd_sc_hd__xor2_2
X_29419_ clknet_leaf_333_clk _03217_ net131 VGND VGND VPWR VPWR C_out\[391\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17364_ _04611_ _04619_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__xnor2_1
X_14576_ _11740_ _11741_ _11739_ VGND VGND VPWR VPWR _11747_ sky130_fd_sc_hd__a21bo_1
XFILLER_60_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19103_ systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[5\] systolic_inst.A_outs\[7\]\[6\]
+ systolic_inst.B_outs\[7\]\[0\] VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__a22oi_1
XFILLER_14_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16315_ _03662_ _03665_ _03693_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__or3_1
XFILLER_174_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13527_ deser_A.shift_reg\[91\] deser_A.shift_reg\[92\] net129 VGND VGND VPWR VPWR
+ _00364_ sky130_fd_sc_hd__mux2_1
X_17295_ _04530_ _04552_ _04553_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__and3_1
XFILLER_201_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19034_ systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[2\]
+ systolic_inst.B_outs\[7\]\[0\] VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__a22oi_1
XPHY_EDGE_ROW_213_Left_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16246_ _03517_ _03626_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_168_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13458_ deser_A.shift_reg\[22\] deser_A.shift_reg\[23\] deser_A.receiving VGND VGND
+ VPWR VPWR _00295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16177_ systolic_inst.B_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[5\] systolic_inst.A_outs\[12\]\[6\]
+ systolic_inst.B_outs\[12\]\[3\] VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_110_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13389_ A_in\[98\] deser_A.word_buffer\[98\] net96 VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15128_ _12241_ _12242_ VGND VGND VPWR VPWR _12244_ sky130_fd_sc_hd__and2b_1
XFILLER_217_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_290_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_290_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19936_ _06895_ _06932_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15059_ _12176_ VGND VGND VPWR VPWR _12177_ sky130_fd_sc_hd__inv_2
XFILLER_25_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19867_ _06830_ _06832_ _06831_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_222_Left_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18818_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[8\]\[3\]
+ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19798_ _06798_ _06797_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__nand2b_1
XFILLER_7_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18749_ _05806_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__nand2_1
XFILLER_97_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21760_ _08556_ _08564_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_218_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20711_ _07622_ _07624_ _07626_ systolic_inst.acc_wires\[5\]\[13\] net109 VGND VGND
+ VPWR VPWR _01631_ sky130_fd_sc_hd__a32o_1
XFILLER_93_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21691_ _08459_ _08461_ _08498_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__a21o_1
XFILLER_180_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23430_ _09993_ _09996_ _10054_ _10055_ VGND VGND VPWR VPWR _10056_ sky130_fd_sc_hd__a211oi_4
X_20642_ net63 _07566_ _07567_ systolic_inst.acc_wires\[5\]\[3\] net107 VGND VGND
+ VPWR VPWR _01621_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_24_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_231_Left_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23361_ _09959_ _09987_ VGND VGND VPWR VPWR _09989_ sky130_fd_sc_hd__xor2_1
XFILLER_165_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20573_ _07435_ _07474_ _07473_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__a21bo_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_227_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25100_ net113 ser_C.shift_reg\[378\] VGND VGND VPWR VPWR _11020_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_227_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22312_ _09025_ _09026_ _09027_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__o21ba_1
XFILLER_178_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26080_ deser_B.serial_word\[35\] deser_B.shift_reg\[35\] net55 VGND VGND VPWR VPWR
+ _03382_ sky130_fd_sc_hd__mux2_1
X_23292_ systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[1\] systolic_inst.A_outs\[0\]\[1\]
+ systolic_inst.B_outs\[0\]\[2\] VGND VGND VPWR VPWR _09923_ sky130_fd_sc_hd__nand4_2
XFILLER_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25031_ C_out\[342\] net97 net77 ser_C.shift_reg\[342\] _10985_ VGND VGND VPWR VPWR
+ _02592_ sky130_fd_sc_hd__a221o_1
X_22243_ _08983_ _08986_ VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22174_ _08916_ _08919_ VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_281_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_281_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21125_ _07955_ _07994_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__or2_1
XFILLER_132_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26982_ clknet_leaf_29_A_in_serial_clk _00780_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_240_Left_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21056_ systolic_inst.A_outs\[4\]\[2\] _11271_ _07850_ VGND VGND VPWR VPWR _07928_
+ sky130_fd_sc_hd__o21ai_1
X_25933_ systolic_inst.acc_wires\[12\]\[25\] C_out\[409\] net21 VGND VGND VPWR VPWR
+ _03235_ sky130_fd_sc_hd__mux2_1
X_28721_ clknet_leaf_310_clk _02519_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20007_ _06924_ _06986_ _06984_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__a21oi_1
X_28652_ clknet_leaf_203_clk _02450_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[200\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_115_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25864_ systolic_inst.acc_wires\[10\]\[20\] C_out\[340\] net11 VGND VGND VPWR VPWR
+ _03166_ sky130_fd_sc_hd__mux2_1
XFILLER_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_203_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24815_ C_out\[234\] net99 net79 ser_C.shift_reg\[234\] _10877_ VGND VGND VPWR VPWR
+ _02484_ sky130_fd_sc_hd__a221o_1
X_27603_ clknet_leaf_33_clk _01401_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_234_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28583_ clknet_leaf_309_clk _02381_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[131\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25795_ systolic_inst.acc_wires\[8\]\[15\] C_out\[271\] net28 VGND VGND VPWR VPWR
+ _03097_ sky130_fd_sc_hd__mux2_1
XFILLER_234_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27534_ clknet_leaf_312_clk _01332_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_195_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24746_ net112 ser_C.shift_reg\[201\] VGND VGND VPWR VPWR _10843_ sky130_fd_sc_hd__and2_1
XFILLER_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21958_ _08737_ _08740_ _08744_ VGND VGND VPWR VPWR _08746_ sky130_fd_sc_hd__a21o_1
XFILLER_242_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27465_ clknet_leaf_237_clk _01263_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_20909_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[5\] _07782_ _07783_
+ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__a22o_1
X_24677_ C_out\[165\] net103 net76 ser_C.shift_reg\[165\] _10808_ VGND VGND VPWR VPWR
+ _02415_ sky130_fd_sc_hd__a221o_1
X_21889_ _08686_ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__inv_2
XFILLER_163_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_212_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29204_ clknet_leaf_206_clk _03002_ net147 VGND VGND VPWR VPWR C_out\[176\] sky130_fd_sc_hd__dfrtp_1
X_14430_ _11575_ _11578_ _11612_ VGND VGND VPWR VPWR _11613_ sky130_fd_sc_hd__a21oi_1
X_26416_ clknet_leaf_5_clk _00223_ net133 VGND VGND VPWR VPWR A_in\[84\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_212_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628_ _10211_ _10213_ VGND VGND VPWR VPWR _10249_ sky130_fd_sc_hd__or2_1
XFILLER_39_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27396_ clknet_leaf_335_clk _01194_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29135_ clknet_leaf_168_clk _02933_ net148 VGND VGND VPWR VPWR C_out\[107\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26347_ clknet_leaf_20_clk _00154_ net135 VGND VGND VPWR VPWR A_in\[15\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _11545_ _11513_ VGND VGND VPWR VPWR _11546_ sky130_fd_sc_hd__and2b_1
XFILLER_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23559_ _10178_ _10179_ _10180_ VGND VGND VPWR VPWR _10182_ sky130_fd_sc_hd__nor3b_1
XFILLER_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16100_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[5\] VGND VGND
+ VPWR VPWR _13095_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ A_in\[21\] deser_A.word_buffer\[21\] net92 VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__mux2_1
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29066_ clknet_leaf_115_clk _02864_ net152 VGND VGND VPWR VPWR C_out\[38\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17080_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[16\]
+ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14292_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[6\]
+ systolic_inst.A_outs\[15\]\[7\] VGND VGND VPWR VPWR _11478_ sky130_fd_sc_hd__and4_1
X_26278_ clknet_leaf_20_A_in_serial_clk _00086_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28017_ clknet_leaf_154_clk _01815_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16031_ systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[5\]
+ systolic_inst.B_outs\[12\]\[0\] VGND VGND VPWR VPWR _13028_ sky130_fd_sc_hd__a22oi_1
X_25229_ ser_C.parallel_data\[441\] net102 net74 ser_C.shift_reg\[441\] _11084_ VGND
+ VGND VPWR VPWR _02691_ sky130_fd_sc_hd__a221o_1
X_13243_ deser_A.word_buffer\[81\] deser_A.serial_word\[81\] net127 VGND VGND VPWR
+ VPWR _00091_ sky130_fd_sc_hd__mux2_1
XFILLER_183_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13174_ deser_A.word_buffer\[12\] deser_A.serial_word\[12\] net127 VGND VGND VPWR
+ VPWR _00022_ sky130_fd_sc_hd__mux2_1
XFILLER_151_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_272_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_272_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_176_Right_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17982_ _05174_ _05173_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__nand2b_1
XFILLER_238_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19721_ _06720_ _06723_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28919_ clknet_leaf_269_clk _02717_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[467\]
+ sky130_fd_sc_hd__dfrtp_1
X_16933_ _04215_ _04218_ _04247_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__o21ai_1
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19652_ _06656_ _06657_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__nand2_1
XFILLER_38_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16864_ _04180_ _04181_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__nand2_1
XFILLER_203_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18603_ _05701_ _05703_ _05700_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__o21ba_1
XFILLER_168_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15815_ _12853_ _12854_ VGND VGND VPWR VPWR _12855_ sky130_fd_sc_hd__and2_1
XFILLER_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19583_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[27\]
+ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16795_ _04112_ _04113_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__xor2_1
XFILLER_206_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15746_ _12795_ _12796_ VGND VGND VPWR VPWR _12797_ sky130_fd_sc_hd__xnor2_1
X_18534_ _05628_ _05663_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_103_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_783 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15677_ _12684_ _12700_ _12698_ VGND VGND VPWR VPWR _12731_ sky130_fd_sc_hd__o21a_1
X_18465_ _05596_ _05597_ _05579_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__a21oi_1
XFILLER_209_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14628_ _11788_ _11791_ VGND VGND VPWR VPWR _11792_ sky130_fd_sc_hd__nand2_1
X_17416_ _04643_ _04644_ _04645_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__o21ba_1
X_18396_ _05547_ _05550_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17347_ _04603_ _04600_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__and2b_1
XFILLER_187_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14559_ net69 _11730_ _11732_ systolic_inst.acc_wires\[15\]\[4\] net107 VGND VGND
+ VPWR VPWR _00982_ sky130_fd_sc_hd__a32o_1
XFILLER_174_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload201 clknet_leaf_69_clk VGND VGND VPWR VPWR clkload201/Y sky130_fd_sc_hd__clkinvlp_4
X_17278_ _04507_ _04536_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__xor2_1
Xclkload212 clknet_leaf_46_clk VGND VGND VPWR VPWR clkload212/Y sky130_fd_sc_hd__inv_8
Xclkload223 clknet_leaf_129_clk VGND VGND VPWR VPWR clkload223/Y sky130_fd_sc_hd__bufinv_16
Xclkload234 clknet_leaf_85_clk VGND VGND VPWR VPWR clkload234/Y sky130_fd_sc_hd__clkinv_2
X_19017_ systolic_inst.A_outs\[7\]\[6\] systolic_inst.A_outs\[6\]\[6\] net119 VGND
+ VGND VPWR VPWR _01464_ sky130_fd_sc_hd__mux2_1
X_16229_ _03559_ _03576_ _03574_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__o21a_1
Xclkload245 clknet_leaf_121_clk VGND VGND VPWR VPWR clkload245/X sky130_fd_sc_hd__clkbuf_4
XFILLER_220_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload256 clknet_leaf_99_clk VGND VGND VPWR VPWR clkload256/Y sky130_fd_sc_hd__bufinv_16
XFILLER_162_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload267 clknet_leaf_137_clk VGND VGND VPWR VPWR clkload267/Y sky130_fd_sc_hd__inv_6
Xclkload278 clknet_leaf_147_clk VGND VGND VPWR VPWR clkload278/Y sky130_fd_sc_hd__clkinv_2
Xclkload289 clknet_leaf_193_clk VGND VGND VPWR VPWR clkload289/Y sky130_fd_sc_hd__inv_6
XFILLER_177_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_263_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_263_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19919_ _06914_ _06915_ _06883_ _06888_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__o211a_1
XFILLER_190_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22930_ _09608_ _09607_ VGND VGND VPWR VPWR _09609_ sky130_fd_sc_hd__nand2b_1
XFILLER_112_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_A_in_serial_clk clknet_2_1__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_25_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22861_ _09539_ _09540_ VGND VGND VPWR VPWR _09542_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_216_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24600_ net110 ser_C.shift_reg\[128\] VGND VGND VPWR VPWR _10770_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_216_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21812_ systolic_inst.A_outs\[3\]\[6\] _11274_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__nor2_1
X_25580_ systolic_inst.acc_wires\[1\]\[24\] C_out\[56\] net53 VGND VGND VPWR VPWR
+ _02882_ sky130_fd_sc_hd__mux2_1
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22792_ _09472_ _09473_ _09440_ _09442_ VGND VGND VPWR VPWR _09475_ sky130_fd_sc_hd__a211o_1
XFILLER_227_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24531_ C_out\[92\] net100 net82 ser_C.shift_reg\[92\] _10735_ VGND VGND VPWR VPWR
+ _02342_ sky130_fd_sc_hd__a221o_1
X_21743_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[10\] _08547_
+ _08549_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__a22o_1
XFILLER_149_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1055 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27250_ clknet_leaf_275_clk _01048_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24462_ net114 ser_C.shift_reg\[59\] VGND VGND VPWR VPWR _10701_ sky130_fd_sc_hd__and2_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21674_ _08443_ _08481_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__nor2_1
XFILLER_75_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26201_ systolic_inst.A_shift\[30\]\[7\] net71 _11333_ A_in\[127\] VGND VGND VPWR
+ VPWR _03491_ sky130_fd_sc_hd__a22o_1
X_23413_ systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[7\] VGND VGND VPWR
+ VPWR _10039_ sky130_fd_sc_hd__and2b_1
XFILLER_138_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20625_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[5\]\[0\]
+ _07551_ _07552_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__and4_1
X_27181_ clknet_leaf_273_clk _00979_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24393_ C_out\[23\] net104 _10643_ ser_C.shift_reg\[23\] _10666_ VGND VGND VPWR VPWR
+ _02273_ sky130_fd_sc_hd__a221o_1
XFILLER_165_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26132_ deser_B.serial_word\[87\] deser_B.shift_reg\[87\] net56 VGND VGND VPWR VPWR
+ _03434_ sky130_fd_sc_hd__mux2_1
XFILLER_193_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23344_ systolic_inst.A_outs\[0\]\[1\] systolic_inst.A_outs\[0\]\[2\] systolic_inst.B_outs\[0\]\[3\]
+ systolic_inst.B_outs\[0\]\[4\] VGND VGND VPWR VPWR _09972_ sky130_fd_sc_hd__and4_1
X_20556_ _07487_ _07488_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__or2_1
XFILLER_180_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26063_ deser_B.serial_word\[18\] deser_B.shift_reg\[18\] net55 VGND VGND VPWR VPWR
+ _03365_ sky130_fd_sc_hd__mux2_1
X_23275_ _09910_ _09914_ _09915_ _11713_ VGND VGND VPWR VPWR _09917_ sky130_fd_sc_hd__a31o_1
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20487_ _07420_ _07421_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__or2_2
XFILLER_180_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25014_ net111 ser_C.shift_reg\[335\] VGND VGND VPWR VPWR _10977_ sky130_fd_sc_hd__and2_1
X_22226_ _08933_ _08935_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__and2b_1
XFILLER_152_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_254_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_254_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_56_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22157_ _08903_ _08904_ VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__or2_1
XFILLER_105_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_205_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21108_ _07952_ _07978_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__nand2_1
XFILLER_120_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22088_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.B_shift\[1\]\[2\] net122 VGND
+ VGND VPWR VPWR _01788_ sky130_fd_sc_hd__mux2_1
X_26965_ clknet_leaf_23_A_in_serial_clk _00763_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_219_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28704_ clknet_leaf_187_clk _02502_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[252\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13930_ deser_A.serial_word\[91\] deser_A.shift_reg\[91\] net57 VGND VGND VPWR VPWR
+ _00756_ sky130_fd_sc_hd__mux2_1
XFILLER_102_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25916_ systolic_inst.acc_wires\[12\]\[8\] C_out\[392\] net18 VGND VGND VPWR VPWR
+ _03218_ sky130_fd_sc_hd__mux2_1
XFILLER_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21039_ _07910_ _07911_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__nor2_1
X_29684_ clknet_leaf_105_clk _03479_ net152 VGND VGND VPWR VPWR ser_C.bit_idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_197_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26896_ clknet_leaf_6_A_in_serial_clk _00694_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_197_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28635_ clknet_leaf_181_clk _02433_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[183\]
+ sky130_fd_sc_hd__dfrtp_1
X_13861_ deser_A.serial_word\[22\] deser_A.shift_reg\[22\] net58 VGND VGND VPWR VPWR
+ _00687_ sky130_fd_sc_hd__mux2_1
XFILLER_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25847_ systolic_inst.acc_wires\[10\]\[3\] C_out\[323\] net14 VGND VGND VPWR VPWR
+ _03149_ sky130_fd_sc_hd__mux2_1
XFILLER_35_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15600_ _12621_ _12623_ _12622_ VGND VGND VPWR VPWR _12656_ sky130_fd_sc_hd__o21ba_1
XFILLER_62_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16580_ systolic_inst.A_outs\[11\]\[5\] systolic_inst.A_outs\[10\]\[5\] net118 VGND
+ VGND VPWR VPWR _01207_ sky130_fd_sc_hd__mux2_1
X_28566_ clknet_leaf_165_clk _02364_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_13792_ B_in\[99\] deser_B.word_buffer\[99\] _00005_ VGND VGND VPWR VPWR _00629_
+ sky130_fd_sc_hd__mux2_1
X_25778_ systolic_inst.acc_wires\[7\]\[30\] C_out\[254\] net43 VGND VGND VPWR VPWR
+ _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_222_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15531_ systolic_inst.A_outs\[13\]\[1\] _11272_ systolic_inst.B_outs\[13\]\[6\] systolic_inst.A_outs\[13\]\[2\]
+ VGND VGND VPWR VPWR _12589_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_203_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24729_ C_out\[191\] net99 net79 ser_C.shift_reg\[191\] _10834_ VGND VGND VPWR VPWR
+ _02441_ sky130_fd_sc_hd__a221o_1
X_27517_ clknet_leaf_212_clk _01315_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28497_ clknet_leaf_117_clk _02295_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _05419_ _05422_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__nand2_1
X_15462_ _12519_ _12521_ VGND VGND VPWR VPWR _12522_ sky130_fd_sc_hd__nor2_1
XFILLER_76_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27448_ clknet_leaf_241_clk _01246_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_188_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17201_ systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[1\] VGND VGND
+ VPWR VPWR _04464_ sky130_fd_sc_hd__nand2_1
XFILLER_141_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14413_ systolic_inst.A_outs\[15\]\[5\] systolic_inst.B_outs\[15\]\[6\] _11273_ systolic_inst.A_outs\[15\]\[4\]
+ VGND VGND VPWR VPWR _11596_ sky130_fd_sc_hd__o2bb2a_1
X_18181_ _05342_ _05365_ _05366_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__or4_1
XFILLER_230_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27379_ clknet_leaf_340_clk _01177_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15393_ _12453_ _12454_ _12444_ VGND VGND VPWR VPWR _12456_ sky130_fd_sc_hd__a21o_1
XFILLER_141_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17132_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[24\]
+ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__nor2_1
X_29118_ clknet_leaf_163_clk _02916_ net151 VGND VGND VPWR VPWR C_out\[90\] sky130_fd_sc_hd__dfrtp_1
XFILLER_129_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14344_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[7\] VGND VGND
+ VPWR VPWR _11529_ sky130_fd_sc_hd__and2b_1
XFILLER_195_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_146_Left_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29049_ clknet_leaf_103_clk _02847_ net151 VGND VGND VPWR VPWR C_out\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_116_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17063_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[11\]\[14\]
+ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__nand2_1
XFILLER_128_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14275_ _11419_ _11460_ VGND VGND VPWR VPWR _11462_ sky130_fd_sc_hd__and2_1
XFILLER_195_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16014_ _12993_ _13010_ _13011_ VGND VGND VPWR VPWR _13012_ sky130_fd_sc_hd__a21oi_1
X_13226_ deser_A.word_buffer\[64\] deser_A.serial_word\[64\] net127 VGND VGND VPWR
+ VPWR _00074_ sky130_fd_sc_hd__mux2_1
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_245_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_245_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13157_ net56 _11305_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__nor2_1
XFILLER_124_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17965_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[6\] VGND VGND VPWR
+ VPWR _05158_ sky130_fd_sc_hd__nand2_1
XFILLER_239_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19704_ _06684_ _06706_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__xnor2_1
XFILLER_239_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16916_ _04204_ _04231_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__xnor2_1
XFILLER_214_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_155_Left_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17896_ _05087_ _05090_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19635_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.A_outs\[6\]\[2\] VGND VGND VPWR
+ VPWR _06642_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16847_ _04057_ _04163_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__nand2_1
XFILLER_19_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19566_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[24\]
+ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__nor2_1
XFILLER_92_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16778_ systolic_inst.B_outs\[11\]\[4\] systolic_inst.A_outs\[11\]\[5\] systolic_inst.A_outs\[11\]\[6\]
+ systolic_inst.B_outs\[11\]\[3\] VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__a22oi_1
XFILLER_225_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18517_ _05645_ _05646_ _05615_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__a21o_1
XFILLER_94_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15729_ _12715_ _12780_ VGND VGND VPWR VPWR _12781_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19497_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[7\]\[14\]
+ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18448_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[2\] VGND VGND VPWR
+ VPWR _05581_ sky130_fd_sc_hd__and2_1
XFILLER_179_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18379_ _05520_ _05522_ _05534_ _05535_ _05528_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__a311oi_4
XFILLER_144_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20410_ _07270_ _07305_ _07307_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_135_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_212_Right_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21390_ _08223_ _08228_ _08234_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__or3b_1
XFILLER_179_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20341_ _07277_ _07278_ _07254_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__a21o_1
XFILLER_31_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23060_ net122 _09733_ _09734_ _09713_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__a31o_1
X_20272_ _07209_ _07212_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22011_ _08790_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__inv_2
XFILLER_118_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_236_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_236_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_241_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_241_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26750_ clknet_leaf_56_clk _00552_ net143 VGND VGND VPWR VPWR B_in\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23962_ _10506_ systolic_inst.B_shift\[9\]\[0\] _11332_ VGND VGND VPWR VPWR _02002_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25701_ systolic_inst.acc_wires\[5\]\[17\] C_out\[177\] net47 VGND VGND VPWR VPWR
+ _03003_ sky130_fd_sc_hd__mux2_1
X_22913_ _09557_ _09591_ VGND VGND VPWR VPWR _09592_ sky130_fd_sc_hd__xor2_1
XFILLER_112_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26681_ clknet_leaf_26_B_in_serial_clk _00484_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_151_1095 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23893_ _10473_ _10477_ _10478_ VGND VGND VPWR VPWR _10479_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25632_ systolic_inst.acc_wires\[3\]\[12\] C_out\[108\] net49 VGND VGND VPWR VPWR
+ _02934_ sky130_fd_sc_hd__mux2_1
XFILLER_83_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28420_ clknet_leaf_20_clk _02218_ VGND VGND VPWR VPWR systolic_inst.A_shift\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_22844_ _09524_ VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__inv_2
XFILLER_72_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28351_ clknet_leaf_342_clk _02149_ VGND VGND VPWR VPWR systolic_inst.A_shift\[24\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25563_ systolic_inst.acc_wires\[1\]\[7\] C_out\[39\] net36 VGND VGND VPWR VPWR _02865_
+ sky130_fd_sc_hd__mux2_1
XFILLER_227_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22775_ systolic_inst.B_outs\[1\]\[3\] systolic_inst.A_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\]
+ systolic_inst.A_outs\[1\]\[2\] VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27302_ clknet_leaf_288_clk _01100_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24514_ net114 ser_C.shift_reg\[85\] VGND VGND VPWR VPWR _10727_ sky130_fd_sc_hd__and2_1
XFILLER_12_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21726_ _08489_ _08497_ _08496_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__a21bo_1
X_28282_ clknet_leaf_134_clk _02080_ VGND VGND VPWR VPWR systolic_inst.B_shift\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25494_ _11225_ _11226_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__nor2_1
X_27233_ clknet_leaf_275_clk _01031_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24445_ C_out\[49\] _11302_ net81 ser_C.shift_reg\[49\] _10692_ VGND VGND VPWR VPWR
+ _02299_ sky130_fd_sc_hd__a221o_1
XFILLER_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21657_ _08447_ _08464_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__xor2_1
XFILLER_36_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20608_ _07514_ _07518_ _07519_ _07538_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__nand4_1
X_27164_ clknet_leaf_273_clk _00962_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24376_ net7 ser_C.shift_reg\[16\] VGND VGND VPWR VPWR _10658_ sky130_fd_sc_hd__and2_1
X_21588_ _08397_ _08398_ _08372_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__o21ai_1
XFILLER_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26115_ deser_B.serial_word\[70\] deser_B.shift_reg\[70\] _00001_ VGND VGND VPWR
+ VPWR _03417_ sky130_fd_sc_hd__mux2_1
XFILLER_181_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23327_ _09952_ _09953_ _09954_ VGND VGND VPWR VPWR _09956_ sky130_fd_sc_hd__a21oi_1
X_27095_ clknet_leaf_6_B_in_serial_clk _00893_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_186_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20539_ _07436_ _07438_ _07437_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__o21ba_1
XFILLER_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26046_ deser_B.serial_word\[1\] deser_B.shift_reg\[1\] net55 VGND VGND VPWR VPWR
+ _03348_ sky130_fd_sc_hd__mux2_1
X_14060_ deser_B.shift_reg\[94\] deser_B.shift_reg\[95\] net126 VGND VGND VPWR VPWR
+ _00886_ sky130_fd_sc_hd__mux2_1
X_23258_ _09899_ _09902_ VGND VGND VPWR VPWR _09903_ sky130_fd_sc_hd__xor2_1
XFILLER_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_227_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_227_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_238_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22209_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[5\] VGND VGND VPWR
+ VPWR _08955_ sky130_fd_sc_hd__nand2_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23189_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[18\]
+ VGND VGND VPWR VPWR _09844_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_145_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27997_ clknet_leaf_117_clk _01795_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14962_ _12081_ _12082_ VGND VGND VPWR VPWR _12083_ sky130_fd_sc_hd__nor2_1
X_17750_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[26\]
+ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__nand2_1
X_26948_ clknet_leaf_19_A_in_serial_clk _00746_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16701_ _11262_ _04022_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13913_ deser_A.serial_word\[74\] deser_A.shift_reg\[74\] net57 VGND VGND VPWR VPWR
+ _00739_ sky130_fd_sc_hd__mux2_1
X_29667_ clknet_leaf_26_B_in_serial_clk _03462_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_17681_ _04905_ _04910_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__a21oi_1
X_14893_ _11978_ _12013_ VGND VGND VPWR VPWR _12016_ sky130_fd_sc_hd__xor2_1
XFILLER_236_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26879_ clknet_leaf_12_A_in_serial_clk _00677_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19420_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[7\]\[3\]
+ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__nand2_1
X_28618_ clknet_leaf_215_clk _02416_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[166\]
+ sky130_fd_sc_hd__dfrtp_1
X_13844_ deser_A.serial_word\[5\] deser_A.shift_reg\[5\] net58 VGND VGND VPWR VPWR
+ _00670_ sky130_fd_sc_hd__mux2_1
X_16632_ _03954_ _03955_ _03948_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__a21oi_1
XFILLER_207_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29598_ clknet_leaf_14_B_in_serial_clk _03393_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19351_ _06410_ _06409_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__nand2b_1
XFILLER_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28549_ clknet_leaf_178_clk _02347_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_13775_ B_in\[82\] deser_B.word_buffer\[82\] net85 VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16563_ net108 systolic_inst.acc_wires\[12\]\[29\] net67 _03910_ VGND VGND VPWR VPWR
+ _01199_ sky130_fd_sc_hd__a22o_1
XFILLER_222_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18302_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[16\]
+ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__nand2_1
XFILLER_206_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15514_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[7\] _12572_ net116
+ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_204_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_175_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19282_ _06238_ _06342_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__nand2_1
XFILLER_149_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16494_ systolic_inst.acc_wires\[12\]\[16\] systolic_inst.acc_wires\[12\]\[17\] systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__o21ai_1
XFILLER_241_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15445_ net107 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[5\] _12504_
+ _12505_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__a22o_1
X_18233_ _05402_ _05406_ _05409_ _05410_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__o211a_1
XFILLER_175_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15376_ net116 _12440_ VGND VGND VPWR VPWR _12441_ sky130_fd_sc_hd__nand2_1
X_18164_ _05262_ _05350_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__or2_1
XFILLER_156_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17115_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[22\]
+ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__or2_1
XFILLER_15_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14327_ net105 systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[8\] _11512_
+ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__a21o_1
XFILLER_183_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18095_ _05283_ _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__nor2_1
Xmax_cap104 _11302_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_12
XFILLER_184_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap115 net121 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_12
XFILLER_209_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap126 deser_B.receiving VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_130_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17046_ _04337_ _04342_ _04343_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand3_1
XFILLER_116_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14258_ _11437_ _11443_ VGND VGND VPWR VPWR _11445_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_218_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_218_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_217_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13209_ deser_A.word_buffer\[47\] deser_A.serial_word\[47\] net127 VGND VGND VPWR
+ VPWR _00057_ sky130_fd_sc_hd__mux2_1
XFILLER_171_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14189_ _11351_ _11361_ _11363_ VGND VGND VPWR VPWR _11378_ sky130_fd_sc_hd__a21o_1
XFILLER_217_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_163_Left_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18997_ _06086_ _06088_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _05108_ _05140_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_867 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17879_ _05050_ _05073_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19618_ systolic_inst.A_outs\[6\]\[6\] systolic_inst.A_outs\[5\]\[6\] net120 VGND
+ VGND VPWR VPWR _01528_ sky130_fd_sc_hd__mux2_1
XFILLER_53_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20890_ _07766_ _07765_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__and2b_1
XFILLER_148_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19549_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[22\]
+ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__or2_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_234_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_234_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22560_ _09279_ _09281_ _09283_ systolic_inst.acc_wires\[2\]\[13\] net109 VGND VGND
+ VPWR VPWR _01823_ sky130_fd_sc_hd__a32o_1
XFILLER_62_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_172_Left_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1096 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21511_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.A_outs\[3\]\[2\] VGND VGND VPWR
+ VPWR _08324_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_230_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_230_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22491_ net65 _09222_ _09224_ systolic_inst.acc_wires\[2\]\[3\] net109 VGND VGND
+ VPWR VPWR _01813_ sky130_fd_sc_hd__a32o_1
XFILLER_107_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24230_ _10600_ systolic_inst.A_shift\[19\]\[6\] net70 VGND VGND VPWR VPWR _02176_
+ sky130_fd_sc_hd__mux2_1
X_21442_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[28\]
+ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__or2_1
XFILLER_33_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24161_ systolic_inst.A_shift\[28\]\[4\] A_in\[100\] net59 VGND VGND VPWR VPWR _10582_
+ sky130_fd_sc_hd__mux2_1
X_21373_ _11258_ systolic_inst.acc_wires\[4\]\[17\] net63 _08220_ VGND VGND VPWR VPWR
+ _01699_ sky130_fd_sc_hd__a22o_1
XFILLER_162_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23112_ net64 _09776_ _09778_ systolic_inst.acc_wires\[1\]\[6\] _11258_ VGND VGND
+ VPWR VPWR _01880_ sky130_fd_sc_hd__a32o_1
XFILLER_194_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20324_ systolic_inst.A_outs\[5\]\[2\] systolic_inst.B_outs\[5\]\[3\] systolic_inst.A_outs\[5\]\[3\]
+ systolic_inst.B_outs\[5\]\[4\] VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__nand4_2
XFILLER_163_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24092_ _10555_ systolic_inst.B_shift\[19\]\[1\] net71 VGND VGND VPWR VPWR _02083_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_209_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_209_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_181_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27920_ clknet_leaf_146_clk _01718_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_23043_ _09627_ _09716_ VGND VGND VPWR VPWR _09718_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20255_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.A_outs\[5\]\[1\] systolic_inst.B_outs\[5\]\[2\]
+ systolic_inst.B_outs\[5\]\[3\] VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_181_Left_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20186_ net62 _07152_ _07153_ systolic_inst.acc_wires\[6\]\[25\] net106 VGND VGND
+ VPWR VPWR _01579_ sky130_fd_sc_hd__a32o_1
X_27851_ clknet_leaf_181_clk _01649_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26802_ clknet_leaf_88_clk _00604_ net5 VGND VGND VPWR VPWR B_in\[74\] sky130_fd_sc_hd__dfrtp_1
XFILLER_131_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27782_ clknet_leaf_187_clk _01580_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_24994_ net111 ser_C.shift_reg\[325\] VGND VGND VPWR VPWR _10967_ sky130_fd_sc_hd__and2_1
XFILLER_229_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29521_ clknet_leaf_256_clk _03319_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[493\]
+ sky130_fd_sc_hd__dfrtp_1
X_26733_ clknet_leaf_97_clk _00535_ net153 VGND VGND VPWR VPWR B_in\[5\] sky130_fd_sc_hd__dfrtp_1
X_23945_ _10501_ systolic_inst.B_shift\[10\]\[4\] _11332_ VGND VGND VPWR VPWR _01990_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26664_ clknet_leaf_4_B_in_serial_clk _00467_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_29452_ clknet_leaf_290_clk _03250_ net136 VGND VGND VPWR VPWR C_out\[424\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23876_ _10463_ _10464_ VGND VGND VPWR VPWR _10465_ sky130_fd_sc_hd__nand2_1
XFILLER_29_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25615_ systolic_inst.acc_wires\[2\]\[27\] C_out\[91\] net51 VGND VGND VPWR VPWR
+ _02917_ sky130_fd_sc_hd__mux2_1
X_28403_ clknet_leaf_33_clk _02201_ VGND VGND VPWR VPWR systolic_inst.A_shift\[16\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_22827_ _09507_ _09508_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__nand2b_1
XFILLER_72_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26595_ clknet_leaf_0_A_in_serial_clk _00398_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[125\]
+ sky130_fd_sc_hd__dfrtp_1
X_29383_ clknet_leaf_245_clk _03181_ net145 VGND VGND VPWR VPWR C_out\[355\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_190_Left_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25546_ systolic_inst.acc_wires\[0\]\[22\] C_out\[22\] net54 VGND VGND VPWR VPWR
+ _02848_ sky130_fd_sc_hd__mux2_1
XFILLER_198_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28334_ clknet_leaf_342_clk _02132_ VGND VGND VPWR VPWR systolic_inst.A_shift\[26\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13560_ deser_A.shift_reg\[124\] deser_A.shift_reg\[125\] net130 VGND VGND VPWR VPWR
+ _00397_ sky130_fd_sc_hd__mux2_1
XFILLER_240_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22758_ _09411_ _09414_ _09441_ VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__o21a_1
XFILLER_197_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21709_ _08443_ _08514_ VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__and2_1
X_28265_ clknet_leaf_52_clk _02063_ VGND VGND VPWR VPWR systolic_inst.B_shift\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_27_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_27_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_73_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25477_ systolic_inst.cycle_cnt\[15\] systolic_inst.cycle_cnt\[14\] _11210_ VGND
+ VGND VPWR VPWR _11215_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_188_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13491_ deser_A.shift_reg\[55\] deser_A.shift_reg\[56\] net130 VGND VGND VPWR VPWR
+ _00328_ sky130_fd_sc_hd__mux2_1
X_22689_ net122 systolic_inst.B_outs\[1\]\[0\] systolic_inst.A_outs\[1\]\[0\] VGND
+ VGND VPWR VPWR _09378_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_188_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15230_ _12329_ _12330_ VGND VGND VPWR VPWR _12332_ sky130_fd_sc_hd__nand2_1
XFILLER_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24428_ net114 ser_C.shift_reg\[42\] VGND VGND VPWR VPWR _10684_ sky130_fd_sc_hd__and2_1
XFILLER_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27216_ clknet_leaf_292_clk _01014_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_28196_ clknet_leaf_47_clk _01994_ VGND VGND VPWR VPWR systolic_inst.B_shift\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15161_ _12272_ VGND VGND VPWR VPWR _12273_ sky130_fd_sc_hd__inv_2
X_27147_ clknet_leaf_4_clk _00945_ VGND VGND VPWR VPWR systolic_inst.A_shift\[21\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_24359_ C_out\[6\] net104 _10643_ ser_C.shift_reg\[6\] _10649_ VGND VGND VPWR VPWR
+ _02256_ sky130_fd_sc_hd__a221o_1
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14112_ systolic_inst.B_shift\[12\]\[4\] net72 _11333_ B_in\[100\] VGND VGND VPWR
+ VPWR _00934_ sky130_fd_sc_hd__a22o_1
XFILLER_153_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27078_ clknet_leaf_27_B_in_serial_clk _00876_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_15092_ _12207_ _12208_ VGND VGND VPWR VPWR _12209_ sky130_fd_sc_hd__nor2_1
XFILLER_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14043_ deser_B.shift_reg\[77\] deser_B.shift_reg\[78\] deser_B.receiving VGND VGND
+ VPWR VPWR _00869_ sky130_fd_sc_hd__mux2_1
XFILLER_181_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26029_ systolic_inst.acc_wires\[15\]\[25\] ser_C.parallel_data\[505\] net37 VGND
+ VGND VPWR VPWR _03331_ sky130_fd_sc_hd__mux2_1
X_18920_ _06021_ _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18851_ _05956_ _05960_ _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__a21o_1
XFILLER_122_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_164_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17802_ net107 systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[0\] _05002_
+ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__a21o_1
X_18782_ _05902_ _05903_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__and2b_1
X_15994_ systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[3\] VGND VGND
+ VPWR VPWR _12993_ sky130_fd_sc_hd__nand2_1
XFILLER_125_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17733_ _04950_ _04954_ _04957_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14945_ _12065_ _12064_ VGND VGND VPWR VPWR _12067_ sky130_fd_sc_hd__nand2b_1
XFILLER_208_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17664_ _04894_ _04898_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__nand2b_1
XFILLER_21_1260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14876_ _11997_ _11998_ VGND VGND VPWR VPWR _11999_ sky130_fd_sc_hd__nor2_1
X_19403_ net119 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[7\]\[0\]
+ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16615_ _03934_ _03939_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__xnor2_1
X_13827_ deser_B.bit_idx\[1\] deser_B.bit_idx\[2\] _11319_ VGND VGND VPWR VPWR _11323_
+ sky130_fd_sc_hd__and3_1
XFILLER_165_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17595_ _04838_ _04839_ _04840_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__a21o_1
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19334_ _06306_ _06365_ _06364_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__a21oi_1
X_13758_ B_in\[65\] deser_B.word_buffer\[65\] net87 VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__mux2_1
X_16546_ _03893_ _03896_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19265_ _06276_ _06293_ _06291_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__o21a_1
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13689_ deser_B.word_buffer\[125\] deser_B.serial_word\[125\] net123 VGND VGND VPWR
+ VPWR _00526_ sky130_fd_sc_hd__mux2_1
X_16477_ _03814_ _03819_ _03820_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__a21boi_1
XFILLER_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18216_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[9\]\[4\]
+ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__nand2_1
X_15428_ systolic_inst.A_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[2\] systolic_inst.B_outs\[13\]\[3\]
+ systolic_inst.B_outs\[13\]\[4\] VGND VGND VPWR VPWR _12489_ sky130_fd_sc_hd__and4_1
X_19196_ _06242_ _06259_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15359_ systolic_inst.A_outs\[13\]\[3\] systolic_inst.A_outs\[12\]\[3\] net115 VGND
+ VGND VPWR VPWR _01077_ sky130_fd_sc_hd__mux2_1
X_18147_ _05292_ _05334_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18078_ _05227_ _05229_ _05228_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17029_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[11\]\[8\]
+ _04329_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__and3_1
XFILLER_217_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20040_ _07026_ _07027_ _07028_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__a21o_1
XFILLER_63_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1002 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21991_ _08772_ _08773_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__nand2_1
XFILLER_27_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_236_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23730_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[0\]\[6\]
+ VGND VGND VPWR VPWR _10341_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_236_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[6\]
+ systolic_inst.B_outs\[4\]\[6\] VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_236_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_232_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _10250_ _10253_ VGND VGND VPWR VPWR _10281_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20873_ systolic_inst.A_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[3\]
+ systolic_inst.B_outs\[4\]\[4\] VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__and4_1
XFILLER_148_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25400_ _11169_ systolic_inst.A_shift\[2\]\[7\] net71 VGND VGND VPWR VPWR _02777_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22612_ _09325_ _09326_ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__and2_1
XFILLER_228_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26380_ clknet_leaf_21_clk _00187_ net133 VGND VGND VPWR VPWR A_in\[48\] sky130_fd_sc_hd__dfrtp_1
X_23592_ _10211_ _10212_ _10148_ _10151_ VGND VGND VPWR VPWR _10214_ sky130_fd_sc_hd__o211a_1
XFILLER_34_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25331_ ser_C.parallel_data\[492\] net97 net77 ser_C.shift_reg\[492\] _11135_ VGND
+ VGND VPWR VPWR _02742_ sky130_fd_sc_hd__a221o_1
X_22543_ _09267_ _09268_ VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28050_ clknet_leaf_128_clk _01848_ net142 VGND VGND VPWR VPWR systolic_inst.A_outs\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_25262_ net111 ser_C.shift_reg\[459\] VGND VGND VPWR VPWR _11101_ sky130_fd_sc_hd__and2_1
XFILLER_10_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22474_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[2\]\[0\]
+ _09208_ _09209_ VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__and4_1
X_27001_ clknet_leaf_15_B_in_serial_clk _00799_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24213_ systolic_inst.A_shift\[21\]\[6\] A_in\[86\] net59 VGND VGND VPWR VPWR _10592_
+ sky130_fd_sc_hd__mux2_1
XFILLER_148_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21425_ _08260_ _08262_ _08264_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__or3_1
XFILLER_135_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25193_ C_out\[423\] net102 net74 ser_C.shift_reg\[423\] _11066_ VGND VGND VPWR VPWR
+ _02673_ sky130_fd_sc_hd__a221o_1
XFILLER_163_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24144_ _10573_ systolic_inst.A_shift\[28\]\[3\] net70 VGND VGND VPWR VPWR _02117_
+ sky130_fd_sc_hd__mux2_1
X_21356_ _08198_ _08202_ _08204_ _08205_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__a211o_1
XFILLER_151_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20307_ _07222_ _07245_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__xor2_1
XFILLER_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24075_ systolic_inst.B_shift\[3\]\[2\] _11332_ net83 systolic_inst.B_shift\[7\]\[2\]
+ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__a22o_1
X_28952_ clknet_leaf_263_clk _02750_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[500\]
+ sky130_fd_sc_hd__dfrtp_1
X_21287_ _08137_ _08141_ _08144_ _08145_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__o211a_1
XFILLER_104_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23026_ _09701_ _09700_ VGND VGND VPWR VPWR _09702_ sky130_fd_sc_hd__and2b_1
X_27903_ clknet_leaf_42_clk _01701_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_20238_ systolic_inst.B_outs\[4\]\[7\] systolic_inst.B_outs\[0\]\[7\] net117 VGND
+ VGND VPWR VPWR _01601_ sky130_fd_sc_hd__mux2_1
X_28883_ clknet_leaf_329_clk _02681_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[431\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27834_ clknet_leaf_145_clk _01632_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_20169_ _07131_ _07135_ _07138_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__nand3_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27765_ clknet_leaf_210_clk _01563_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24977_ C_out\[315\] net103 net76 ser_C.shift_reg\[315\] _10958_ VGND VGND VPWR VPWR
+ _02565_ sky130_fd_sc_hd__a221o_1
XFILLER_58_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29504_ clknet_leaf_266_clk _03302_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[476\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26716_ clknet_leaf_29_B_in_serial_clk _00519_ net135 VGND VGND VPWR VPWR deser_B.word_buffer\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14730_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[30\]
+ VGND VGND VPWR VPWR _11878_ sky130_fd_sc_hd__nand2_1
X_23928_ systolic_inst.A_shift\[3\]\[0\] net71 _11333_ A_in\[24\] VGND VGND VPWR VPWR
+ _01978_ sky130_fd_sc_hd__a22o_1
X_27696_ clknet_leaf_196_clk _01494_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14661_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[20\]
+ VGND VGND VPWR VPWR _11819_ sky130_fd_sc_hd__or2_1
X_29435_ clknet_leaf_335_clk _03233_ net131 VGND VGND VPWR VPWR C_out\[407\] sky130_fd_sc_hd__dfrtp_1
X_23859_ net64 _10449_ _10450_ systolic_inst.acc_wires\[0\]\[25\] _11258_ VGND VGND
+ VPWR VPWR _01955_ sky130_fd_sc_hd__a32o_1
X_26647_ clknet_leaf_20_B_in_serial_clk _00450_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13612_ deser_B.word_buffer\[48\] deser_B.serial_word\[48\] net124 VGND VGND VPWR
+ VPWR _00449_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _03763_ _03766_ _03768_ _03770_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__o211a_1
XFILLER_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29366_ clknet_leaf_202_clk _03164_ net147 VGND VGND VPWR VPWR C_out\[338\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14592_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[15\]\[10\]
+ VGND VGND VPWR VPWR _11760_ sky130_fd_sc_hd__nand2_1
X_17380_ _04635_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__nor2_1
X_26578_ clknet_leaf_28_A_in_serial_clk _00381_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16331_ _03709_ _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__and2b_1
X_13543_ deser_A.shift_reg\[107\] deser_A.shift_reg\[108\] net129 VGND VGND VPWR VPWR
+ _00380_ sky130_fd_sc_hd__mux2_1
X_28317_ clknet_leaf_2_clk _02115_ VGND VGND VPWR VPWR systolic_inst.A_shift\[28\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25529_ systolic_inst.acc_wires\[0\]\[5\] C_out\[5\] net33 VGND VGND VPWR VPWR _02831_
+ sky130_fd_sc_hd__mux2_1
X_29297_ clknet_leaf_310_clk _03095_ net142 VGND VGND VPWR VPWR C_out\[269\] sky130_fd_sc_hd__dfrtp_1
XFILLER_186_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19050_ _06114_ _06119_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__nand2_1
X_16262_ _03603_ _03605_ _03642_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__nand3_1
X_28248_ clknet_leaf_80_clk _02046_ VGND VGND VPWR VPWR systolic_inst.B_shift\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13474_ deser_A.shift_reg\[38\] deser_A.shift_reg\[39\] deser_A.receiving VGND VGND
+ VPWR VPWR _00311_ sky130_fd_sc_hd__mux2_1
XFILLER_16_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15213_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[14\]\[9\]
+ _12312_ VGND VGND VPWR VPWR _12317_ sky130_fd_sc_hd__a21oi_1
X_18001_ systolic_inst.B_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[5\]
+ systolic_inst.A_outs\[9\]\[6\] VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__and4_1
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16193_ _03559_ _03576_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__xor2_1
XFILLER_154_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28179_ clknet_leaf_62_clk _01977_ VGND VGND VPWR VPWR systolic_inst.B_shift\[18\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15144_ net107 _12248_ _12258_ VGND VGND VPWR VPWR _12259_ sky130_fd_sc_hd__or3_1
XFILLER_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19952_ _06883_ _06888_ _06916_ _06947_ _06914_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_112_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15075_ _12192_ _12191_ VGND VGND VPWR VPWR _12193_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_166_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14026_ deser_B.shift_reg\[60\] deser_B.shift_reg\[61\] deser_B.receiving VGND VGND
+ VPWR VPWR _00852_ sky130_fd_sc_hd__mux2_1
X_18903_ _06001_ _06005_ _06007_ _06008_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__a211o_1
X_19883_ _06820_ _06845_ _06844_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__a21boi_1
XFILLER_150_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_27__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_27__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_18834_ _05940_ _05944_ _05947_ _05948_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__o211a_1
XFILLER_228_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18765_ _05856_ _05861_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__or3_1
X_15977_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.A_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\]
+ systolic_inst.A_outs\[12\]\[1\] VGND VGND VPWR VPWR _12978_ sky130_fd_sc_hd__and4_1
XFILLER_83_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17716_ _11712_ _04943_ _04944_ systolic_inst.acc_wires\[10\]\[20\] net106 VGND VGND
+ VPWR VPWR _01318_ sky130_fd_sc_hd__a32o_1
XFILLER_208_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14928_ _12040_ _12048_ VGND VGND VPWR VPWR _12050_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18696_ _05821_ _05820_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__and2b_1
XFILLER_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17647_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[10\]\[11\]
+ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__nand2_1
XFILLER_224_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14859_ _11938_ _11940_ _11982_ VGND VGND VPWR VPWR _11983_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17578_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[10\]\[1\]
+ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__and2_1
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19317_ systolic_inst.A_outs\[7\]\[5\] systolic_inst.B_outs\[7\]\[6\] systolic_inst.A_outs\[7\]\[6\]
+ systolic_inst.B_outs\[7\]\[7\] VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__and4b_1
X_16529_ systolic_inst.acc_wires\[12\]\[22\] systolic_inst.acc_wires\[12\]\[23\] systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__o21a_1
XFILLER_220_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19248_ systolic_inst.A_outs\[7\]\[6\] _06310_ _06309_ VGND VGND VPWR VPWR _06311_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_108_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19179_ systolic_inst.B_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[5\]
+ systolic_inst.B_outs\[7\]\[3\] VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__a22oi_1
XFILLER_30_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21210_ _08042_ _08043_ _08045_ _08046_ _08030_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_22_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22190_ _08906_ _08935_ _08936_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__nand3_1
XFILLER_191_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_225_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_225_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21141_ _08000_ _08010_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21072_ _07941_ _07942_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20023_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[6\]\[2\]
+ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__nand2_1
X_24900_ net110 ser_C.shift_reg\[278\] VGND VGND VPWR VPWR _10920_ sky130_fd_sc_hd__and2_1
X_25880_ systolic_inst.acc_wires\[11\]\[4\] C_out\[356\] net38 VGND VGND VPWR VPWR
+ _03182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_238_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24831_ C_out\[242\] net98 net78 ser_C.shift_reg\[242\] _10885_ VGND VGND VPWR VPWR
+ _02492_ sky130_fd_sc_hd__a221o_1
XFILLER_41_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24762_ net113 ser_C.shift_reg\[209\] VGND VGND VPWR VPWR _10851_ sky130_fd_sc_hd__and2_1
X_27550_ clknet_leaf_299_clk _01348_ net139 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_100_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21974_ _08731_ _08733_ _08735_ _08738_ _08758_ VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__o311a_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23713_ _10326_ VGND VGND VPWR VPWR _10327_ sky130_fd_sc_hd__inv_2
X_26501_ clknet_leaf_12_A_in_serial_clk _00304_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27481_ clknet_leaf_41_clk _01279_ net142 VGND VGND VPWR VPWR systolic_inst.B_outs\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_27_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20925_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[5\] _07800_ net117
+ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__mux2_1
X_24693_ C_out\[173\] net104 net76 ser_C.shift_reg\[173\] _10816_ VGND VGND VPWR VPWR
+ _02423_ sky130_fd_sc_hd__a221o_1
XFILLER_27_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29220_ clknet_leaf_207_clk _03018_ net147 VGND VGND VPWR VPWR C_out\[192\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23644_ _10195_ _10263_ VGND VGND VPWR VPWR _10264_ sky130_fd_sc_hd__or2_1
X_26432_ clknet_leaf_0_clk _00239_ net134 VGND VGND VPWR VPWR A_in\[100\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20856_ _07725_ _07733_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__and2_1
XFILLER_214_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29151_ clknet_leaf_172_clk _02949_ net148 VGND VGND VPWR VPWR C_out\[123\] sky130_fd_sc_hd__dfrtp_1
X_26363_ clknet_leaf_19_clk _00170_ net133 VGND VGND VPWR VPWR A_in\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_167_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23575_ _11267_ systolic_inst.B_outs\[0\]\[7\] _10120_ VGND VGND VPWR VPWR _10197_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_23_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20787_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[25\]
+ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_214_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28102_ clknet_leaf_111_clk _01900_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_214_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25314_ net112 ser_C.shift_reg\[485\] VGND VGND VPWR VPWR _11127_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_214_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22526_ _09249_ _09252_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__nand2_1
XFILLER_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29082_ clknet_leaf_110_clk _02880_ net151 VGND VGND VPWR VPWR C_out\[54\] sky130_fd_sc_hd__dfrtp_1
XFILLER_195_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26294_ clknet_leaf_2_A_in_serial_clk _00102_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28033_ clknet_leaf_158_clk _01831_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_210_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25245_ ser_C.parallel_data\[449\] net102 net74 ser_C.shift_reg\[449\] _11092_ VGND
+ VGND VPWR VPWR _02699_ sky130_fd_sc_hd__a221o_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22457_ _09193_ _09194_ VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_210_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21408_ net63 _08249_ _08250_ systolic_inst.acc_wires\[4\]\[22\] _11258_ VGND VGND
+ VPWR VPWR _01704_ sky130_fd_sc_hd__a32o_1
XFILLER_202_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13190_ deser_A.word_buffer\[28\] deser_A.serial_word\[28\] net128 VGND VGND VPWR
+ VPWR _00038_ sky130_fd_sc_hd__mux2_1
X_25176_ net111 ser_C.shift_reg\[416\] VGND VGND VPWR VPWR _11058_ sky130_fd_sc_hd__and2_1
XFILLER_203_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22388_ _09127_ _09128_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__nor2_1
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24127_ systolic_inst.A_shift\[30\]\[3\] A_in\[115\] net59 VGND VGND VPWR VPWR _10565_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21339_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[4\]\[13\]
+ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__or2_1
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24058_ _10546_ systolic_inst.B_shift\[15\]\[0\] net70 VGND VGND VPWR VPWR _02058_
+ sky130_fd_sc_hd__mux2_1
X_28935_ clknet_leaf_261_clk _02733_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23009_ net109 systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[12\] _09683_
+ _09685_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__a22o_1
X_15900_ _12919_ _12920_ VGND VGND VPWR VPWR _12928_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_161_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28866_ clknet_leaf_332_clk _02664_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[414\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16880_ _04056_ _04196_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__or2_1
XFILLER_103_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27817_ clknet_leaf_143_clk _01615_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_15831_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[13\]\[12\]
+ VGND VGND VPWR VPWR _12869_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28797_ clknet_leaf_234_clk _02595_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[345\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18550_ _05641_ _05677_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__xor2_1
X_27748_ clknet_leaf_209_clk _01546_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15762_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[13\]\[0\]
+ _12804_ _12802_ VGND VGND VPWR VPWR _12810_ sky130_fd_sc_hd__a31o_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17501_ _04721_ _04723_ _04752_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__nand3_1
XFILLER_233_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14713_ net105 systolic_inst.acc_wires\[15\]\[27\] net69 _11863_ VGND VGND VPWR VPWR
+ _01005_ sky130_fd_sc_hd__a22o_1
X_18481_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[5\] _05610_ _05611_
+ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_206_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27679_ clknet_leaf_234_clk _01477_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15693_ systolic_inst.B_outs\[13\]\[6\] systolic_inst.A_outs\[13\]\[7\] VGND VGND
+ VPWR VPWR _12746_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_159_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29418_ clknet_leaf_333_clk _03216_ net131 VGND VGND VPWR VPWR C_out\[390\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17432_ _04678_ _04686_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__nand2_1
X_14644_ net107 systolic_inst.acc_wires\[15\]\[16\] _11803_ _11805_ VGND VGND VPWR
+ VPWR _00994_ sky130_fd_sc_hd__a22o_1
XFILLER_205_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14575_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[15\]\[7\]
+ VGND VGND VPWR VPWR _11746_ sky130_fd_sc_hd__or2_1
X_29349_ clknet_leaf_294_clk _03147_ net138 VGND VGND VPWR VPWR C_out\[321\] sky130_fd_sc_hd__dfrtp_1
X_17363_ _04611_ _04619_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__nand2_1
XFILLER_92_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19102_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[3\] _06153_ _06151_
+ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__a31o_1
X_16314_ _03662_ _03665_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__o21ai_1
XFILLER_242_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13526_ deser_A.shift_reg\[90\] deser_A.shift_reg\[91\] net129 VGND VGND VPWR VPWR
+ _00363_ sky130_fd_sc_hd__mux2_1
X_17294_ _04550_ _04551_ _04521_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__a21o_1
XFILLER_186_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19033_ net105 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _06104_ sky130_fd_sc_hd__and2_1
X_13457_ deser_A.shift_reg\[21\] deser_A.shift_reg\[22\] deser_A.receiving VGND VGND
+ VPWR VPWR _00294_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16245_ _03517_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__or2_1
XFILLER_220_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16176_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[7\] VGND VGND
+ VPWR VPWR _03560_ sky130_fd_sc_hd__nand2_4
X_13388_ A_in\[97\] deser_A.word_buffer\[97\] net96 VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15127_ _12242_ _12241_ VGND VGND VPWR VPWR _12243_ sky130_fd_sc_hd__and2b_1
XFILLER_142_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19935_ _06929_ _06930_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__xnor2_1
X_15058_ _12174_ _12175_ VGND VGND VPWR VPWR _12176_ sky130_fd_sc_hd__nand2_1
XFILLER_141_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_220_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_220_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14009_ deser_B.shift_reg\[43\] deser_B.shift_reg\[44\] net125 VGND VGND VPWR VPWR
+ _00835_ sky130_fd_sc_hd__mux2_1
XFILLER_123_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19866_ _06861_ _06864_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__xnor2_1
XFILLER_229_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18817_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[8\]\[3\]
+ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__nand2_1
XFILLER_233_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19797_ systolic_inst.A_outs\[6\]\[2\] systolic_inst.B_outs\[6\]\[5\] _06760_ _06759_
+ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_108_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18748_ _05869_ _05870_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__xnor2_1
XFILLER_237_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_218_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18679_ _05768_ _05804_ systolic_inst.A_outs\[8\]\[7\] VGND VGND VPWR VPWR _05805_
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_218_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_218_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20710_ _11713_ _07625_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__nor2_1
XFILLER_91_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21690_ _08489_ _08497_ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20641_ _07562_ _07563_ _07564_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__a21o_1
XFILLER_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23360_ _09959_ _09987_ VGND VGND VPWR VPWR _09988_ sky130_fd_sc_hd__nand2_1
X_20572_ _07502_ _07503_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22311_ net122 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[9\] _09053_
+ _09054_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_227_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23291_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.A_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\]
+ systolic_inst.A_outs\[0\]\[0\] VGND VGND VPWR VPWR _09922_ sky130_fd_sc_hd__a22o_1
XFILLER_192_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25030_ net112 ser_C.shift_reg\[343\] VGND VGND VPWR VPWR _10985_ sky130_fd_sc_hd__and2_1
X_22242_ _08986_ _08983_ VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__and2b_1
XFILLER_30_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22173_ _08919_ _08916_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__and2b_1
XFILLER_191_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21124_ _07989_ _07993_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_58_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26981_ clknet_leaf_29_A_in_serial_clk _00779_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_236_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28720_ clknet_leaf_310_clk _02518_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21055_ systolic_inst.A_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[6\] VGND VGND VPWR
+ VPWR _07927_ sky130_fd_sc_hd__nand2_1
X_25932_ systolic_inst.acc_wires\[12\]\[24\] C_out\[408\] net17 VGND VGND VPWR VPWR
+ _03234_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20006_ _06782_ _06920_ _06991_ _06989_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__a31o_1
XFILLER_219_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28651_ clknet_leaf_202_clk _02449_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[199\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_5_10__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_10__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25863_ systolic_inst.acc_wires\[10\]\[19\] C_out\[339\] net11 VGND VGND VPWR VPWR
+ _03165_ sky130_fd_sc_hd__mux2_1
XFILLER_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27602_ clknet_leaf_319_clk _01400_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_234_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24814_ net113 ser_C.shift_reg\[235\] VGND VGND VPWR VPWR _10877_ sky130_fd_sc_hd__and2_1
XFILLER_74_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28582_ clknet_leaf_308_clk _02380_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[130\]
+ sky130_fd_sc_hd__dfrtp_1
X_25794_ systolic_inst.acc_wires\[8\]\[14\] C_out\[270\] net28 VGND VGND VPWR VPWR
+ _03096_ sky130_fd_sc_hd__mux2_1
XFILLER_228_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27533_ clknet_leaf_312_clk _01331_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_21957_ _08737_ _08740_ _08744_ VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_195_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24745_ C_out\[199\] net97 net80 ser_C.shift_reg\[199\] _10842_ VGND VGND VPWR VPWR
+ _02449_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_226_Right_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20908_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[5\] _07782_ _07783_
+ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__nand4_2
X_24676_ net111 ser_C.shift_reg\[166\] VGND VGND VPWR VPWR _10808_ sky130_fd_sc_hd__and2_1
X_27464_ clknet_leaf_238_clk _01262_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_230_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21888_ _08676_ _08680_ _08683_ _08684_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__o211a_1
XFILLER_163_1318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29203_ clknet_leaf_145_clk _03001_ net149 VGND VGND VPWR VPWR C_out\[175\] sky130_fd_sc_hd__dfrtp_1
X_23627_ _10246_ _10247_ VGND VGND VPWR VPWR _10248_ sky130_fd_sc_hd__nand2_1
XFILLER_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26415_ clknet_leaf_5_clk _00222_ net131 VGND VGND VPWR VPWR A_in\[83\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_212_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ systolic_inst.B_outs\[3\]\[4\] systolic_inst.B_shift\[3\]\[4\] net120 VGND
+ VGND VPWR VPWR _01662_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_212_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27395_ clknet_leaf_336_clk _01193_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_204_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29134_ clknet_leaf_170_clk _02932_ net148 VGND VGND VPWR VPWR C_out\[106\] sky130_fd_sc_hd__dfrtp_1
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _11514_ _11543_ VGND VGND VPWR VPWR _11545_ sky130_fd_sc_hd__xnor2_1
X_23558_ _10178_ _10179_ _10180_ VGND VGND VPWR VPWR _10181_ sky130_fd_sc_hd__o21bai_1
X_26346_ clknet_leaf_20_clk _00153_ net135 VGND VGND VPWR VPWR A_in\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ A_in\[20\] deser_A.word_buffer\[20\] net92 VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__mux2_1
XFILLER_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22509_ _09237_ _09238_ _09239_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__a21o_1
XFILLER_195_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29065_ clknet_leaf_115_clk _02863_ net152 VGND VGND VPWR VPWR C_out\[37\] sky130_fd_sc_hd__dfrtp_1
XFILLER_195_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14291_ systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[6\] systolic_inst.A_outs\[15\]\[7\]
+ systolic_inst.B_outs\[15\]\[1\] VGND VGND VPWR VPWR _11477_ sky130_fd_sc_hd__a22o_1
X_26277_ clknet_leaf_20_A_in_serial_clk _00085_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_156_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23489_ _10111_ _10112_ VGND VGND VPWR VPWR _10113_ sky130_fd_sc_hd__nand2_1
XFILLER_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28016_ clknet_leaf_152_clk _01814_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_16030_ _13004_ _13006_ _13005_ VGND VGND VPWR VPWR _13027_ sky130_fd_sc_hd__a21bo_1
X_13242_ deser_A.word_buffer\[80\] deser_A.serial_word\[80\] net127 VGND VGND VPWR
+ VPWR _00090_ sky130_fd_sc_hd__mux2_1
XFILLER_109_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25228_ net111 ser_C.shift_reg\[442\] VGND VGND VPWR VPWR _11084_ sky130_fd_sc_hd__and2_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13173_ deser_A.word_buffer\[11\] deser_A.serial_word\[11\] net128 VGND VGND VPWR
+ VPWR _00021_ sky130_fd_sc_hd__mux2_1
X_25159_ C_out\[406\] net101 net73 ser_C.shift_reg\[406\] _11049_ VGND VGND VPWR VPWR
+ _02656_ sky130_fd_sc_hd__a221o_1
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17981_ _05118_ _05133_ _05132_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_148_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19720_ _06721_ _06722_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__or2_1
XFILLER_117_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28918_ clknet_leaf_282_clk _02716_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16932_ _04215_ _04218_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__nor3_1
XFILLER_137_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19651_ _06654_ _06655_ _06643_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__a21o_1
X_28849_ clknet_leaf_338_clk _02647_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[397\]
+ sky130_fd_sc_hd__dfrtp_1
X_16863_ _04141_ _04143_ _04179_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__nand3_1
XFILLER_78_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18602_ _05692_ _05698_ _05697_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__a21o_1
X_15814_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[13\]\[10\]
+ VGND VGND VPWR VPWR _12854_ sky130_fd_sc_hd__or2_1
XFILLER_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19582_ net106 systolic_inst.acc_wires\[7\]\[26\] net62 _06612_ VGND VGND VPWR VPWR
+ _01516_ sky130_fd_sc_hd__a22o_1
X_16794_ _04112_ _04113_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__and2b_1
XFILLER_93_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18533_ _05657_ _05661_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_103_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _12713_ _12775_ VGND VGND VPWR VPWR _12796_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_A_in_serial_clk clknet_2_3__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_12_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_46_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18464_ _05594_ _05595_ _05573_ _05576_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_64_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15676_ _12716_ _12729_ VGND VGND VPWR VPWR _12730_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_64_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17415_ net105 _04668_ _04669_ _04670_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__o31a_1
XFILLER_33_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14627_ _11783_ _11790_ VGND VGND VPWR VPWR _11791_ sky130_fd_sc_hd__nand2_1
X_18395_ _05548_ _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__nand2_1
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17346_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] _04602_ VGND
+ VGND VPWR VPWR _04603_ sky130_fd_sc_hd__a21o_1
X_14558_ _11731_ VGND VGND VPWR VPWR _11732_ sky130_fd_sc_hd__inv_2
XFILLER_201_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13509_ deser_A.shift_reg\[73\] deser_A.shift_reg\[74\] net129 VGND VGND VPWR VPWR
+ _00346_ sky130_fd_sc_hd__mux2_1
X_17277_ _04531_ _04534_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__xnor2_1
Xclkload202 clknet_leaf_70_clk VGND VGND VPWR VPWR clkload202/X sky130_fd_sc_hd__clkbuf_4
X_14489_ _11620_ _11669_ VGND VGND VPWR VPWR _11670_ sky130_fd_sc_hd__xnor2_1
Xclkload213 clknet_leaf_47_clk VGND VGND VPWR VPWR clkload213/X sky130_fd_sc_hd__clkbuf_4
Xclkload224 clknet_leaf_134_clk VGND VGND VPWR VPWR clkload224/X sky130_fd_sc_hd__clkbuf_8
X_19016_ systolic_inst.A_outs\[7\]\[5\] systolic_inst.A_outs\[6\]\[5\] net119 VGND
+ VGND VPWR VPWR _01463_ sky130_fd_sc_hd__mux2_1
X_16228_ _03592_ _03610_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__xor2_1
Xclkload235 clknet_leaf_86_clk VGND VGND VPWR VPWR clkload235/X sky130_fd_sc_hd__clkbuf_4
Xclkload246 clknet_leaf_122_clk VGND VGND VPWR VPWR clkload246/Y sky130_fd_sc_hd__bufinv_16
Xclkload257 clknet_leaf_100_clk VGND VGND VPWR VPWR clkload257/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload268 clknet_leaf_138_clk VGND VGND VPWR VPWR clkload268/Y sky130_fd_sc_hd__inv_4
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload279 clknet_leaf_206_clk VGND VGND VPWR VPWR clkload279/Y sky130_fd_sc_hd__clkinv_4
XFILLER_155_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16159_ _03543_ _03513_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__nand2b_1
XFILLER_170_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19918_ _06915_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__inv_2
XFILLER_130_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19849_ _06847_ _06848_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__nor2_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22860_ _09539_ _09540_ VGND VGND VPWR VPWR _09541_ sky130_fd_sc_hd__nand2b_1
XFILLER_3_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21811_ systolic_inst.B_outs\[3\]\[6\] systolic_inst.A_outs\[3\]\[7\] VGND VGND VPWR
+ VPWR _08615_ sky130_fd_sc_hd__nand2_1
XFILLER_225_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22791_ _09440_ _09442_ _09472_ _09473_ VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__o211a_1
XFILLER_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24530_ net114 ser_C.shift_reg\[93\] VGND VGND VPWR VPWR _10735_ sky130_fd_sc_hd__and2_1
XFILLER_240_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21742_ net106 _08548_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__nor2_1
XFILLER_64_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24461_ C_out\[57\] net100 net82 ser_C.shift_reg\[57\] _10700_ VGND VGND VPWR VPWR
+ _02307_ sky130_fd_sc_hd__a221o_1
X_21673_ _08449_ _08451_ _08448_ VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_190_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23412_ _10034_ _10037_ VGND VGND VPWR VPWR _10038_ sky130_fd_sc_hd__xnor2_1
X_26200_ systolic_inst.A_shift\[30\]\[6\] net71 _11333_ A_in\[126\] VGND VGND VPWR
+ VPWR _03490_ sky130_fd_sc_hd__a22o_1
XFILLER_123_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20624_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[5\]\[1\]
+ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__or2_1
X_27180_ clknet_leaf_273_clk _00978_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24392_ net7 ser_C.shift_reg\[24\] VGND VGND VPWR VPWR _10666_ sky130_fd_sc_hd__and2_1
XFILLER_123_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26131_ deser_B.serial_word\[86\] deser_B.shift_reg\[86\] net56 VGND VGND VPWR VPWR
+ _03433_ sky130_fd_sc_hd__mux2_1
X_23343_ systolic_inst.A_outs\[0\]\[2\] systolic_inst.B_outs\[0\]\[3\] VGND VGND VPWR
+ VPWR _09971_ sky130_fd_sc_hd__nand2_1
XFILLER_177_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20555_ _07485_ _07486_ VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__and2_1
XFILLER_197_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26062_ deser_B.serial_word\[17\] deser_B.shift_reg\[17\] net55 VGND VGND VPWR VPWR
+ _03364_ sky130_fd_sc_hd__mux2_1
X_23274_ _09910_ _09914_ _09915_ VGND VGND VPWR VPWR _09916_ sky130_fd_sc_hd__a21oi_1
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20486_ _07359_ _07385_ _07384_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__a21boi_1
XFILLER_121_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25013_ C_out\[333\] net97 net80 ser_C.shift_reg\[333\] _10976_ VGND VGND VPWR VPWR
+ _02583_ sky130_fd_sc_hd__a221o_1
X_22225_ _08954_ _08970_ VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22156_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[5\] _08901_ _08902_
+ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_205_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_205_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21107_ _07976_ _07977_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__and2_1
XFILLER_191_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22087_ systolic_inst.B_outs\[1\]\[1\] systolic_inst.B_shift\[1\]\[1\] net122 VGND
+ VGND VPWR VPWR _01787_ sky130_fd_sc_hd__mux2_1
X_26964_ clknet_leaf_22_A_in_serial_clk _00762_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28703_ clknet_leaf_188_clk _02501_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[251\]
+ sky130_fd_sc_hd__dfrtp_1
X_25915_ systolic_inst.acc_wires\[12\]\[7\] C_out\[391\] net18 VGND VGND VPWR VPWR
+ _03217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21038_ _07868_ _07870_ _07909_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__nor3_1
X_29683_ clknet_leaf_106_clk _03478_ net152 VGND VGND VPWR VPWR ser_C.bit_idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_197_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26895_ clknet_leaf_7_A_in_serial_clk _00693_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_143_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_197_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28634_ clknet_leaf_181_clk _02432_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[182\]
+ sky130_fd_sc_hd__dfrtp_1
X_13860_ deser_A.serial_word\[21\] deser_A.shift_reg\[21\] net58 VGND VGND VPWR VPWR
+ _00686_ sky130_fd_sc_hd__mux2_1
X_25846_ systolic_inst.acc_wires\[10\]\[2\] C_out\[322\] net14 VGND VGND VPWR VPWR
+ _03148_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28565_ clknet_leaf_167_clk _02363_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13791_ B_in\[98\] deser_B.word_buffer\[98\] _00005_ VGND VGND VPWR VPWR _00628_
+ sky130_fd_sc_hd__mux2_1
X_22989_ _09627_ _09665_ VGND VGND VPWR VPWR _09666_ sky130_fd_sc_hd__xnor2_1
X_25777_ systolic_inst.acc_wires\[7\]\[29\] C_out\[253\] net43 VGND VGND VPWR VPWR
+ _03079_ sky130_fd_sc_hd__mux2_1
XFILLER_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27516_ clknet_leaf_225_clk _01314_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_15530_ systolic_inst.A_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[2\] systolic_inst.B_outs\[13\]\[6\]
+ systolic_inst.B_outs\[13\]\[7\] VGND VGND VPWR VPWR _12588_ sky130_fd_sc_hd__and4b_1
X_24728_ net113 ser_C.shift_reg\[192\] VGND VGND VPWR VPWR _10834_ sky130_fd_sc_hd__and2_1
XFILLER_63_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28496_ clknet_leaf_117_clk _02294_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_67_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.A_outs\[13\]\[1\] systolic_inst.B_outs\[13\]\[5\]
+ systolic_inst.B_outs\[13\]\[6\] VGND VGND VPWR VPWR _12521_ sky130_fd_sc_hd__and4_1
XFILLER_76_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27447_ clknet_leaf_241_clk _01245_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_190_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_190_clk
+ sky130_fd_sc_hd__clkbuf_8
X_24659_ C_out\[156\] net104 _10643_ ser_C.shift_reg\[156\] _10799_ VGND VGND VPWR
+ VPWR _02406_ sky130_fd_sc_hd__a221o_1
XFILLER_230_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17200_ net107 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[1\] _04461_
+ _04463_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__a22o_1
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14412_ systolic_inst.A_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[5\] systolic_inst.B_outs\[15\]\[6\]
+ systolic_inst.B_outs\[15\]\[7\] VGND VGND VPWR VPWR _11595_ sky130_fd_sc_hd__and4b_1
X_18180_ _05341_ _05313_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__and2b_1
XFILLER_204_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27378_ clknet_leaf_341_clk _01176_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15392_ _12444_ _12453_ _12454_ VGND VGND VPWR VPWR _12455_ sky130_fd_sc_hd__nand3_1
XFILLER_184_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29117_ clknet_leaf_159_clk _02915_ net151 VGND VGND VPWR VPWR C_out\[89\] sky130_fd_sc_hd__dfrtp_1
XFILLER_168_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17131_ _04399_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__nor2_1
X_14343_ systolic_inst.A_outs\[15\]\[4\] systolic_inst.B_outs\[15\]\[5\] VGND VGND
+ VPWR VPWR _11528_ sky130_fd_sc_hd__nand2_1
X_26329_ clknet_leaf_1_A_in_serial_clk _00137_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_204_1178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29048_ clknet_leaf_102_clk _02846_ net151 VGND VGND VPWR VPWR C_out\[20\] sky130_fd_sc_hd__dfrtp_1
X_14274_ _11419_ _11460_ VGND VGND VPWR VPWR _11461_ sky130_fd_sc_hd__or2_1
X_17062_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[11\]\[14\]
+ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__or2_1
XFILLER_195_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16013_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.B_outs\[12\]\[1\] systolic_inst.A_outs\[12\]\[3\]
+ systolic_inst.A_outs\[12\]\[4\] VGND VGND VPWR VPWR _13011_ sky130_fd_sc_hd__and4_1
X_13225_ deser_A.word_buffer\[63\] deser_A.serial_word\[63\] net127 VGND VGND VPWR
+ VPWR _00073_ sky130_fd_sc_hd__mux2_1
XFILLER_152_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13156_ net3 deser_B.receiving VGND VGND VPWR VPWR _11305_ sky130_fd_sc_hd__nor2_1
XFILLER_135_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17964_ _05155_ _05156_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__nor2_1
XFILLER_111_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19703_ _06684_ _06706_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__nand2b_1
X_16915_ _04229_ _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__nor2_1
XFILLER_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17895_ _05088_ _05089_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_105_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19634_ systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[1\] VGND VGND VPWR
+ VPWR _06641_ sky130_fd_sc_hd__nand2_1
XFILLER_38_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16846_ _04057_ _04163_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__or2_1
XFILLER_4_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19565_ _06577_ _06597_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16777_ systolic_inst.B_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[7\] VGND VGND
+ VPWR VPWR _04097_ sky130_fd_sc_hd__nand2_4
X_13989_ deser_B.shift_reg\[23\] deser_B.shift_reg\[24\] net125 VGND VGND VPWR VPWR
+ _00815_ sky130_fd_sc_hd__mux2_1
XFILLER_98_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18516_ _05615_ _05645_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__nand3_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15728_ _12778_ _12779_ VGND VGND VPWR VPWR _12780_ sky130_fd_sc_hd__nor2_1
X_19496_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[7\]\[14\]
+ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__or2_1
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18447_ net108 _05578_ _05579_ _05580_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__o31ai_1
X_15659_ _12576_ _12712_ VGND VGND VPWR VPWR _12713_ sky130_fd_sc_hd__or2_1
XFILLER_221_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_181_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_181_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_146_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18378_ systolic_inst.acc_wires\[9\]\[26\] systolic_inst.acc_wires\[9\]\[27\] systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__o21a_1
XFILLER_105_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17329_ _04546_ _04584_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_135_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20340_ _07254_ _07277_ _07278_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_96_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20271_ _07210_ _07211_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__nand2_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22010_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[21\]
+ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_19_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_241_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_241_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_7_A_in_serial_clk clknet_2_2__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_7_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_130_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23961_ systolic_inst.B_shift\[13\]\[0\] B_in\[40\] _00008_ VGND VGND VPWR VPWR _10506_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25700_ systolic_inst.acc_wires\[5\]\[16\] C_out\[176\] net47 VGND VGND VPWR VPWR
+ _03002_ sky130_fd_sc_hd__mux2_1
XFILLER_111_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22912_ systolic_inst.A_outs\[1\]\[6\] _09590_ _09589_ VGND VGND VPWR VPWR _09591_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_99_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23892_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[31\]
+ VGND VGND VPWR VPWR _10478_ sky130_fd_sc_hd__xnor2_1
X_26680_ clknet_leaf_26_B_in_serial_clk _00483_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25631_ systolic_inst.acc_wires\[3\]\[11\] C_out\[107\] net49 VGND VGND VPWR VPWR
+ _02933_ sky130_fd_sc_hd__mux2_1
X_22843_ _09480_ _09523_ VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_192_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28350_ clknet_leaf_342_clk _02148_ VGND VGND VPWR VPWR systolic_inst.A_shift\[24\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25562_ systolic_inst.acc_wires\[1\]\[6\] C_out\[38\] net36 VGND VGND VPWR VPWR _02864_
+ sky130_fd_sc_hd__mux2_1
X_22774_ systolic_inst.A_outs\[1\]\[2\] systolic_inst.B_outs\[1\]\[3\] systolic_inst.A_outs\[1\]\[3\]
+ systolic_inst.B_outs\[1\]\[4\] VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_49_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27301_ clknet_leaf_290_clk _01099_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24513_ C_out\[83\] net100 net82 ser_C.shift_reg\[83\] _10726_ VGND VGND VPWR VPWR
+ _02333_ sky130_fd_sc_hd__a221o_1
X_21725_ _08530_ _08531_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__nand2_1
XFILLER_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25493_ systolic_inst.cycle_cnt\[20\] _11279_ _11223_ systolic_inst.cycle_cnt\[19\]
+ VGND VGND VPWR VPWR _11226_ sky130_fd_sc_hd__a22oi_1
X_28281_ clknet_leaf_134_clk _02079_ VGND VGND VPWR VPWR systolic_inst.B_shift\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_172_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_172_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_169_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27232_ clknet_leaf_274_clk _01030_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24444_ net114 ser_C.shift_reg\[50\] VGND VGND VPWR VPWR _10692_ sky130_fd_sc_hd__and2_1
X_21656_ _08447_ _08464_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__or2_1
XFILLER_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20607_ _07536_ _07537_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__xnor2_1
X_24375_ C_out\[14\] net104 _10643_ ser_C.shift_reg\[14\] _10657_ VGND VGND VPWR VPWR
+ _02264_ sky130_fd_sc_hd__a221o_1
X_27163_ clknet_leaf_297_clk _00961_ net138 VGND VGND VPWR VPWR systolic_inst.B_outs\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_21587_ _08395_ _08396_ _08365_ _08368_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__o211a_1
XFILLER_197_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26114_ deser_B.serial_word\[69\] deser_B.shift_reg\[69\] _00001_ VGND VGND VPWR
+ VPWR _03416_ sky130_fd_sc_hd__mux2_1
X_23326_ _09952_ _09953_ _09954_ VGND VGND VPWR VPWR _09955_ sky130_fd_sc_hd__and3_1
X_20538_ _07468_ _07469_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__xnor2_1
X_27094_ clknet_leaf_6_B_in_serial_clk _00892_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_186_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_186_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23257_ _09900_ _09901_ VGND VGND VPWR VPWR _09902_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_207_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26045_ deser_B.serial_word\[0\] deser_B.shift_reg\[0\] net55 VGND VGND VPWR VPWR
+ _03347_ sky130_fd_sc_hd__mux2_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20469_ _07402_ _07403_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__nor2_1
XFILLER_84_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22208_ _08918_ _08953_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_234_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23188_ net109 systolic_inst.acc_wires\[1\]\[17\] net65 _09843_ VGND VGND VPWR VPWR
+ _01891_ sky130_fd_sc_hd__a22o_1
XFILLER_238_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_8__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_199_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22139_ _08886_ _08887_ _08870_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__a21oi_1
X_27996_ clknet_leaf_117_clk _01794_ net152 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14961_ systolic_inst.A_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[6\] _11264_ systolic_inst.A_outs\[14\]\[2\]
+ VGND VGND VPWR VPWR _12082_ sky130_fd_sc_hd__o2bb2a_1
X_26947_ clknet_leaf_19_A_in_serial_clk _00745_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16700_ _04020_ _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__nand2_1
XFILLER_236_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13912_ deser_A.serial_word\[73\] deser_A.shift_reg\[73\] net57 VGND VGND VPWR VPWR
+ _00738_ sky130_fd_sc_hd__mux2_1
XFILLER_208_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29666_ clknet_leaf_2_B_in_serial_clk _03461_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17680_ _04912_ _04913_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__or2_1
X_26878_ clknet_leaf_13_A_in_serial_clk _00676_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14892_ _11978_ _12013_ VGND VGND VPWR VPWR _12015_ sky130_fd_sc_hd__and2_1
XFILLER_235_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28617_ clknet_leaf_215_clk _02415_ net149 VGND VGND VPWR VPWR ser_C.shift_reg\[165\]
+ sky130_fd_sc_hd__dfrtp_1
X_16631_ _03948_ _03954_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__and3_1
X_13843_ deser_A.serial_word\[4\] deser_A.shift_reg\[4\] net58 VGND VGND VPWR VPWR
+ _00669_ sky130_fd_sc_hd__mux2_1
X_25829_ systolic_inst.acc_wires\[9\]\[17\] C_out\[305\] net15 VGND VGND VPWR VPWR
+ _03131_ sky130_fd_sc_hd__mux2_1
XFILLER_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29597_ clknet_leaf_14_B_in_serial_clk _03392_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19350_ _06377_ _06380_ _06378_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__o21ba_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28548_ clknet_leaf_178_clk _02346_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_16562_ _03908_ _03909_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__xnor2_1
X_13774_ B_in\[81\] deser_B.word_buffer\[81\] net86 VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18301_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[16\]
+ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_139_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15513_ _12570_ _12571_ VGND VGND VPWR VPWR _12572_ sky130_fd_sc_hd__xor2_1
X_19281_ _06238_ _06342_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__or2_1
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_163_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_163_clk
+ sky130_fd_sc_hd__clkbuf_8
X_28479_ clknet_leaf_110_clk _02277_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_175_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16493_ _03850_ _03851_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__nand2_1
XFILLER_206_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18232_ _05409_ _05410_ _05402_ _05406_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__a211o_1
XFILLER_128_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15444_ _12502_ _12503_ net116 VGND VGND VPWR VPWR _12505_ sky130_fd_sc_hd__o21a_1
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18163_ _05347_ _05348_ _05349_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15375_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[1\]
+ systolic_inst.B_outs\[13\]\[0\] VGND VGND VPWR VPWR _12440_ sky130_fd_sc_hd__a22o_1
XFILLER_106_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17114_ _04405_ _04404_ systolic_inst.acc_wires\[11\]\[21\] net105 VGND VGND VPWR
+ VPWR _01255_ sky130_fd_sc_hd__a2bb2o_1
X_14326_ net118 _11510_ _11511_ VGND VGND VPWR VPWR _11512_ sky130_fd_sc_hd__and3_1
X_18094_ _05243_ _05245_ _05281_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap116 net117 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_130_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap127 net128 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_12
X_17045_ net105 systolic_inst.acc_wires\[11\]\[11\] net69 _04346_ VGND VGND VPWR VPWR
+ _01245_ sky130_fd_sc_hd__a22o_1
X_14257_ _11443_ _11437_ VGND VGND VPWR VPWR _11444_ sky130_fd_sc_hd__and2b_1
Xmax_cap138 net139 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_16
Xmax_cap149 net152 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_16
XFILLER_174_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13208_ deser_A.word_buffer\[46\] deser_A.serial_word\[46\] net127 VGND VGND VPWR
+ VPWR _00056_ sky130_fd_sc_hd__mux2_1
XFILLER_217_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14188_ net107 systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[4\] _11377_
+ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__a21o_1
XFILLER_98_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13139_ systolic_inst.cycle_cnt\[7\] systolic_inst.cycle_cnt\[6\] systolic_inst.cycle_cnt\[5\]
+ systolic_inst.cycle_cnt\[4\] VGND VGND VPWR VPWR _11292_ sky130_fd_sc_hd__or4_1
XFILLER_217_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18996_ _06081_ _06084_ _06083_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__o21a_1
XFILLER_225_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17947_ _05108_ _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__and2b_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17878_ _05050_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__nand2b_1
XFILLER_187_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19617_ systolic_inst.A_outs\[6\]\[5\] systolic_inst.A_outs\[5\]\[5\] net120 VGND
+ VGND VPWR VPWR _01527_ sky130_fd_sc_hd__mux2_1
X_16829_ _04130_ _04147_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__xor2_1
XFILLER_96_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19548_ _06583_ _06582_ systolic_inst.acc_wires\[7\]\[21\] net105 VGND VGND VPWR
+ VPWR _01511_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_234_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_234_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_154_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_154_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19479_ net105 systolic_inst.acc_wires\[7\]\[11\] net62 _06524_ VGND VGND VPWR VPWR
+ _01501_ sky130_fd_sc_hd__a22o_1
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21510_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[3\] _08323_ net122
+ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__mux2_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_230_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22490_ _09223_ VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__inv_2
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21441_ _08262_ _08264_ _08276_ _08277_ _08270_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__a311oi_4
XFILLER_72_1384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24160_ _10581_ systolic_inst.A_shift\[27\]\[3\] net70 VGND VGND VPWR VPWR _02125_
+ sky130_fd_sc_hd__mux2_1
X_21372_ _08218_ _08219_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_B_in_serial_clk clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_14_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_68_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23111_ _09777_ VGND VGND VPWR VPWR _09778_ sky130_fd_sc_hd__inv_2
XFILLER_135_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20323_ _07230_ _07260_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__xor2_1
X_24091_ systolic_inst.B_shift\[23\]\[1\] B_in\[57\] net59 VGND VGND VPWR VPWR _10555_
+ sky130_fd_sc_hd__mux2_1
XFILLER_200_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23042_ _09627_ _09716_ VGND VGND VPWR VPWR _09717_ sky130_fd_sc_hd__nor2_1
XFILLER_66_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_181_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20254_ systolic_inst.A_outs\[5\]\[1\] systolic_inst.B_outs\[5\]\[2\] systolic_inst.B_outs\[5\]\[3\]
+ systolic_inst.A_outs\[5\]\[0\] VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__a22oi_1
XFILLER_235_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_181_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27850_ clknet_leaf_181_clk _01648_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_118_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20185_ _07146_ _07149_ _07151_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__o21ai_1
XFILLER_153_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26801_ clknet_leaf_89_clk _00603_ net5 VGND VGND VPWR VPWR B_in\[73\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27781_ clknet_leaf_186_clk _01579_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24993_ C_out\[323\] net97 net80 ser_C.shift_reg\[323\] _10966_ VGND VGND VPWR VPWR
+ _02573_ sky130_fd_sc_hd__a221o_1
XFILLER_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29520_ clknet_leaf_256_clk _03318_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[492\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_215_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26732_ clknet_leaf_79_clk _00534_ net144 VGND VGND VPWR VPWR B_in\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_229_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23944_ systolic_inst.B_shift\[14\]\[4\] B_in\[20\] net59 VGND VGND VPWR VPWR _10501_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29451_ clknet_leaf_290_clk _03249_ net139 VGND VGND VPWR VPWR C_out\[423\] sky130_fd_sc_hd__dfrtp_1
X_26663_ clknet_leaf_4_B_in_serial_clk _00466_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_179_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23875_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[28\]
+ VGND VGND VPWR VPWR _10464_ sky130_fd_sc_hd__nand2_1
XFILLER_57_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28402_ clknet_leaf_32_clk _02200_ VGND VGND VPWR VPWR systolic_inst.A_shift\[16\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25614_ systolic_inst.acc_wires\[2\]\[26\] C_out\[90\] net51 VGND VGND VPWR VPWR
+ _02916_ sky130_fd_sc_hd__mux2_1
X_22826_ _09505_ _09506_ _09470_ _09472_ VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__o211ai_1
X_29382_ clknet_leaf_245_clk _03180_ net145 VGND VGND VPWR VPWR C_out\[354\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26594_ clknet_leaf_30_A_in_serial_clk _00397_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_1251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28333_ clknet_leaf_342_clk _02131_ VGND VGND VPWR VPWR systolic_inst.A_shift\[26\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25545_ systolic_inst.acc_wires\[0\]\[21\] C_out\[21\] net54 VGND VGND VPWR VPWR
+ _02847_ sky130_fd_sc_hd__mux2_1
XFILLER_13_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22757_ _09416_ _09439_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_145_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21708_ _08443_ _08514_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__nor2_1
X_28264_ clknet_leaf_53_clk _02062_ VGND VGND VPWR VPWR systolic_inst.B_shift\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13490_ deser_A.shift_reg\[54\] deser_A.shift_reg\[55\] net130 VGND VGND VPWR VPWR
+ _00327_ sky130_fd_sc_hd__mux2_1
X_25476_ systolic_inst.cycle_cnt\[14\] _11306_ _11210_ systolic_inst.cycle_cnt\[15\]
+ VGND VGND VPWR VPWR _11214_ sky130_fd_sc_hd__a31o_1
X_22688_ systolic_inst.B_outs\[0\]\[7\] systolic_inst.B_shift\[0\]\[7\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__mux2_1
XFILLER_157_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27215_ clknet_leaf_292_clk _01013_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_24427_ C_out\[40\] _11302_ net81 ser_C.shift_reg\[40\] _10683_ VGND VGND VPWR VPWR
+ _02290_ sky130_fd_sc_hd__a221o_1
X_21639_ systolic_inst.B_outs\[3\]\[3\] systolic_inst.B_outs\[3\]\[4\] systolic_inst.A_outs\[3\]\[4\]
+ systolic_inst.A_outs\[3\]\[5\] VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__and4_1
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28195_ clknet_leaf_56_clk _01993_ VGND VGND VPWR VPWR systolic_inst.B_shift\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15160_ _12262_ _12265_ _12269_ _12270_ VGND VGND VPWR VPWR _12272_ sky130_fd_sc_hd__o211a_1
X_27146_ clknet_leaf_8_clk _00944_ VGND VGND VPWR VPWR systolic_inst.A_shift\[21\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24358_ net7 ser_C.shift_reg\[7\] VGND VGND VPWR VPWR _10649_ sky130_fd_sc_hd__and2_1
XFILLER_165_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14111_ systolic_inst.B_shift\[12\]\[3\] net72 _11333_ B_in\[99\] VGND VGND VPWR
+ VPWR _00933_ sky130_fd_sc_hd__a22o_1
X_23309_ _09925_ _09938_ VGND VGND VPWR VPWR _09939_ sky130_fd_sc_hd__or2_1
XFILLER_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15091_ _12205_ _12206_ VGND VGND VPWR VPWR _12208_ sky130_fd_sc_hd__nor2_1
X_27077_ clknet_leaf_26_B_in_serial_clk _00875_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24289_ systolic_inst.A_shift\[12\]\[0\] A_in\[48\] net59 VGND VGND VPWR VPWR _10618_
+ sky130_fd_sc_hd__mux2_1
XFILLER_141_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14042_ deser_B.shift_reg\[76\] deser_B.shift_reg\[77\] deser_B.receiving VGND VGND
+ VPWR VPWR _00868_ sky130_fd_sc_hd__mux2_1
XFILLER_5_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26028_ systolic_inst.acc_wires\[15\]\[24\] ser_C.parallel_data\[504\] net37 VGND
+ VGND VPWR VPWR _03330_ sky130_fd_sc_hd__mux2_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18850_ _05961_ _05962_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__nand2_1
XFILLER_84_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17801_ net116 systolic_inst.B_outs\[9\]\[0\] systolic_inst.A_outs\[9\]\[0\] VGND
+ VGND VPWR VPWR _05002_ sky130_fd_sc_hd__and3_1
XFILLER_171_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_164_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18781_ _05903_ _05902_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__and2b_1
X_27979_ clknet_leaf_168_clk _01777_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_121_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15993_ _12990_ _12991_ VGND VGND VPWR VPWR _12992_ sky130_fd_sc_hd__or2_1
XFILLER_121_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17732_ _04950_ _04954_ _04957_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__nand3_1
X_14944_ _12065_ _12064_ VGND VGND VPWR VPWR _12066_ sky130_fd_sc_hd__and2b_1
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29649_ clknet_leaf_5_B_in_serial_clk _03444_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_17663_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[10\]\[12\]
+ _04896_ _04898_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__a211o_1
X_14875_ _11992_ _11996_ VGND VGND VPWR VPWR _11998_ sky130_fd_sc_hd__and2_1
XFILLER_63_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19402_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[7\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__a21o_1
XFILLER_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16614_ _03934_ _03939_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__nand2_1
X_13826_ _11320_ _11322_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__nor2_1
X_17594_ _04833_ _04834_ _04832_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__a21bo_1
XFILLER_211_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19333_ _06343_ _06392_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__xor2_1
X_16545_ _03886_ _03888_ _03895_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13757_ B_in\[64\] deser_B.word_buffer\[64\] net87 VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_136_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_206_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19264_ _06308_ _06326_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__xor2_1
XFILLER_149_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16476_ _03807_ _03809_ _03810_ _03815_ _03836_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__o311a_1
X_13688_ deser_B.word_buffer\[124\] deser_B.serial_word\[124\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__mux2_1
X_18215_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[9\]\[4\]
+ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__and2_1
XFILLER_15_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15427_ _12470_ _12487_ VGND VGND VPWR VPWR _12488_ sky130_fd_sc_hd__xor2_1
X_19195_ _06242_ _06259_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__or2_1
XFILLER_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18146_ _05331_ _05332_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__xor2_1
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15358_ systolic_inst.A_outs\[13\]\[2\] systolic_inst.A_outs\[12\]\[2\] net115 VGND
+ VGND VPWR VPWR _01076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14309_ _11492_ _11493_ VGND VGND VPWR VPWR _11495_ sky130_fd_sc_hd__xor2_1
XFILLER_176_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18077_ _05263_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15289_ _12381_ VGND VGND VPWR VPWR _12382_ sky130_fd_sc_hd__inv_2
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17028_ _04327_ _04329_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__nand2_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xload_slew141 net142 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_16
XFILLER_100_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xload_slew152 net5 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_16
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18979_ _06065_ _06067_ _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__a21o_1
XFILLER_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21990_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[18\]
+ VGND VGND VPWR VPWR _08773_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_236_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20941_ _07815_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_236_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23660_ _10278_ _10279_ VGND VGND VPWR VPWR _10280_ sky130_fd_sc_hd__and2_1
X_20872_ _07749_ _07748_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[3\]
+ net108 VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_46_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22611_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[22\]
+ VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_127_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
X_23591_ _10148_ _10151_ _10211_ _10212_ VGND VGND VPWR VPWR _10213_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22542_ _09260_ _09262_ _09258_ VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__a21bo_1
X_25330_ net112 ser_C.shift_reg\[493\] VGND VGND VPWR VPWR _11135_ sky130_fd_sc_hd__and2_1
XFILLER_195_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22473_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[2\]\[1\]
+ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__or2_1
X_25261_ ser_C.parallel_data\[457\] net102 net74 ser_C.shift_reg\[457\] _11100_ VGND
+ VGND VPWR VPWR _02707_ sky130_fd_sc_hd__a221o_1
XFILLER_33_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27000_ clknet_leaf_16_B_in_serial_clk _00798_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_210_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21424_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[25\]
+ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__xor2_2
X_24212_ _10591_ systolic_inst.A_shift\[20\]\[5\] net70 VGND VGND VPWR VPWR _02167_
+ sky130_fd_sc_hd__mux2_1
X_25192_ net111 ser_C.shift_reg\[424\] VGND VGND VPWR VPWR _11066_ sky130_fd_sc_hd__and2_1
X_24143_ systolic_inst.A_shift\[29\]\[3\] A_in\[107\] net59 VGND VGND VPWR VPWR _10573_
+ sky130_fd_sc_hd__mux2_1
X_21355_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[15\]
+ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__and2_1
XFILLER_194_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20306_ _07222_ _07245_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__and2_1
XFILLER_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24074_ systolic_inst.B_shift\[3\]\[1\] net70 net83 systolic_inst.B_shift\[7\]\[1\]
+ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__a22o_1
X_28951_ clknet_leaf_264_clk _02749_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_163_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21286_ _08144_ _08145_ _08137_ _08141_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__a211o_1
XFILLER_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23025_ _09655_ _09669_ _09667_ VGND VGND VPWR VPWR _09701_ sky130_fd_sc_hd__o21a_1
X_27902_ clknet_leaf_41_clk _01700_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20237_ systolic_inst.B_outs\[4\]\[6\] systolic_inst.B_outs\[0\]\[6\] net117 VGND
+ VGND VPWR VPWR _01600_ sky130_fd_sc_hd__mux2_1
XFILLER_131_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28882_ clknet_leaf_330_clk _02680_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[430\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_31_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27833_ clknet_leaf_142_clk _01631_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_162_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20168_ _07137_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__inv_2
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27764_ clknet_leaf_210_clk _01562_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_20099_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[6\]\[13\]
+ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__xor2_1
X_24976_ net111 ser_C.shift_reg\[316\] VGND VGND VPWR VPWR _10958_ sky130_fd_sc_hd__and2_1
XFILLER_183_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29503_ clknet_leaf_266_clk _03301_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[475\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26715_ clknet_leaf_27_B_in_serial_clk _00518_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23927_ _10496_ systolic_inst.B_shift\[18\]\[7\] net71 VGND VGND VPWR VPWR _01977_
+ sky130_fd_sc_hd__mux2_1
X_27695_ clknet_leaf_236_clk _01493_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29434_ clknet_leaf_335_clk _03232_ net131 VGND VGND VPWR VPWR C_out\[406\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26646_ clknet_leaf_18_B_in_serial_clk _00449_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_14660_ net107 systolic_inst.acc_wires\[15\]\[19\] net69 _11818_ VGND VGND VPWR VPWR
+ _00997_ sky130_fd_sc_hd__a22o_1
X_23858_ _10444_ _10446_ _10448_ VGND VGND VPWR VPWR _10450_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13611_ deser_B.word_buffer\[47\] deser_B.serial_word\[47\] net124 VGND VGND VPWR
+ VPWR _00448_ sky130_fd_sc_hd__mux2_1
X_22809_ systolic_inst.A_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\] systolic_inst.B_outs\[1\]\[5\]
+ systolic_inst.A_outs\[1\]\[2\] VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__a22o_1
X_29365_ clknet_leaf_212_clk _03163_ net147 VGND VGND VPWR VPWR C_out\[337\] sky130_fd_sc_hd__dfrtp_1
XFILLER_207_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_118_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_26_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26577_ clknet_leaf_28_A_in_serial_clk _00380_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_14591_ _11755_ _11757_ _11759_ systolic_inst.acc_wires\[15\]\[9\] net105 VGND VGND
+ VPWR VPWR _00987_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23789_ _10389_ _10391_ VGND VGND VPWR VPWR _10392_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_172_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_B_in_serial_clk clknet_2_2__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_9_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_97_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16330_ _03676_ _03678_ _03708_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__or3_1
XFILLER_38_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28316_ clknet_leaf_4_clk _02114_ VGND VGND VPWR VPWR systolic_inst.A_shift\[28\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25528_ systolic_inst.acc_wires\[0\]\[4\] C_out\[4\] net33 VGND VGND VPWR VPWR _02830_
+ sky130_fd_sc_hd__mux2_1
X_13542_ deser_A.shift_reg\[106\] deser_A.shift_reg\[107\] net129 VGND VGND VPWR VPWR
+ _00379_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29296_ clknet_leaf_316_clk _03094_ net137 VGND VGND VPWR VPWR C_out\[268\] sky130_fd_sc_hd__dfrtp_1
XFILLER_213_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28247_ clknet_leaf_80_clk _02045_ VGND VGND VPWR VPWR systolic_inst.B_shift\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16261_ _03603_ _03605_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__a21o_1
X_25459_ systolic_inst.ce_local _11199_ _11202_ VGND VGND VPWR VPWR _11203_ sky130_fd_sc_hd__and3_1
XFILLER_158_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13473_ deser_A.shift_reg\[37\] deser_A.shift_reg\[38\] deser_A.receiving VGND VGND
+ VPWR VPWR _00310_ sky130_fd_sc_hd__mux2_1
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18000_ systolic_inst.B_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[5\] systolic_inst.A_outs\[9\]\[6\]
+ systolic_inst.B_outs\[9\]\[3\] VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__a22oi_1
XFILLER_12_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15212_ _12314_ _12315_ VGND VGND VPWR VPWR _12316_ sky130_fd_sc_hd__and2_1
XFILLER_51_1254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28178_ clknet_leaf_55_clk _01976_ VGND VGND VPWR VPWR systolic_inst.B_shift\[18\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16192_ _03574_ _03575_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__nand2_1
XFILLER_103_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15143_ _12254_ _12257_ VGND VGND VPWR VPWR _12258_ sky130_fd_sc_hd__xnor2_1
X_27129_ clknet_leaf_16_clk _00927_ VGND VGND VPWR VPWR systolic_inst.A_shift\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19951_ _06883_ _06888_ _06916_ _06914_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__a31o_1
XFILLER_138_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15074_ _12143_ _12159_ _12157_ VGND VGND VPWR VPWR _12192_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_166_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14025_ deser_B.shift_reg\[59\] deser_B.shift_reg\[60\] deser_B.receiving VGND VGND
+ VPWR VPWR _00851_ sky130_fd_sc_hd__mux2_1
X_18902_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[15\]
+ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__and2_1
XFILLER_45_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19882_ _06879_ _06880_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__nand2_1
XFILLER_45_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18833_ _05947_ _05948_ _05940_ _05944_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__a211o_1
XFILLER_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18764_ _05885_ _05886_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__nor2_1
XFILLER_23_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15976_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[0\] _12977_
+ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__a21o_1
XFILLER_48_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _04941_ _04942_ _04939_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__o21ai_2
XFILLER_97_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14927_ _12040_ _12048_ VGND VGND VPWR VPWR _12049_ sky130_fd_sc_hd__nand2_1
XFILLER_23_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18695_ _05766_ _05784_ _05783_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__o21a_1
XFILLER_208_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17646_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[10\]\[11\]
+ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__or2_1
XFILLER_184_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14858_ _11951_ _11981_ VGND VGND VPWR VPWR _11982_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13809_ B_in\[116\] deser_B.word_buffer\[116\] net87 VGND VGND VPWR VPWR _00646_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_109_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_189_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17577_ net120 _04824_ _04825_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__a21oi_1
XFILLER_225_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14789_ systolic_inst.A_outs\[14\]\[1\] systolic_inst.B_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[4\]
+ systolic_inst.A_outs\[14\]\[0\] VGND VGND VPWR VPWR _11915_ sky130_fd_sc_hd__a22o_1
XFILLER_223_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19316_ systolic_inst.B_outs\[7\]\[6\] systolic_inst.A_outs\[7\]\[6\] _11261_ systolic_inst.A_outs\[7\]\[5\]
+ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16528_ _03860_ _03867_ _03872_ _03878_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__and4_1
XFILLER_232_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19247_ systolic_inst.B_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[7\]
+ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_119_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16459_ _03814_ _03817_ _03821_ net67 VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__o31a_1
XFILLER_118_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19178_ systolic_inst.B_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[4\]
+ systolic_inst.A_outs\[7\]\[5\] VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__and4_1
XFILLER_121_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18129_ _05315_ _05316_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__nor2_1
XFILLER_145_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21140_ _08008_ _08009_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_225_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_225_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21071_ _07942_ _07941_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__nand2b_1
XFILLER_141_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20022_ net68 _07012_ _07013_ systolic_inst.acc_wires\[6\]\[1\] net106 VGND VGND
+ VPWR VPWR _01555_ sky130_fd_sc_hd__a32o_1
XFILLER_28_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_207_Right_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24830_ net113 ser_C.shift_reg\[243\] VGND VGND VPWR VPWR _10885_ sky130_fd_sc_hd__and2_1
XFILLER_230_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_176_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24761_ C_out\[207\] net99 net79 ser_C.shift_reg\[207\] _10850_ VGND VGND VPWR VPWR
+ _02457_ sky130_fd_sc_hd__a221o_1
X_21973_ _08741_ _08742_ _08757_ VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__and3_1
XFILLER_132_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_348_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_348_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26500_ clknet_leaf_6_A_in_serial_clk _00303_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_23712_ _10322_ _10323_ _10324_ VGND VGND VPWR VPWR _10326_ sky130_fd_sc_hd__and3_1
X_27480_ clknet_leaf_307_clk _01278_ net141 VGND VGND VPWR VPWR systolic_inst.B_outs\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_20924_ _07772_ _07798_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__xnor2_1
XFILLER_242_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24692_ net112 ser_C.shift_reg\[174\] VGND VGND VPWR VPWR _10816_ sky130_fd_sc_hd__and2_1
XFILLER_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26431_ clknet_leaf_0_clk _00238_ net131 VGND VGND VPWR VPWR A_in\[99\] sky130_fd_sc_hd__dfrtp_1
X_23643_ systolic_inst.B_outs\[0\]\[6\] systolic_inst.A_outs\[0\]\[7\] _10193_ VGND
+ VGND VPWR VPWR _10263_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20855_ _07725_ _07733_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__or2_1
XFILLER_230_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29150_ clknet_leaf_174_clk _02948_ net148 VGND VGND VPWR VPWR C_out\[122\] sky130_fd_sc_hd__dfrtp_1
XFILLER_168_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26362_ clknet_leaf_17_clk _00169_ net134 VGND VGND VPWR VPWR A_in\[30\] sky130_fd_sc_hd__dfrtp_1
X_20786_ _07690_ _07689_ systolic_inst.acc_wires\[5\]\[24\] net106 VGND VGND VPWR
+ VPWR _01642_ sky130_fd_sc_hd__a2bb2o_1
X_23574_ systolic_inst.A_outs\[0\]\[5\] _10195_ _10194_ VGND VGND VPWR VPWR _10196_
+ sky130_fd_sc_hd__a21o_1
X_28101_ clknet_leaf_111_clk _01899_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_214_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25313_ ser_C.parallel_data\[483\] net102 net74 ser_C.shift_reg\[483\] _11126_ VGND
+ VGND VPWR VPWR _02733_ sky130_fd_sc_hd__a221o_1
X_29081_ clknet_leaf_109_clk _02879_ net150 VGND VGND VPWR VPWR C_out\[53\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_214_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22525_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[2\]\[8\]
+ _09250_ _09252_ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_214_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26293_ clknet_leaf_2_A_in_serial_clk _00101_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_28032_ clknet_leaf_159_clk _01830_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_155_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_210_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25244_ net111 ser_C.shift_reg\[450\] VGND VGND VPWR VPWR _11092_ sky130_fd_sc_hd__and2_1
X_22456_ _09194_ _09193_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_210_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21407_ _08246_ _08247_ _08248_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__or3_1
X_22387_ systolic_inst.A_outs\[2\]\[5\] systolic_inst.B_outs\[2\]\[6\] systolic_inst.A_outs\[2\]\[6\]
+ systolic_inst.B_outs\[2\]\[7\] VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__and4b_1
XFILLER_182_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25175_ C_out\[414\] net101 net73 ser_C.shift_reg\[414\] _11057_ VGND VGND VPWR VPWR
+ _02664_ sky130_fd_sc_hd__a221o_1
XFILLER_157_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21338_ _11258_ systolic_inst.acc_wires\[4\]\[12\] net63 _08190_ VGND VGND VPWR VPWR
+ _01694_ sky130_fd_sc_hd__a22o_1
XFILLER_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24126_ _10564_ systolic_inst.A_shift\[29\]\[2\] net71 VGND VGND VPWR VPWR _02108_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24057_ systolic_inst.B_shift\[19\]\[0\] B_in\[24\] net59 VGND VGND VPWR VPWR _10546_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28934_ clknet_leaf_264_clk _02732_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[482\]
+ sky130_fd_sc_hd__dfrtp_1
X_21269_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[4\]\[3\]
+ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__and2_1
XFILLER_173_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23008_ net109 _09684_ VGND VGND VPWR VPWR _09685_ sky130_fd_sc_hd__nor2_1
XFILLER_172_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28865_ clknet_leaf_332_clk _02663_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[413\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_237_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_A_in_serial_clk clknet_2_1__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_20_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_27816_ clknet_leaf_143_clk _01614_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15830_ _12853_ _12859_ _12861_ VGND VGND VPWR VPWR _12868_ sky130_fd_sc_hd__o21a_1
XFILLER_103_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28796_ clknet_leaf_233_clk _02594_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[344\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_237_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27747_ clknet_leaf_209_clk _01545_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15761_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[13\]\[2\]
+ VGND VGND VPWR VPWR _12809_ sky130_fd_sc_hd__or2_1
X_24959_ C_out\[306\] net103 net76 ser_C.shift_reg\[306\] _10949_ VGND VGND VPWR VPWR
+ _02556_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_339_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_339_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17500_ _04721_ _04723_ _04752_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__a21o_1
XFILLER_18_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14712_ _11861_ _11862_ VGND VGND VPWR VPWR _11863_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18480_ _05610_ _05611_ systolic_inst.A_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[5\]
+ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__and4bb_1
X_27678_ clknet_leaf_234_clk _01476_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_15692_ net108 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[12\] _12743_
+ _12745_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__a22o_1
XFILLER_79_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29417_ clknet_leaf_333_clk _03215_ net131 VGND VGND VPWR VPWR C_out\[389\] sky130_fd_sc_hd__dfrtp_1
X_17431_ _04683_ _04684_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__xnor2_1
XFILLER_221_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26629_ clknet_leaf_19_B_in_serial_clk _00432_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ net61 _11804_ VGND VGND VPWR VPWR _11805_ sky130_fd_sc_hd__nor2_1
XFILLER_207_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29348_ clknet_leaf_296_clk _03146_ net138 VGND VGND VPWR VPWR C_out\[320\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17362_ _04616_ _04617_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_101_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14574_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[15\]\[7\]
+ VGND VGND VPWR VPWR _11745_ sky130_fd_sc_hd__nand2_1
XFILLER_53_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19101_ systolic_inst.A_outs\[7\]\[4\] _06131_ _06149_ _06148_ _06145_ VGND VGND
+ VPWR VPWR _06168_ sky130_fd_sc_hd__a32o_1
XFILLER_198_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16313_ _03664_ _03691_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13525_ deser_A.shift_reg\[89\] deser_A.shift_reg\[90\] net129 VGND VGND VPWR VPWR
+ _00362_ sky130_fd_sc_hd__mux2_1
X_29279_ clknet_leaf_188_clk _03077_ net148 VGND VGND VPWR VPWR C_out\[251\] sky130_fd_sc_hd__dfrtp_1
X_17293_ _04521_ _04550_ _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__nand3_1
XFILLER_203_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19032_ _06103_ _06101_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[1\]
+ net105 VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__a2bb2o_1
X_16244_ systolic_inst.A_outs\[12\]\[6\] _03594_ _03595_ _03560_ VGND VGND VPWR VPWR
+ _03626_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_174_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13456_ deser_A.shift_reg\[20\] deser_A.shift_reg\[21\] deser_A.receiving VGND VGND
+ VPWR VPWR _00293_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_168_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16175_ _03557_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__or2_1
XFILLER_177_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13387_ A_in\[96\] deser_A.word_buffer\[96\] net96 VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15126_ _12176_ _12219_ _12218_ VGND VGND VPWR VPWR _12242_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19934_ _06930_ _06929_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__nand2b_1
XFILLER_138_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15057_ _12030_ _12173_ VGND VGND VPWR VPWR _12175_ sky130_fd_sc_hd__nand2_1
XFILLER_218_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14008_ deser_B.shift_reg\[42\] deser_B.shift_reg\[43\] net125 VGND VGND VPWR VPWR
+ _00834_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_220_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19865_ _06862_ _06863_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__nor2_1
XFILLER_110_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18816_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[8\]\[3\]
+ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__and2_1
XFILLER_233_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19796_ _06793_ _06796_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_108_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15959_ systolic_inst.A_outs\[12\]\[0\] systolic_inst.A_shift\[24\]\[0\] net115 VGND
+ VGND VPWR VPWR _01138_ sky130_fd_sc_hd__mux2_1
X_18747_ _05870_ _05869_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__nand2b_1
XFILLER_110_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18678_ systolic_inst.B_outs\[8\]\[3\] systolic_inst.B_outs\[8\]\[4\] VGND VGND VPWR
+ VPWR _05804_ sky130_fd_sc_hd__or2_1
XFILLER_224_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_218_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_218_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17629_ _04862_ _04865_ _04868_ net60 VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__a31o_1
XFILLER_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20640_ _07565_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20571_ _07435_ _07501_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22310_ _09051_ _09052_ net122 VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_227_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23290_ _09921_ _09919_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[1\]
+ _11258_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_227_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22241_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] _08985_ VGND
+ VGND VPWR VPWR _08986_ sky130_fd_sc_hd__a21o_1
XFILLER_192_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22172_ _08917_ _08918_ VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__or2_1
XFILLER_191_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21123_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\] _07992_ VGND
+ VGND VPWR VPWR _07993_ sky130_fd_sc_hd__a21o_1
X_26980_ clknet_leaf_28_A_in_serial_clk _00778_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21054_ _07923_ _07925_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__xor2_1
X_25931_ systolic_inst.acc_wires\[12\]\[23\] C_out\[407\] net17 VGND VGND VPWR VPWR
+ _03233_ sky130_fd_sc_hd__mux2_1
XFILLER_160_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20005_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[14\] _06999_ net119
+ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28650_ clknet_leaf_202_clk _02448_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[198\]
+ sky130_fd_sc_hd__dfrtp_1
X_25862_ systolic_inst.acc_wires\[10\]\[18\] C_out\[338\] net11 VGND VGND VPWR VPWR
+ _03164_ sky130_fd_sc_hd__mux2_1
XFILLER_219_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27601_ clknet_leaf_319_clk _01399_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_98_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24813_ C_out\[233\] net99 net79 ser_C.shift_reg\[233\] _10876_ VGND VGND VPWR VPWR
+ _02483_ sky130_fd_sc_hd__a221o_1
XFILLER_80_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28581_ clknet_leaf_311_clk _02379_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[129\]
+ sky130_fd_sc_hd__dfrtp_1
X_25793_ systolic_inst.acc_wires\[8\]\[13\] C_out\[269\] net29 VGND VGND VPWR VPWR
+ _03095_ sky130_fd_sc_hd__mux2_1
XFILLER_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27532_ clknet_leaf_314_clk _01330_ net141 VGND VGND VPWR VPWR systolic_inst.A_outs\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_24744_ net112 ser_C.shift_reg\[200\] VGND VGND VPWR VPWR _10842_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21956_ _08741_ _08742_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_195_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_190_Right_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_195_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_999 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27463_ clknet_leaf_195_clk _01261_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20907_ _07780_ _07781_ _07758_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__a21bo_1
X_24675_ C_out\[164\] net103 net76 ser_C.shift_reg\[164\] _10807_ VGND VGND VPWR VPWR
+ _02414_ sky130_fd_sc_hd__a221o_1
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21887_ _08683_ _08684_ _08676_ _08680_ VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__a211o_1
X_29202_ clknet_leaf_145_clk _03000_ net149 VGND VGND VPWR VPWR C_out\[174\] sky130_fd_sc_hd__dfrtp_1
X_26414_ clknet_leaf_29_clk _00221_ net131 VGND VGND VPWR VPWR A_in\[82\] sky130_fd_sc_hd__dfrtp_1
X_23626_ _10244_ _10245_ _10220_ VGND VGND VPWR VPWR _10247_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_212_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ systolic_inst.B_outs\[3\]\[3\] systolic_inst.B_shift\[3\]\[3\] net120 VGND
+ VGND VPWR VPWR _01661_ sky130_fd_sc_hd__mux2_1
X_27394_ clknet_leaf_335_clk _01192_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29133_ clknet_leaf_169_clk _02931_ net148 VGND VGND VPWR VPWR C_out\[105\] sky130_fd_sc_hd__dfrtp_1
X_26345_ clknet_leaf_23_clk _00152_ net135 VGND VGND VPWR VPWR A_in\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23557_ _10099_ _10102_ _10138_ _10139_ VGND VGND VPWR VPWR _10180_ sky130_fd_sc_hd__o31a_1
XFILLER_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20769_ _07674_ _07675_ _07673_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__o21ai_1
XFILLER_168_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13310_ A_in\[19\] deser_A.word_buffer\[19\] net91 VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__mux2_1
X_29064_ clknet_leaf_114_clk _02862_ net150 VGND VGND VPWR VPWR C_out\[36\] sky130_fd_sc_hd__dfrtp_1
X_22508_ _09232_ _09233_ _09231_ VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_150_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14290_ _11447_ _11449_ _11448_ VGND VGND VPWR VPWR _11476_ sky130_fd_sc_hd__o21bai_1
X_26276_ clknet_leaf_19_A_in_serial_clk _00084_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_210_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23488_ _10066_ _10110_ VGND VGND VPWR VPWR _10112_ sky130_fd_sc_hd__or2_1
XFILLER_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28015_ clknet_leaf_155_clk _01813_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25227_ ser_C.parallel_data\[440\] net101 net73 ser_C.shift_reg\[440\] _11083_ VGND
+ VGND VPWR VPWR _02690_ sky130_fd_sc_hd__a221o_1
X_13241_ deser_A.word_buffer\[79\] deser_A.serial_word\[79\] net127 VGND VGND VPWR
+ VPWR _00089_ sky130_fd_sc_hd__mux2_1
X_22439_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[13\] _09178_ net122
+ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__mux2_1
XFILLER_109_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13172_ deser_A.word_buffer\[10\] deser_A.serial_word\[10\] net128 VGND VGND VPWR
+ VPWR _00020_ sky130_fd_sc_hd__mux2_1
X_25158_ net110 ser_C.shift_reg\[407\] VGND VGND VPWR VPWR _11049_ sky130_fd_sc_hd__and2_1
XFILLER_48_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24109_ systolic_inst.B_shift\[1\]\[4\] _11332_ net83 systolic_inst.B_shift\[5\]\[4\]
+ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__a22o_1
XFILLER_237_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17980_ _05154_ _05171_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__xor2_1
XFILLER_215_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25089_ C_out\[371\] net98 net78 ser_C.shift_reg\[371\] _11014_ VGND VGND VPWR VPWR
+ _02621_ sky130_fd_sc_hd__a221o_1
XFILLER_78_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16931_ _04198_ _04246_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28917_ clknet_leaf_270_clk _02715_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_1006 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19650_ _06643_ _06654_ _06655_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__nand3_1
XFILLER_46_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16862_ _04141_ _04143_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__a21o_1
X_28848_ clknet_leaf_338_clk _02646_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15813_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[13\]\[10\]
+ VGND VGND VPWR VPWR _12853_ sky130_fd_sc_hd__nand2_1
X_18601_ net117 _05727_ _05728_ _05729_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__a31o_1
X_19581_ _06609_ _06611_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28779_ clknet_leaf_230_clk _02577_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[327\]
+ sky130_fd_sc_hd__dfrtp_1
X_16793_ _04066_ _04074_ _04073_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__a21o_1
XFILLER_20_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18532_ _05661_ _05657_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__nand2b_1
X_15744_ _12716_ _12780_ _12778_ VGND VGND VPWR VPWR _12795_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18463_ _05573_ _05576_ _05594_ _05595_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__a211o_1
XFILLER_221_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15675_ _12727_ _12728_ VGND VGND VPWR VPWR _12729_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ net118 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[9\] VGND
+ VGND VPWR VPWR _04670_ sky130_fd_sc_hd__or2_1
XFILLER_21_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14626_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[15\]\[13\]
+ _11784_ VGND VGND VPWR VPWR _11790_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18394_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[30\]
+ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__or2_1
XFILLER_57_1260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[7\]
+ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__o21ai_2
XFILLER_222_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14557_ _11727_ _11728_ _11729_ VGND VGND VPWR VPWR _11731_ sky130_fd_sc_hd__and3_1
XFILLER_159_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_clk clknet_5_24__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13508_ deser_A.shift_reg\[72\] deser_A.shift_reg\[73\] net129 VGND VGND VPWR VPWR
+ _00345_ sky130_fd_sc_hd__mux2_1
X_17276_ _04534_ _04531_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__and2b_1
XFILLER_158_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14488_ _11667_ _11668_ VGND VGND VPWR VPWR _11669_ sky130_fd_sc_hd__nor2_1
XFILLER_179_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload203 clknet_leaf_74_clk VGND VGND VPWR VPWR clkload203/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19015_ systolic_inst.A_outs\[7\]\[4\] systolic_inst.A_outs\[6\]\[4\] net119 VGND
+ VGND VPWR VPWR _01462_ sky130_fd_sc_hd__mux2_1
XFILLER_31_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload214 clknet_leaf_48_clk VGND VGND VPWR VPWR clkload214/X sky130_fd_sc_hd__clkbuf_8
X_16227_ _03607_ _03608_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__xor2_1
Xclkload225 clknet_leaf_135_clk VGND VGND VPWR VPWR clkload225/Y sky130_fd_sc_hd__bufinv_16
X_13439_ deser_A.shift_reg\[3\] deser_A.shift_reg\[4\] deser_A.receiving VGND VGND
+ VPWR VPWR _00276_ sky130_fd_sc_hd__mux2_1
Xclkload236 clknet_leaf_81_clk VGND VGND VPWR VPWR clkload236/Y sky130_fd_sc_hd__clkinv_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload247 clknet_leaf_123_clk VGND VGND VPWR VPWR clkload247/X sky130_fd_sc_hd__clkbuf_8
XFILLER_115_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload258 clknet_leaf_101_clk VGND VGND VPWR VPWR clkload258/Y sky130_fd_sc_hd__inv_6
Xclkload269 clknet_leaf_140_clk VGND VGND VPWR VPWR clkload269/Y sky130_fd_sc_hd__clkinv_2
X_16158_ _03540_ _03541_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__xor2_1
XFILLER_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15109_ _12193_ _12196_ _12225_ VGND VGND VPWR VPWR _12226_ sky130_fd_sc_hd__o21a_1
XFILLER_177_1094 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16089_ _13044_ _13075_ _13077_ VGND VGND VPWR VPWR _13084_ sky130_fd_sc_hd__o21ba_1
XFILLER_103_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19917_ _06877_ _06879_ _06913_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__a21oi_1
XFILLER_218_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19848_ _06808_ _06810_ _06846_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__and3_1
XFILLER_25_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19779_ systolic_inst.B_outs\[6\]\[7\] _06744_ _06745_ VGND VGND VPWR VPWR _06780_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_3_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21810_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[12\] _08614_ net122
+ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__mux2_1
XFILLER_37_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22790_ _09470_ _09471_ _09448_ VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__a21o_1
XFILLER_225_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21741_ _08473_ _08477_ _08507_ _08509_ _08545_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__o311a_1
XFILLER_224_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24460_ net114 ser_C.shift_reg\[58\] VGND VGND VPWR VPWR _10700_ sky130_fd_sc_hd__and2_1
XFILLER_212_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21672_ _08440_ _08446_ _08445_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__a21o_1
XFILLER_240_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23411_ _10035_ _10036_ VGND VGND VPWR VPWR _10037_ sky130_fd_sc_hd__nor2_1
XFILLER_162_1352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20623_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[5\]\[1\]
+ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__nand2_1
X_24391_ C_out\[22\] net104 _10643_ ser_C.shift_reg\[22\] _10665_ VGND VGND VPWR VPWR
+ _02272_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_31_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_123_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26130_ deser_B.serial_word\[85\] deser_B.shift_reg\[85\] net56 VGND VGND VPWR VPWR
+ _03432_ sky130_fd_sc_hd__mux2_1
X_23342_ _09968_ _09969_ VGND VGND VPWR VPWR _09970_ sky130_fd_sc_hd__nand2_1
X_20554_ _07485_ _07486_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__nor2_1
XFILLER_123_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26061_ deser_B.serial_word\[16\] deser_B.shift_reg\[16\] net55 VGND VGND VPWR VPWR
+ _03363_ sky130_fd_sc_hd__mux2_1
XFILLER_164_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23273_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[31\]
+ VGND VGND VPWR VPWR _09915_ sky130_fd_sc_hd__xnor2_1
X_20485_ _07361_ _07418_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25012_ net111 ser_C.shift_reg\[334\] VGND VGND VPWR VPWR _10976_ sky130_fd_sc_hd__and2_1
X_22224_ _08931_ _08967_ VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__xor2_1
XFILLER_121_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22155_ _08901_ _08902_ systolic_inst.A_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[5\]
+ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_5_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21106_ _07937_ _07939_ _07975_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_205_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22086_ systolic_inst.B_outs\[1\]\[0\] systolic_inst.B_shift\[1\]\[0\] net122 VGND
+ VGND VPWR VPWR _01786_ sky130_fd_sc_hd__mux2_1
X_26963_ clknet_leaf_23_A_in_serial_clk _00761_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[96\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_98_clk clknet_5_22__leaf_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
X_28702_ clknet_leaf_188_clk _02500_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[250\]
+ sky130_fd_sc_hd__dfrtp_1
X_25914_ systolic_inst.acc_wires\[12\]\[6\] C_out\[390\] net18 VGND VGND VPWR VPWR
+ _03216_ sky130_fd_sc_hd__mux2_1
X_21037_ _07868_ _07870_ _07909_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__o21a_1
X_29682_ clknet_leaf_106_clk _03477_ net152 VGND VGND VPWR VPWR ser_C.bit_idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_219_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26894_ clknet_leaf_7_A_in_serial_clk _00692_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_197_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28633_ clknet_leaf_181_clk _02431_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[181\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25845_ systolic_inst.acc_wires\[10\]\[1\] C_out\[321\] net14 VGND VGND VPWR VPWR
+ _03147_ sky130_fd_sc_hd__mux2_1
XFILLER_235_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28564_ clknet_leaf_168_clk _02362_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_13790_ B_in\[97\] deser_B.word_buffer\[97\] net89 VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__mux2_1
X_25776_ systolic_inst.acc_wires\[7\]\[28\] C_out\[252\] net44 VGND VGND VPWR VPWR
+ _03078_ sky130_fd_sc_hd__mux2_1
X_22988_ _09662_ _09663_ VGND VGND VPWR VPWR _09665_ sky130_fd_sc_hd__xnor2_1
XFILLER_210_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27515_ clknet_leaf_225_clk _01313_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24727_ C_out\[190\] net99 net79 ser_C.shift_reg\[190\] _10833_ VGND VGND VPWR VPWR
+ _02440_ sky130_fd_sc_hd__a221o_1
XFILLER_215_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28495_ clknet_leaf_117_clk _02293_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_21939_ _08718_ _08724_ _08728_ VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__a21o_1
XFILLER_231_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15460_ systolic_inst.A_outs\[13\]\[1\] systolic_inst.B_outs\[13\]\[6\] VGND VGND
+ VPWR VPWR _12520_ sky130_fd_sc_hd__nand2_1
X_27446_ clknet_leaf_241_clk _01244_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_230_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24658_ net7 ser_C.shift_reg\[157\] VGND VGND VPWR VPWR _10799_ sky130_fd_sc_hd__and2_1
XFILLER_54_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14411_ systolic_inst.B_outs\[15\]\[5\] systolic_inst.A_outs\[15\]\[6\] VGND VGND
+ VPWR VPWR _11594_ sky130_fd_sc_hd__nand2_1
XFILLER_70_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23609_ _11268_ systolic_inst.B_outs\[0\]\[7\] _10120_ VGND VGND VPWR VPWR _10230_
+ sky130_fd_sc_hd__and3_1
X_27377_ clknet_leaf_333_clk _01175_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_15391_ systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[3\]
+ systolic_inst.B_outs\[13\]\[0\] VGND VGND VPWR VPWR _12454_ sky130_fd_sc_hd__a22o_1
X_24589_ C_out\[121\] net100 net82 ser_C.shift_reg\[121\] _10764_ VGND VGND VPWR VPWR
+ _02371_ sky130_fd_sc_hd__a221o_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
X_29116_ clknet_leaf_159_clk _02914_ net151 VGND VGND VPWR VPWR C_out\[88\] sky130_fd_sc_hd__dfrtp_1
XFILLER_204_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17130_ systolic_inst.acc_wires\[11\]\[20\] systolic_inst.acc_wires\[11\]\[21\] systolic_inst.acc_wires\[11\]\[22\]
+ systolic_inst.acc_wires\[11\]\[23\] systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__o41a_1
X_14342_ _11447_ _11526_ VGND VGND VPWR VPWR _11527_ sky130_fd_sc_hd__xnor2_1
X_26328_ clknet_leaf_0_A_in_serial_clk _00136_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_29047_ clknet_leaf_102_clk _02845_ net151 VGND VGND VPWR VPWR C_out\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17061_ _04356_ _04358_ _04360_ systolic_inst.acc_wires\[11\]\[13\] net105 VGND VGND
+ VPWR VPWR _01247_ sky130_fd_sc_hd__a32o_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14273_ _11451_ _11459_ VGND VGND VPWR VPWR _11460_ sky130_fd_sc_hd__xnor2_1
X_26259_ clknet_leaf_6_A_in_serial_clk _00067_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_171_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16012_ systolic_inst.B_outs\[12\]\[0\] systolic_inst.A_outs\[12\]\[4\] VGND VGND
+ VPWR VPWR _13010_ sky130_fd_sc_hd__nand2_1
X_13224_ deser_A.word_buffer\[62\] deser_A.serial_word\[62\] net128 VGND VGND VPWR
+ VPWR _00072_ sky130_fd_sc_hd__mux2_1
XFILLER_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13155_ deser_A.serial_toggle_sync2 deser_A.serial_toggle_sync1 VGND VGND VPWR VPWR
+ _00003_ sky130_fd_sc_hd__xor2_4
XFILLER_139_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17963_ systolic_inst.B_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[5\]
+ systolic_inst.B_outs\[9\]\[3\] VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__a22oi_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_89_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
X_19702_ _06704_ _06705_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__and2_1
XFILLER_111_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16914_ _04227_ _04228_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__nor2_1
XFILLER_211_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17894_ systolic_inst.B_outs\[9\]\[3\] systolic_inst.A_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\]
+ systolic_inst.A_outs\[9\]\[2\] VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_105_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19633_ _06640_ _06638_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[1\]
+ net106 VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_238_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16845_ systolic_inst.A_outs\[11\]\[6\] _04132_ _04133_ _04097_ VGND VGND VPWR VPWR
+ _04163_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_225_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19564_ systolic_inst.acc_wires\[7\]\[20\] systolic_inst.acc_wires\[7\]\[21\] systolic_inst.acc_wires\[7\]\[22\]
+ systolic_inst.acc_wires\[7\]\[23\] systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__o41a_1
X_16776_ _04094_ _04095_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__or2_1
XFILLER_98_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13988_ deser_B.shift_reg\[22\] deser_B.shift_reg\[23\] net125 VGND VGND VPWR VPWR
+ _00814_ sky130_fd_sc_hd__mux2_1
XFILLER_19_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15727_ _12751_ _12754_ _12777_ VGND VGND VPWR VPWR _12779_ sky130_fd_sc_hd__and3_1
X_18515_ _05643_ _05644_ _05632_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__o21bai_1
XFILLER_80_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19495_ net62 _06535_ _06538_ systolic_inst.acc_wires\[7\]\[13\] net105 VGND VGND
+ VPWR VPWR _01503_ sky130_fd_sc_hd__a32o_1
XFILLER_146_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15658_ systolic_inst.B_outs\[13\]\[2\] systolic_inst.A_outs\[13\]\[7\] _12685_ _12648_
+ VGND VGND VPWR VPWR _12712_ sky130_fd_sc_hd__a31o_1
X_18446_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[3\] VGND
+ VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nand2_1
XFILLER_59_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_B_in_serial_clk clknet_2_1__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_22_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_34_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14609_ _11760_ _11766_ _11768_ VGND VGND VPWR VPWR _11775_ sky130_fd_sc_hd__o21a_1
X_18377_ _05527_ _05531_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__nor2_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15589_ _12577_ _12643_ VGND VGND VPWR VPWR _12645_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_13_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_202_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17328_ _04546_ _04584_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__and2_1
XFILLER_239_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17259_ _04516_ _04517_ systolic_inst.A_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[5\]
+ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_96_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20270_ systolic_inst.A_outs\[5\]\[1\] systolic_inst.B_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\]
+ systolic_inst.A_outs\[5\]\[0\] VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__a22o_1
XFILLER_66_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_219_Left_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_241_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_241_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_241_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23960_ systolic_inst.B_shift\[11\]\[7\] _11332_ net83 systolic_inst.B_shift\[15\]\[7\]
+ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__a22o_1
XFILLER_124_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_200_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22911_ systolic_inst.B_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[7\]
+ VGND VGND VPWR VPWR _09590_ sky130_fd_sc_hd__and3_1
XFILLER_217_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23891_ net64 _10476_ _10477_ systolic_inst.acc_wires\[0\]\[30\] _11258_ VGND VGND
+ VPWR VPWR _01960_ sky130_fd_sc_hd__a32o_1
X_25630_ systolic_inst.acc_wires\[3\]\[10\] C_out\[106\] net48 VGND VGND VPWR VPWR
+ _02932_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22842_ _09521_ _09522_ VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_192_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_228_Left_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25561_ systolic_inst.acc_wires\[1\]\[5\] C_out\[37\] net36 VGND VGND VPWR VPWR _02863_
+ sky130_fd_sc_hd__mux2_1
XFILLER_227_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22773_ _09424_ _09454_ VGND VGND VPWR VPWR _09456_ sky130_fd_sc_hd__xor2_1
XFILLER_140_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27300_ clknet_leaf_290_clk _01098_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24512_ net112 ser_C.shift_reg\[84\] VGND VGND VPWR VPWR _10726_ sky130_fd_sc_hd__and2_1
X_21724_ _08521_ _08529_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__or2_1
X_28280_ clknet_leaf_134_clk _02078_ VGND VGND VPWR VPWR systolic_inst.B_shift\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25492_ systolic_inst.cycle_cnt\[20\] systolic_inst.cycle_cnt\[19\] _11223_ VGND
+ VGND VPWR VPWR _11225_ sky130_fd_sc_hd__and3_1
XFILLER_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27231_ clknet_leaf_274_clk _01029_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_24443_ C_out\[48\] _11302_ net81 ser_C.shift_reg\[48\] _10691_ VGND VGND VPWR VPWR
+ _02298_ sky130_fd_sc_hd__a221o_1
XFILLER_71_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21655_ _08462_ _08463_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20606_ _07323_ _07461_ _07512_ _07510_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__a31o_1
XFILLER_123_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27162_ clknet_leaf_297_clk _00960_ net138 VGND VGND VPWR VPWR systolic_inst.B_outs\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_24374_ net7 ser_C.shift_reg\[15\] VGND VGND VPWR VPWR _10657_ sky130_fd_sc_hd__and2_1
XFILLER_165_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21586_ _08365_ _08368_ _08395_ _08396_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__a211oi_2
XFILLER_162_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26113_ deser_B.serial_word\[68\] deser_B.shift_reg\[68\] _00001_ VGND VGND VPWR
+ VPWR _03415_ sky130_fd_sc_hd__mux2_1
XFILLER_137_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23325_ systolic_inst.A_outs\[0\]\[0\] systolic_inst.B_outs\[0\]\[3\] _09933_ _09932_
+ VGND VGND VPWR VPWR _09954_ sky130_fd_sc_hd__a31o_1
XFILLER_123_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27093_ clknet_leaf_5_B_in_serial_clk _00891_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20537_ systolic_inst.B_outs\[5\]\[5\] systolic_inst.A_outs\[5\]\[7\] _07468_ VGND
+ VGND VPWR VPWR _07470_ sky130_fd_sc_hd__and3_1
XFILLER_197_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_186_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26044_ net9 ser_C.shift_reg\[0\] net114 VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_237_Left_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23256_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[28\]
+ VGND VGND VPWR VPWR _09901_ sky130_fd_sc_hd__nand2_1
X_20468_ systolic_inst.A_outs\[5\]\[4\] systolic_inst.B_outs\[5\]\[6\] _11276_ systolic_inst.A_outs\[5\]\[3\]
+ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_207_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22207_ _08947_ _08951_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__xnor2_1
X_23187_ _09840_ _09842_ VGND VGND VPWR VPWR _09843_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20399_ _07333_ _07334_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__xnor2_1
XFILLER_234_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_145_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22138_ _08884_ _08885_ _08864_ _08867_ VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_199_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27995_ clknet_leaf_127_clk _01793_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14960_ systolic_inst.A_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[3\] systolic_inst.B_outs\[14\]\[6\]
+ systolic_inst.B_outs\[14\]\[7\] VGND VGND VPWR VPWR _12081_ sky130_fd_sc_hd__and4b_1
X_26946_ clknet_leaf_19_A_in_serial_clk _00744_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_22069_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[30\]
+ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_141_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13911_ deser_A.serial_word\[72\] deser_A.shift_reg\[72\] net57 VGND VGND VPWR VPWR
+ _00737_ sky130_fd_sc_hd__mux2_1
XFILLER_102_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29665_ clknet_leaf_3_B_in_serial_clk _03460_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_26877_ clknet_leaf_13_A_in_serial_clk _00675_ net144 VGND VGND VPWR VPWR deser_A.serial_word\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14891_ _11978_ _12013_ VGND VGND VPWR VPWR _12014_ sky130_fd_sc_hd__or2_1
XFILLER_74_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16630_ _03935_ _03952_ _03953_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__or3_1
X_13842_ deser_A.serial_word\[3\] deser_A.shift_reg\[3\] net58 VGND VGND VPWR VPWR
+ _00668_ sky130_fd_sc_hd__mux2_1
X_28616_ clknet_leaf_216_clk _02414_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[164\]
+ sky130_fd_sc_hd__dfrtp_1
X_25828_ systolic_inst.acc_wires\[9\]\[16\] C_out\[304\] net15 VGND VGND VPWR VPWR
+ _03130_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29596_ clknet_leaf_14_B_in_serial_clk _03391_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16561_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[28\]
+ _03906_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__a21oi_1
X_28547_ clknet_leaf_165_clk _02345_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_13773_ B_in\[80\] deser_B.word_buffer\[80\] net86 VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__mux2_1
X_25759_ systolic_inst.acc_wires\[7\]\[11\] C_out\[235\] net42 VGND VGND VPWR VPWR
+ _03061_ sky130_fd_sc_hd__mux2_1
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18300_ _05467_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__and2_1
X_15512_ _12502_ _12503_ _12535_ _12533_ VGND VGND VPWR VPWR _12571_ sky130_fd_sc_hd__a31o_1
X_19280_ systolic_inst.A_outs\[7\]\[6\] _06310_ _06311_ _06277_ VGND VGND VPWR VPWR
+ _06342_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_139_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28478_ clknet_leaf_110_clk _02276_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_203_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16492_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[18\]
+ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_175_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18231_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[9\]\[6\]
+ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__or2_1
X_15443_ _12502_ _12503_ VGND VGND VPWR VPWR _12504_ sky130_fd_sc_hd__nand2_1
X_27429_ clknet_leaf_242_clk _01227_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_176_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18162_ _11263_ systolic_inst.A_outs\[9\]\[7\] _05296_ _05320_ VGND VGND VPWR VPWR
+ _05349_ sky130_fd_sc_hd__o211a_1
X_15374_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.A_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\]
+ systolic_inst.A_outs\[13\]\[1\] VGND VGND VPWR VPWR _12439_ sky130_fd_sc_hd__and4_1
XFILLER_184_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17113_ _04395_ _04401_ _04402_ net60 VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__a31o_1
XFILLER_7_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14325_ _11470_ _11472_ _11509_ VGND VGND VPWR VPWR _11511_ sky130_fd_sc_hd__or3_1
X_18093_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__inv_2
XFILLER_157_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap117 net121 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_130_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17044_ _04344_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_130_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14256_ _11441_ _11442_ VGND VGND VPWR VPWR _11443_ sky130_fd_sc_hd__or2_1
XFILLER_172_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap128 deser_A.serial_word_ready VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_12
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap139 net140 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_91_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13207_ deser_A.word_buffer\[45\] deser_A.serial_word\[45\] net127 VGND VGND VPWR
+ VPWR _00055_ sky130_fd_sc_hd__mux2_1
XFILLER_171_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14187_ _11376_ _11375_ VGND VGND VPWR VPWR _11377_ sky130_fd_sc_hd__and2b_1
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13138_ systolic_inst.cycle_cnt\[15\] systolic_inst.cycle_cnt\[14\] systolic_inst.cycle_cnt\[13\]
+ systolic_inst.cycle_cnt\[12\] VGND VGND VPWR VPWR _11291_ sky130_fd_sc_hd__or4_1
XFILLER_135_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18995_ _06086_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__inv_2
XFILLER_174_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17946_ _05109_ _05138_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17877_ _05071_ _05072_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__and2_1
XFILLER_187_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19616_ systolic_inst.A_outs\[6\]\[4\] systolic_inst.A_outs\[5\]\[4\] net120 VGND
+ VGND VPWR VPWR _01526_ sky130_fd_sc_hd__mux2_1
X_16828_ _04145_ _04146_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__nand2_1
XFILLER_241_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19547_ _06573_ _06579_ _06580_ net60 VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_85_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16759_ _04026_ _04041_ _04040_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__o21a_1
XFILLER_185_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_234_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_234_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19478_ _06522_ _06523_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18429_ _05561_ _05562_ _05557_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_44_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21440_ systolic_inst.acc_wires\[4\]\[26\] systolic_inst.acc_wires\[4\]\[27\] systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__o21a_1
XFILLER_147_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_86_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21371_ _08211_ _08214_ _08213_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__o21a_1
XFILLER_120_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23110_ _09773_ _09774_ _09775_ VGND VGND VPWR VPWR _09777_ sky130_fd_sc_hd__and3_1
XFILLER_200_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20322_ _07230_ _07260_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__nand2_1
XFILLER_194_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24090_ _10554_ systolic_inst.B_shift\[19\]\[0\] net71 VGND VGND VPWR VPWR _02082_
+ sky130_fd_sc_hd__mux2_1
XFILLER_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23041_ systolic_inst.B_outs\[1\]\[5\] systolic_inst.B_outs\[1\]\[6\] systolic_inst.A_outs\[1\]\[7\]
+ _09715_ VGND VGND VPWR VPWR _09716_ sky130_fd_sc_hd__a31o_1
X_20253_ net116 _07194_ _07195_ _07188_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_181_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20184_ _07146_ _07149_ _07151_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_38_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26800_ clknet_leaf_88_clk _00602_ net153 VGND VGND VPWR VPWR B_in\[72\] sky130_fd_sc_hd__dfrtp_1
XFILLER_192_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27780_ clknet_leaf_186_clk _01578_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24992_ net111 ser_C.shift_reg\[324\] VGND VGND VPWR VPWR _10966_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_95_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26731_ clknet_leaf_78_clk _00533_ net144 VGND VGND VPWR VPWR B_in\[3\] sky130_fd_sc_hd__dfrtp_1
X_23943_ _10500_ systolic_inst.B_shift\[10\]\[3\] _11332_ VGND VGND VPWR VPWR _01989_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29450_ clknet_leaf_293_clk _03248_ net139 VGND VGND VPWR VPWR C_out\[422\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_179_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26662_ clknet_leaf_2_B_in_serial_clk _00465_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_23874_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[28\]
+ VGND VGND VPWR VPWR _10463_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_179_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25613_ systolic_inst.acc_wires\[2\]\[25\] C_out\[89\] net51 VGND VGND VPWR VPWR
+ _02915_ sky130_fd_sc_hd__mux2_1
X_28401_ clknet_leaf_32_clk _02199_ VGND VGND VPWR VPWR systolic_inst.A_shift\[16\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_22825_ _09470_ _09472_ _09505_ _09506_ VGND VGND VPWR VPWR _09507_ sky130_fd_sc_hd__a211oi_1
X_29381_ clknet_leaf_247_clk _03179_ net145 VGND VGND VPWR VPWR C_out\[353\] sky130_fd_sc_hd__dfrtp_1
XFILLER_226_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26593_ clknet_leaf_30_A_in_serial_clk _00396_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28332_ clknet_leaf_3_clk _02130_ VGND VGND VPWR VPWR systolic_inst.A_shift\[26\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25544_ systolic_inst.acc_wires\[0\]\[20\] C_out\[20\] net54 VGND VGND VPWR VPWR
+ _02846_ sky130_fd_sc_hd__mux2_1
XFILLER_241_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22756_ _09416_ _09439_ VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__and2_1
XFILLER_13_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21707_ _08485_ _08486_ _08487_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__o21ba_1
X_28263_ clknet_leaf_53_clk _02061_ VGND VGND VPWR VPWR systolic_inst.B_shift\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25475_ _11211_ _11212_ systolic_inst.cycle_cnt\[14\] VGND VGND VPWR VPWR _02808_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22687_ systolic_inst.B_outs\[0\]\[6\] systolic_inst.B_shift\[0\]\[6\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__mux2_1
XFILLER_200_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27214_ clknet_leaf_294_clk _01012_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_24426_ net114 ser_C.shift_reg\[41\] VGND VGND VPWR VPWR _10683_ sky130_fd_sc_hd__and2_1
X_21638_ _08440_ _08446_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__xnor2_1
X_28194_ clknet_leaf_49_clk _01992_ VGND VGND VPWR VPWR systolic_inst.B_shift\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27145_ clknet_leaf_7_clk _00943_ VGND VGND VPWR VPWR systolic_inst.A_shift\[21\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_24357_ C_out\[5\] net104 _10643_ ser_C.shift_reg\[5\] _10648_ VGND VGND VPWR VPWR
+ _02255_ sky130_fd_sc_hd__a221o_1
X_21569_ _08378_ _08379_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__or2_1
XFILLER_197_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14110_ systolic_inst.B_shift\[12\]\[2\] net72 _11333_ B_in\[98\] VGND VGND VPWR
+ VPWR _00932_ sky130_fd_sc_hd__a22o_1
X_23308_ _09935_ _09936_ VGND VGND VPWR VPWR _09938_ sky130_fd_sc_hd__xor2_1
X_27076_ clknet_leaf_26_B_in_serial_clk _00874_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_15090_ _12205_ _12206_ VGND VGND VPWR VPWR _12207_ sky130_fd_sc_hd__and2_1
X_24288_ _10617_ systolic_inst.B_shift\[23\]\[7\] net72 VGND VGND VPWR VPWR _02217_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14041_ deser_B.shift_reg\[75\] deser_B.shift_reg\[76\] deser_B.receiving VGND VGND
+ VPWR VPWR _00867_ sky130_fd_sc_hd__mux2_1
X_26027_ systolic_inst.acc_wires\[15\]\[23\] ser_C.parallel_data\[503\] net37 VGND
+ VGND VPWR VPWR _03329_ sky130_fd_sc_hd__mux2_1
XFILLER_107_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23239_ _09881_ _09883_ _09885_ VGND VGND VPWR VPWR _09887_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17800_ systolic_inst.B_outs\[8\]\[7\] systolic_inst.B_outs\[4\]\[7\] net121 VGND
+ VGND VPWR VPWR _01345_ sky130_fd_sc_hd__mux2_1
XFILLER_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ systolic_inst.A_outs\[12\]\[0\] systolic_inst.A_outs\[12\]\[1\] systolic_inst.B_outs\[12\]\[2\]
+ systolic_inst.B_outs\[12\]\[3\] VGND VGND VPWR VPWR _12991_ sky130_fd_sc_hd__and4_1
X_18780_ _05835_ _05878_ _05877_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__o21a_1
X_27978_ clknet_leaf_165_clk _01776_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14943_ _12023_ _12025_ VGND VGND VPWR VPWR _12065_ sky130_fd_sc_hd__and2_1
X_17731_ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__inv_2
X_26929_ clknet_leaf_5_A_in_serial_clk _00727_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29648_ clknet_leaf_1_B_in_serial_clk _03443_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14874_ _11992_ _11996_ VGND VGND VPWR VPWR _11997_ sky130_fd_sc_hd__nor2_1
X_17662_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[10\]\[13\]
+ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__xor2_1
XFILLER_85_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19401_ net105 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] _06451_
+ _06458_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13825_ deser_B.bit_idx\[1\] _11319_ _11321_ VGND VGND VPWR VPWR _11322_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16613_ _03937_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__and2_1
XFILLER_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17593_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[10\]\[3\]
+ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__or2_1
X_29579_ clknet_leaf_23_B_in_serial_clk _03374_ net137 VGND VGND VPWR VPWR deser_B.serial_word\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19332_ _06343_ _06392_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__and2b_1
X_16544_ systolic_inst.acc_wires\[12\]\[24\] systolic_inst.acc_wires\[12\]\[25\] systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__o21a_1
XFILLER_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13756_ B_in\[63\] deser_B.word_buffer\[63\] net87 VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__mux2_1
XFILLER_71_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19263_ _06323_ _06324_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__xor2_1
XFILLER_143_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16475_ _03821_ _03834_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__and2_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13687_ deser_B.word_buffer\[123\] deser_B.serial_word\[123\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15426_ _12483_ _12486_ VGND VGND VPWR VPWR _12487_ sky130_fd_sc_hd__xor2_1
X_18214_ net66 _05393_ _05395_ systolic_inst.acc_wires\[9\]\[3\] net107 VGND VGND
+ VPWR VPWR _01365_ sky130_fd_sc_hd__a32o_1
X_19194_ _06257_ _06258_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15357_ systolic_inst.A_outs\[13\]\[1\] systolic_inst.A_outs\[12\]\[1\] net115 VGND
+ VGND VPWR VPWR _01075_ sky130_fd_sc_hd__mux2_1
X_18145_ _05331_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__nand2b_1
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14308_ _11492_ _11493_ VGND VGND VPWR VPWR _11494_ sky130_fd_sc_hd__and2_1
XFILLER_129_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18076_ _05264_ _05265_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__nor2_1
X_15288_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[21\]
+ VGND VGND VPWR VPWR _12381_ sky130_fd_sc_hd__xnor2_2
XFILLER_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17027_ _04326_ _04329_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_242_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14239_ _11423_ _11424_ _11395_ VGND VGND VPWR VPWR _11427_ sky130_fd_sc_hd__a21o_1
XFILLER_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xload_slew142 net144 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18978_ systolic_inst.acc_wires\[8\]\[24\] systolic_inst.acc_wires\[8\]\[25\] systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__o21a_1
XFILLER_100_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _05119_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20940_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[6\] systolic_inst.B_outs\[4\]\[6\]
+ systolic_inst.A_outs\[4\]\[0\] VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_236_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_236_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20871_ _07735_ _07747_ net117 VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__o21ai_1
XFILLER_241_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22610_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[22\]
+ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__or2_1
XFILLER_228_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23590_ _10167_ _10170_ _10210_ VGND VGND VPWR VPWR _10212_ sky130_fd_sc_hd__nor3_1
XFILLER_35_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22541_ _09265_ _09266_ VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__nand2_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_224_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25260_ net111 ser_C.shift_reg\[458\] VGND VGND VPWR VPWR _11100_ sky130_fd_sc_hd__and2_1
X_22472_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[2\]\[1\]
+ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__nand2_1
XFILLER_33_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24211_ systolic_inst.A_shift\[21\]\[5\] A_in\[85\] net59 VGND VGND VPWR VPWR _10591_
+ sky130_fd_sc_hd__mux2_1
X_21423_ _08263_ _08262_ systolic_inst.acc_wires\[4\]\[24\] _11258_ VGND VGND VPWR
+ VPWR _01706_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25191_ C_out\[422\] net102 net74 ser_C.shift_reg\[422\] _11065_ VGND VGND VPWR VPWR
+ _02672_ sky130_fd_sc_hd__a221o_1
XFILLER_108_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24142_ _10572_ systolic_inst.A_shift\[28\]\[2\] net70 VGND VGND VPWR VPWR _02116_
+ sky130_fd_sc_hd__mux2_1
X_21354_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[15\]
+ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__nor2_1
XFILLER_120_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20305_ _07233_ _07243_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__xor2_1
XFILLER_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24073_ systolic_inst.B_shift\[3\]\[0\] net70 net83 systolic_inst.B_shift\[7\]\[0\]
+ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__a22o_1
X_28950_ clknet_leaf_261_clk _02748_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[498\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21285_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[4\]\[5\]
+ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__or2_1
XFILLER_239_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23024_ _09656_ _09699_ VGND VGND VPWR VPWR _09700_ sky130_fd_sc_hd__xnor2_1
X_27901_ clknet_leaf_42_clk _01699_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20236_ systolic_inst.B_outs\[4\]\[5\] systolic_inst.B_outs\[0\]\[5\] net117 VGND
+ VGND VPWR VPWR _01599_ sky130_fd_sc_hd__mux2_1
XFILLER_235_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28881_ clknet_leaf_288_clk _02679_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[429\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20167_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[23\]
+ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__xor2_1
X_27832_ clknet_leaf_142_clk _01630_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20098_ net106 systolic_inst.acc_wires\[6\]\[12\] net68 _07078_ VGND VGND VPWR VPWR
+ _01566_ sky130_fd_sc_hd__a22o_1
X_27763_ clknet_leaf_211_clk _01561_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24975_ C_out\[314\] net103 net76 ser_C.shift_reg\[314\] _10957_ VGND VGND VPWR VPWR
+ _02564_ sky130_fd_sc_hd__a221o_1
XFILLER_44_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29502_ clknet_leaf_267_clk _03300_ net138 VGND VGND VPWR VPWR ser_C.parallel_data\[474\]
+ sky130_fd_sc_hd__dfrtp_1
X_26714_ clknet_leaf_27_B_in_serial_clk _00517_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_23926_ systolic_inst.B_shift\[22\]\[7\] B_in\[87\] net59 VGND VGND VPWR VPWR _10496_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27694_ clknet_leaf_234_clk _01492_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26645_ clknet_leaf_16_B_in_serial_clk _00448_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_29433_ clknet_leaf_336_clk _03231_ net131 VGND VGND VPWR VPWR C_out\[405\] sky130_fd_sc_hd__dfrtp_1
X_23857_ _10444_ _10446_ _10448_ VGND VGND VPWR VPWR _10449_ sky130_fd_sc_hd__or3_1
XFILLER_166_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13610_ deser_B.word_buffer\[46\] deser_B.serial_word\[46\] net124 VGND VGND VPWR
+ VPWR _00447_ sky130_fd_sc_hd__mux2_1
X_22808_ systolic_inst.A_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\]
+ systolic_inst.B_outs\[1\]\[5\] VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__and4_1
XFILLER_77_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29364_ clknet_leaf_225_clk _03162_ net147 VGND VGND VPWR VPWR C_out\[336\] sky130_fd_sc_hd__dfrtp_1
X_26576_ clknet_leaf_24_A_in_serial_clk _00379_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_14590_ net61 _11758_ VGND VGND VPWR VPWR _11759_ sky130_fd_sc_hd__nor2_1
XFILLER_60_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23788_ _10384_ _10390_ VGND VGND VPWR VPWR _10391_ sky130_fd_sc_hd__nand2_1
XFILLER_198_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_172_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25527_ systolic_inst.acc_wires\[0\]\[3\] C_out\[3\] net33 VGND VGND VPWR VPWR _02829_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13541_ deser_A.shift_reg\[105\] deser_A.shift_reg\[106\] net129 VGND VGND VPWR VPWR
+ _00378_ sky130_fd_sc_hd__mux2_1
X_28315_ clknet_leaf_11_clk _02113_ VGND VGND VPWR VPWR systolic_inst.A_shift\[29\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22739_ systolic_inst.B_outs\[1\]\[1\] systolic_inst.A_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[5\]
+ systolic_inst.B_outs\[1\]\[0\] VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__a22oi_1
X_29295_ clknet_leaf_316_clk _03093_ net137 VGND VGND VPWR VPWR C_out\[267\] sky130_fd_sc_hd__dfrtp_1
XFILLER_129_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28246_ clknet_leaf_77_clk _02044_ VGND VGND VPWR VPWR systolic_inst.B_shift\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16260_ _03632_ _03640_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__xnor2_1
X_25458_ systolic_inst.cycle_cnt\[9\] systolic_inst.cycle_cnt\[8\] VGND VGND VPWR
+ VPWR _11202_ sky130_fd_sc_hd__and2_1
XFILLER_9_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13472_ deser_A.shift_reg\[36\] deser_A.shift_reg\[37\] deser_A.receiving VGND VGND
+ VPWR VPWR _00309_ sky130_fd_sc_hd__mux2_1
XFILLER_186_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15211_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[14\]\[10\]
+ VGND VGND VPWR VPWR _12315_ sky130_fd_sc_hd__or2_1
X_24409_ C_out\[31\] _11302_ net81 ser_C.shift_reg\[31\] _10674_ VGND VGND VPWR VPWR
+ _02281_ sky130_fd_sc_hd__a221o_1
XFILLER_187_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28177_ clknet_leaf_54_clk _01975_ VGND VGND VPWR VPWR systolic_inst.B_shift\[18\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16191_ _03533_ _03535_ _03573_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__nand3_1
X_25389_ systolic_inst.A_shift\[3\]\[2\] A_in\[18\] net59 VGND VGND VPWR VPWR _11164_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15142_ _12255_ _12256_ VGND VGND VPWR VPWR _12257_ sky130_fd_sc_hd__xnor2_1
X_27128_ clknet_leaf_15_clk _00926_ VGND VGND VPWR VPWR systolic_inst.A_shift\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27059_ clknet_leaf_4_B_in_serial_clk _00857_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_19950_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__inv_2
XFILLER_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15073_ _12177_ _12190_ VGND VGND VPWR VPWR _12191_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_112_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14024_ deser_B.shift_reg\[58\] deser_B.shift_reg\[59\] net125 VGND VGND VPWR VPWR
+ _00850_ sky130_fd_sc_hd__mux2_1
X_18901_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[15\]
+ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__nor2_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19881_ _06822_ _06878_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__or2_1
XFILLER_122_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18832_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[8\]\[5\]
+ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__or2_1
XFILLER_136_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18763_ _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__inv_2
X_15975_ net115 systolic_inst.B_outs\[12\]\[0\] systolic_inst.A_outs\[12\]\[0\] VGND
+ VGND VPWR VPWR _12977_ sky130_fd_sc_hd__and3_1
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _04939_ _04941_ _04942_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__or3_1
X_14926_ _12045_ _12046_ VGND VGND VPWR VPWR _12048_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18694_ _05803_ _05819_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__xor2_1
XFILLER_48_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17645_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[10\]\[11\]
+ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__nor2_1
XFILLER_224_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14857_ _11968_ _11980_ VGND VGND VPWR VPWR _11981_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_82_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13808_ B_in\[115\] deser_B.word_buffer\[115\] net87 VGND VGND VPWR VPWR _00645_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_231_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14788_ systolic_inst.A_outs\[14\]\[0\] systolic_inst.A_outs\[14\]\[1\] systolic_inst.B_outs\[14\]\[3\]
+ systolic_inst.B_outs\[14\]\[4\] VGND VGND VPWR VPWR _11914_ sky130_fd_sc_hd__nand4_1
XFILLER_63_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17576_ net120 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[10\]\[0\]
+ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19315_ _06375_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__inv_2
XFILLER_147_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13739_ B_in\[46\] deser_B.word_buffer\[46\] net84 VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__mux2_1
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16527_ _03880_ _03879_ systolic_inst.acc_wires\[12\]\[23\] net108 VGND VGND VPWR
+ VPWR _01193_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19246_ systolic_inst.B_outs\[7\]\[4\] systolic_inst.A_outs\[7\]\[6\] systolic_inst.A_outs\[7\]\[7\]
+ systolic_inst.B_outs\[7\]\[3\] VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16458_ _03814_ _03817_ _03821_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15409_ _12451_ _12468_ _12470_ VGND VGND VPWR VPWR _12471_ sky130_fd_sc_hd__and3_1
XFILLER_176_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19177_ _06235_ _06241_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16389_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[12\]\[4\]
+ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__nand2_1
XFILLER_185_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_229_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18128_ _05249_ _05252_ _05284_ _05315_ _05282_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__o311a_1
XFILLER_172_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_293_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_293_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_225_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18059_ _05247_ _05248_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_225_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21070_ _07896_ _07897_ _07899_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__o21ba_1
XFILLER_160_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20021_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[6\]\[0\]
+ _07009_ _07010_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__a22o_1
XFILLER_63_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_232_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24760_ net113 ser_C.shift_reg\[208\] VGND VGND VPWR VPWR _10850_ sky130_fd_sc_hd__and2_1
X_21972_ _08749_ _08754_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_176_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_169_Left_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23711_ _10322_ _10323_ _10324_ VGND VGND VPWR VPWR _10325_ sky130_fd_sc_hd__a21o_1
XFILLER_82_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20923_ _07796_ _07797_ _07772_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__and3b_1
X_24691_ C_out\[172\] net104 net76 ser_C.shift_reg\[172\] _10815_ VGND VGND VPWR VPWR
+ _02422_ sky130_fd_sc_hd__a221o_1
XFILLER_148_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26430_ clknet_leaf_2_clk _00237_ net131 VGND VGND VPWR VPWR A_in\[98\] sky130_fd_sc_hd__dfrtp_1
X_23642_ _10260_ _10261_ VGND VGND VPWR VPWR _10262_ sky130_fd_sc_hd__nand2b_1
XFILLER_199_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20854_ _07731_ _07732_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__nor2_1
XFILLER_109_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26361_ clknet_leaf_17_clk _00168_ net134 VGND VGND VPWR VPWR A_in\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23573_ systolic_inst.B_outs\[0\]\[6\] _10193_ VGND VGND VPWR VPWR _10195_ sky130_fd_sc_hd__and2_1
XFILLER_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20785_ _07683_ _07685_ _07688_ net60 VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__a31o_1
X_28100_ clknet_leaf_111_clk _01898_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_165_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25312_ net112 ser_C.shift_reg\[484\] VGND VGND VPWR VPWR _11126_ sky130_fd_sc_hd__and2_1
X_29080_ clknet_leaf_109_clk _02878_ net150 VGND VGND VPWR VPWR C_out\[52\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_214_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22524_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[2\]\[9\]
+ VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__xor2_1
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26292_ clknet_leaf_1_A_in_serial_clk _00100_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28031_ clknet_leaf_160_clk _01829_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_25243_ ser_C.parallel_data\[448\] net102 net74 ser_C.shift_reg\[448\] _11091_ VGND
+ VGND VPWR VPWR _02698_ sky130_fd_sc_hd__a221o_1
X_22455_ _09124_ _09171_ _09170_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__o21ba_1
XFILLER_10_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_178_Left_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21406_ _08247_ _08248_ _08246_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__o21ai_1
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25174_ net110 ser_C.shift_reg\[415\] VGND VGND VPWR VPWR _11057_ sky130_fd_sc_hd__and2_1
XFILLER_198_1170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22386_ systolic_inst.B_outs\[2\]\[6\] systolic_inst.A_outs\[2\]\[6\] _11265_ systolic_inst.A_outs\[2\]\[5\]
+ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_159_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1004 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_284_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_284_clk
+ sky130_fd_sc_hd__clkbuf_8
X_24125_ systolic_inst.A_shift\[30\]\[2\] A_in\[114\] net59 VGND VGND VPWR VPWR _10564_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21337_ _08186_ _08189_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__xor2_1
XFILLER_163_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24056_ _10545_ systolic_inst.B_shift\[0\]\[7\] _11332_ VGND VGND VPWR VPWR _02057_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28933_ clknet_leaf_264_clk _02731_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21268_ net63 _08128_ _08130_ systolic_inst.acc_wires\[4\]\[2\] net108 VGND VGND
+ VPWR VPWR _01684_ sky130_fd_sc_hd__a32o_1
XFILLER_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23007_ _09614_ _09619_ _09648_ _09681_ _09647_ VGND VGND VPWR VPWR _09684_ sky130_fd_sc_hd__a311oi_4
XFILLER_132_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20219_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[31\]
+ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28864_ clknet_leaf_332_clk _02662_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[412\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21199_ _08041_ _08065_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__and2_1
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27815_ clknet_leaf_143_clk _01613_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_187_Left_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28795_ clknet_leaf_233_clk _02593_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[343\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15760_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[13\]\[2\]
+ VGND VGND VPWR VPWR _12808_ sky130_fd_sc_hd__nand2_1
X_27746_ clknet_leaf_211_clk _01544_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24958_ net110 ser_C.shift_reg\[307\] VGND VGND VPWR VPWR _10949_ sky130_fd_sc_hd__and2_1
XFILLER_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14711_ _11855_ _11859_ _11856_ VGND VGND VPWR VPWR _11862_ sky130_fd_sc_hd__a21bo_1
X_23909_ _10487_ systolic_inst.B_shift\[13\]\[6\] net72 VGND VGND VPWR VPWR _01968_
+ sky130_fd_sc_hd__mux2_1
X_15691_ net108 _12744_ VGND VGND VPWR VPWR _12745_ sky130_fd_sc_hd__nor2_1
X_27677_ clknet_leaf_201_clk _01475_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24889_ C_out\[271\] net103 net75 ser_C.shift_reg\[271\] _10914_ VGND VGND VPWR VPWR
+ _02521_ sky130_fd_sc_hd__a221o_1
XFILLER_205_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14642_ _11801_ _11802_ VGND VGND VPWR VPWR _11804_ sky130_fd_sc_hd__nor2_1
X_29416_ clknet_leaf_328_clk _03214_ net136 VGND VGND VPWR VPWR C_out\[388\] sky130_fd_sc_hd__dfrtp_1
XFILLER_61_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17430_ _04684_ _04683_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__nand2b_1
XFILLER_233_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26628_ clknet_leaf_19_B_in_serial_clk _00431_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_159_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14573_ net69 _11742_ _11744_ systolic_inst.acc_wires\[15\]\[6\] net105 VGND VGND
+ VPWR VPWR _00984_ sky130_fd_sc_hd__a32o_1
X_17361_ _04617_ _04616_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__nand2b_1
X_29347_ clknet_leaf_224_clk _03145_ net140 VGND VGND VPWR VPWR C_out\[319\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26559_ clknet_leaf_2_A_in_serial_clk _00362_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19100_ net105 systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[5\] _06166_
+ _06167_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__a22o_1
X_16312_ _03664_ _03691_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__nand2b_1
X_13524_ deser_A.shift_reg\[88\] deser_A.shift_reg\[89\] net129 VGND VGND VPWR VPWR
+ _00361_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17292_ _04548_ _04549_ _04537_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__o21bai_1
XFILLER_198_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29278_ clknet_leaf_188_clk _03076_ net148 VGND VGND VPWR VPWR C_out\[250\] sky130_fd_sc_hd__dfrtp_1
X_19031_ net119 _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__nand2_1
X_16243_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[10\] _03625_
+ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__a21o_1
X_28229_ clknet_leaf_48_clk _02027_ VGND VGND VPWR VPWR systolic_inst.B_shift\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13455_ deser_A.shift_reg\[19\] deser_A.shift_reg\[20\] deser_A.receiving VGND VGND
+ VPWR VPWR _00292_ sky130_fd_sc_hd__mux2_1
XFILLER_16_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16174_ _03517_ _03556_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__and2_1
X_13386_ A_in\[95\] deser_A.word_buffer\[95\] net94 VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_275_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_275_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15125_ _12176_ _12240_ VGND VGND VPWR VPWR _12241_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_110_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19933_ _06896_ _06898_ _06897_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__o21ba_1
XFILLER_138_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15056_ _12030_ _12173_ VGND VGND VPWR VPWR _12174_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_220_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14007_ deser_B.shift_reg\[41\] deser_B.shift_reg\[42\] deser_B.receiving VGND VGND
+ VPWR VPWR _00833_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_220_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19864_ systolic_inst.A_outs\[6\]\[4\] systolic_inst.B_outs\[6\]\[6\] _11278_ systolic_inst.A_outs\[6\]\[3\]
+ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18815_ net63 _05931_ _05933_ systolic_inst.acc_wires\[8\]\[2\] net108 VGND VGND
+ VPWR VPWR _01428_ sky130_fd_sc_hd__a32o_1
X_19795_ _06794_ _06795_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18746_ _05836_ _05839_ _05837_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__o21ba_1
XFILLER_97_1200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15958_ _12976_ _12975_ systolic_inst.acc_wires\[13\]\[31\] net107 VGND VGND VPWR
+ VPWR _01137_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_69_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14909_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[7\]
+ VGND VGND VPWR VPWR _12031_ sky130_fd_sc_hd__o21ai_2
XFILLER_97_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18677_ _05801_ _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__nand2_1
X_15889_ _12916_ _12917_ _12914_ VGND VGND VPWR VPWR _12919_ sky130_fd_sc_hd__o21ai_2
XFILLER_58_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17628_ _04868_ _04867_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__and2b_1
XFILLER_197_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17559_ _04740_ _04809_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20570_ _07435_ _07501_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19229_ _06291_ _06292_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__nand2_1
XFILLER_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_227_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_240_Right_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_227_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22240_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[7\]
+ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__o21ai_2
XFILLER_30_1125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_266_clk clknet_5_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_266_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_200_Left_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22171_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[5\]
+ systolic_inst.A_outs\[2\]\[6\] VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__and4_1
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21122_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\] systolic_inst.A_outs\[4\]\[7\]
+ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21053_ systolic_inst.A_outs\[4\]\[4\] _07884_ _07924_ VGND VGND VPWR VPWR _07925_
+ sky130_fd_sc_hd__a21bo_1
X_25930_ systolic_inst.acc_wires\[12\]\[22\] C_out\[406\] net17 VGND VGND VPWR VPWR
+ _03232_ sky130_fd_sc_hd__mux2_1
XFILLER_113_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20004_ _06995_ _06997_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_54_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25861_ systolic_inst.acc_wires\[10\]\[17\] C_out\[337\] net11 VGND VGND VPWR VPWR
+ _03163_ sky130_fd_sc_hd__mux2_1
XFILLER_101_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24812_ net113 ser_C.shift_reg\[234\] VGND VGND VPWR VPWR _10876_ sky130_fd_sc_hd__and2_1
X_27600_ clknet_leaf_319_clk _01398_ net136 VGND VGND VPWR VPWR systolic_inst.A_outs\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_228_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25792_ systolic_inst.acc_wires\[8\]\[12\] C_out\[268\] net29 VGND VGND VPWR VPWR
+ _03094_ sky130_fd_sc_hd__mux2_1
X_28580_ clknet_leaf_311_clk _02378_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[128\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_234_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24743_ C_out\[198\] net97 net80 ser_C.shift_reg\[198\] _10841_ VGND VGND VPWR VPWR
+ _02448_ sky130_fd_sc_hd__a221o_1
XFILLER_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27531_ clknet_leaf_243_clk _01329_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_21955_ _08742_ VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27462_ clknet_leaf_195_clk _01260_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20906_ _07758_ _07780_ _07781_ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__nand3b_2
XFILLER_203_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24674_ net110 ser_C.shift_reg\[165\] VGND VGND VPWR VPWR _10807_ sky130_fd_sc_hd__and2_1
X_21886_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[3\]\[3\]
+ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__or2_1
XFILLER_128_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29201_ clknet_leaf_142_clk _02999_ net149 VGND VGND VPWR VPWR C_out\[173\] sky130_fd_sc_hd__dfrtp_1
X_23625_ _10220_ _10244_ _10245_ VGND VGND VPWR VPWR _10246_ sky130_fd_sc_hd__nand3_1
X_26413_ clknet_leaf_29_clk _00220_ net133 VGND VGND VPWR VPWR A_in\[81\] sky130_fd_sc_hd__dfrtp_1
X_20837_ systolic_inst.B_outs\[3\]\[2\] systolic_inst.B_shift\[3\]\[2\] net120 VGND
+ VGND VPWR VPWR _01660_ sky130_fd_sc_hd__mux2_1
X_27393_ clknet_leaf_336_clk _01191_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29132_ clknet_leaf_169_clk _02930_ net148 VGND VGND VPWR VPWR C_out\[104\] sky130_fd_sc_hd__dfrtp_1
XFILLER_168_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26344_ clknet_leaf_60_clk _00151_ net135 VGND VGND VPWR VPWR A_in\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_204_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23556_ _10175_ _10177_ _10134_ _10136_ VGND VGND VPWR VPWR _10179_ sky130_fd_sc_hd__o211a_1
X_20768_ _07666_ _07667_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__nor2_1
XFILLER_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29063_ clknet_leaf_114_clk _02861_ net150 VGND VGND VPWR VPWR C_out\[35\] sky130_fd_sc_hd__dfrtp_1
X_22507_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[2\]\[6\]
+ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__or2_1
XFILLER_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26275_ clknet_leaf_17_A_in_serial_clk _00083_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23487_ _10066_ _10110_ VGND VGND VPWR VPWR _10111_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20699_ _07601_ _07607_ _07609_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__o21a_1
XFILLER_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28014_ clknet_leaf_112_clk _01812_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_25226_ net110 ser_C.shift_reg\[441\] VGND VGND VPWR VPWR _11083_ sky130_fd_sc_hd__and2_1
X_13240_ deser_A.word_buffer\[78\] deser_A.serial_word\[78\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__mux2_1
X_22438_ _09176_ _09177_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_257_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_257_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13171_ deser_A.word_buffer\[9\] deser_A.serial_word\[9\] net128 VGND VGND VPWR VPWR
+ _00019_ sky130_fd_sc_hd__mux2_1
X_25157_ C_out\[405\] net101 net73 ser_C.shift_reg\[405\] _11048_ VGND VGND VPWR VPWR
+ _02655_ sky130_fd_sc_hd__a221o_1
X_22369_ _09058_ _09076_ _09075_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__o21a_1
XFILLER_100_1359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24108_ systolic_inst.B_shift\[1\]\[3\] _11332_ net83 systolic_inst.B_shift\[5\]\[3\]
+ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__a22o_1
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25088_ net113 ser_C.shift_reg\[372\] VGND VGND VPWR VPWR _11014_ sky130_fd_sc_hd__and2_1
XFILLER_215_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24039_ systolic_inst.B_shift\[8\]\[7\] B_in\[39\] _00008_ VGND VGND VPWR VPWR _10537_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28916_ clknet_leaf_282_clk _02714_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[464\]
+ sky130_fd_sc_hd__dfrtp_1
X_16930_ _04244_ _04245_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__nor2_1
XFILLER_78_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_A_in_serial_clk clknet_2_0__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_2_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28847_ clknet_leaf_338_clk _02645_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[395\]
+ sky130_fd_sc_hd__dfrtp_1
X_16861_ _04169_ _04177_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18600_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[8\] VGND
+ VGND VPWR VPWR _05729_ sky130_fd_sc_hd__and2_1
X_15812_ _12848_ _12850_ _12852_ systolic_inst.acc_wires\[13\]\[9\] net107 VGND VGND
+ VPWR VPWR _01115_ sky130_fd_sc_hd__a32o_1
X_19580_ _06602_ _06604_ _06610_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__a21o_1
XFILLER_19_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28778_ clknet_leaf_229_clk _02576_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[326\]
+ sky130_fd_sc_hd__dfrtp_1
X_16792_ _04110_ _04111_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__nand2_1
XFILLER_237_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_30_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_219_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18531_ _11259_ _05660_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__xnor2_1
XFILLER_234_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27729_ clknet_leaf_143_clk _01527_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_15743_ _12576_ _12712_ _12785_ _12783_ VGND VGND VPWR VPWR _12794_ sky130_fd_sc_hd__a31oi_1
XFILLER_46_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18462_ _05592_ _05593_ _05585_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__a21oi_1
XFILLER_206_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15674_ _12694_ _12696_ _12726_ VGND VGND VPWR VPWR _12728_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_64_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _04665_ _04666_ _04667_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__and3_1
XFILLER_159_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14625_ _11786_ _11787_ VGND VGND VPWR VPWR _11789_ sky130_fd_sc_hd__nand2_1
XFILLER_57_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18393_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[30\]
+ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__nand2_1
XFILLER_57_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14556_ _11727_ _11728_ _11729_ VGND VGND VPWR VPWR _11730_ sky130_fd_sc_hd__a21o_1
X_17344_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[7\]
+ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__o21a_1
XFILLER_144_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ deser_A.shift_reg\[71\] deser_A.shift_reg\[72\] net129 VGND VGND VPWR VPWR
+ _00344_ sky130_fd_sc_hd__mux2_1
XFILLER_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14487_ _11665_ _11666_ VGND VGND VPWR VPWR _11668_ sky130_fd_sc_hd__and2b_1
X_17275_ _04532_ _04533_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__or2_1
XFILLER_179_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload204 clknet_leaf_76_clk VGND VGND VPWR VPWR clkload204/Y sky130_fd_sc_hd__inv_6
XFILLER_146_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19014_ systolic_inst.A_outs\[7\]\[3\] systolic_inst.A_outs\[6\]\[3\] net119 VGND
+ VGND VPWR VPWR _01461_ sky130_fd_sc_hd__mux2_1
XFILLER_179_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload215 clknet_leaf_58_clk VGND VGND VPWR VPWR clkload215/Y sky130_fd_sc_hd__clkinv_4
X_13438_ deser_A.shift_reg\[2\] deser_A.shift_reg\[3\] deser_A.receiving VGND VGND
+ VPWR VPWR _00275_ sky130_fd_sc_hd__mux2_1
X_16226_ _03607_ _03608_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__nand2b_1
XFILLER_139_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload226 clknet_leaf_136_clk VGND VGND VPWR VPWR clkload226/Y sky130_fd_sc_hd__inv_6
Xclkload237 clknet_leaf_82_clk VGND VGND VPWR VPWR clkload237/X sky130_fd_sc_hd__clkbuf_4
Xclkload248 clknet_leaf_124_clk VGND VGND VPWR VPWR clkload248/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_248_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_248_clk
+ sky130_fd_sc_hd__clkbuf_8
Xclkload259 clknet_leaf_102_clk VGND VGND VPWR VPWR clkload259/Y sky130_fd_sc_hd__clkinvlp_4
X_16157_ _03541_ _03540_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__nand2b_1
X_13369_ A_in\[78\] deser_A.word_buffer\[78\] net96 VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__mux2_1
XFILLER_154_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15108_ _12175_ _12224_ VGND VGND VPWR VPWR _12225_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16088_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[6\] _13081_
+ _13083_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__a22o_1
XFILLER_103_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19916_ _06877_ _06879_ _06913_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__and3_1
X_15039_ _12118_ _12120_ _12156_ VGND VGND VPWR VPWR _12158_ sky130_fd_sc_hd__nand3_1
XFILLER_25_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19847_ _06808_ _06810_ _06846_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19778_ _06714_ _06750_ _06748_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__a21o_1
XFILLER_231_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18729_ _05764_ _05823_ _05822_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__a21oi_1
Xwire12 net13 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_8
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21740_ _08545_ _08546_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__or2_1
XFILLER_3_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21671_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[8\] _08479_ net122
+ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_190_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23410_ systolic_inst.A_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[4\]
+ systolic_inst.B_outs\[0\]\[3\] VGND VGND VPWR VPWR _10036_ sky130_fd_sc_hd__a22oi_1
X_20622_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[5\]\[1\]
+ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__and2_1
X_24390_ net7 ser_C.shift_reg\[23\] VGND VGND VPWR VPWR _10665_ sky130_fd_sc_hd__and2_1
XFILLER_162_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23341_ _09966_ _09967_ _09947_ VGND VGND VPWR VPWR _09969_ sky130_fd_sc_hd__a21bo_1
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20553_ _07394_ _07453_ _07451_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26060_ deser_B.serial_word\[15\] deser_B.shift_reg\[15\] net55 VGND VGND VPWR VPWR
+ _03362_ sky130_fd_sc_hd__mux2_1
X_23272_ net65 _09913_ _09914_ systolic_inst.acc_wires\[1\]\[30\] net109 VGND VGND
+ VPWR VPWR _01904_ sky130_fd_sc_hd__a32o_1
XFILLER_153_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20484_ _07361_ _07418_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__nand2_1
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25011_ C_out\[332\] net97 net80 ser_C.shift_reg\[332\] _10975_ VGND VGND VPWR VPWR
+ _02582_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_239_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_239_clk
+ sky130_fd_sc_hd__clkbuf_8
X_22223_ _08931_ _08967_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__and2_1
XFILLER_192_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22154_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[3\] _08898_ _08899_
+ VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_191_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21105_ _07937_ _07939_ _07975_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_205_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22085_ systolic_inst.A_outs\[2\]\[7\] systolic_inst.A_outs\[1\]\[7\] net122 VGND
+ VGND VPWR VPWR _01785_ sky130_fd_sc_hd__mux2_1
XFILLER_134_1411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26962_ clknet_leaf_25_A_in_serial_clk _00760_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_205_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28701_ clknet_leaf_188_clk _02499_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[249\]
+ sky130_fd_sc_hd__dfrtp_1
X_25913_ systolic_inst.acc_wires\[12\]\[5\] C_out\[389\] net18 VGND VGND VPWR VPWR
+ _03215_ sky130_fd_sc_hd__mux2_1
X_21036_ _07907_ _07908_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__nor2_1
X_29681_ clknet_leaf_106_clk _03476_ net151 VGND VGND VPWR VPWR ser_C.bit_idx\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_26893_ clknet_leaf_7_A_in_serial_clk _00691_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28632_ clknet_leaf_181_clk _02430_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[180\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_143_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25844_ systolic_inst.acc_wires\[10\]\[0\] C_out\[320\] net14 VGND VGND VPWR VPWR
+ _03146_ sky130_fd_sc_hd__mux2_1
XFILLER_86_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28563_ clknet_leaf_167_clk _02361_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_234_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22987_ _09663_ _09662_ VGND VGND VPWR VPWR _09664_ sky130_fd_sc_hd__nand2b_1
X_25775_ systolic_inst.acc_wires\[7\]\[27\] C_out\[251\] net44 VGND VGND VPWR VPWR
+ _03077_ sky130_fd_sc_hd__mux2_1
XFILLER_43_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27514_ clknet_leaf_225_clk _01312_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_21938_ _08725_ _08726_ VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__nand2_1
X_24726_ net113 ser_C.shift_reg\[191\] VGND VGND VPWR VPWR _10833_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_156_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28494_ clknet_leaf_117_clk _02292_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24657_ C_out\[155\] net104 _10643_ ser_C.shift_reg\[155\] _10798_ VGND VGND VPWR
+ VPWR _02405_ sky130_fd_sc_hd__a221o_1
XFILLER_128_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27445_ clknet_leaf_242_clk _01243_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_21869_ net122 _08668_ _08669_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_106_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14410_ _11447_ _11592_ VGND VGND VPWR VPWR _11593_ sky130_fd_sc_hd__xnor2_4
XFILLER_208_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23608_ _11268_ systolic_inst.B_outs\[0\]\[7\] _10120_ VGND VGND VPWR VPWR _10229_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15390_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[2\]
+ systolic_inst.A_outs\[13\]\[3\] VGND VGND VPWR VPWR _12453_ sky130_fd_sc_hd__nand4_2
X_24588_ net114 ser_C.shift_reg\[122\] VGND VGND VPWR VPWR _10764_ sky130_fd_sc_hd__and2_1
X_27376_ clknet_leaf_328_clk _01174_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_230_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29115_ clknet_leaf_158_clk _02913_ net151 VGND VGND VPWR VPWR C_out\[87\] sky130_fd_sc_hd__dfrtp_1
X_14341_ _11524_ _11525_ VGND VGND VPWR VPWR _11526_ sky130_fd_sc_hd__nor2_1
X_23539_ _10080_ _10122_ _10160_ VGND VGND VPWR VPWR _10162_ sky130_fd_sc_hd__nor3_1
X_26327_ clknet_leaf_0_A_in_serial_clk _00135_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_211_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17060_ net60 _04359_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__nor2_1
X_29046_ clknet_leaf_101_clk _02844_ net151 VGND VGND VPWR VPWR C_out\[18\] sky130_fd_sc_hd__dfrtp_1
X_14272_ _11417_ _11456_ VGND VGND VPWR VPWR _11459_ sky130_fd_sc_hd__xor2_1
X_26258_ clknet_leaf_4_A_in_serial_clk _00066_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_184_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16011_ _13008_ VGND VGND VPWR VPWR _13009_ sky130_fd_sc_hd__inv_2
XFILLER_183_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25209_ C_out\[431\] net101 net73 ser_C.shift_reg\[431\] _11074_ VGND VGND VPWR VPWR
+ _02681_ sky130_fd_sc_hd__a221o_1
X_13223_ deser_A.word_buffer\[61\] deser_A.serial_word\[61\] net128 VGND VGND VPWR
+ VPWR _00071_ sky130_fd_sc_hd__mux2_1
X_26189_ _11302_ _11254_ VGND VGND VPWR VPWR _11255_ sky130_fd_sc_hd__nor2_1
XFILLER_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13154_ net58 _11304_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__nor2_1
XFILLER_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17962_ systolic_inst.B_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[4\]
+ systolic_inst.A_outs\[9\]\[5\] VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_109_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19701_ _06675_ _06703_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__or2_1
X_16913_ _04227_ _04228_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__and2_1
X_17893_ systolic_inst.A_outs\[9\]\[2\] systolic_inst.B_outs\[9\]\[3\] systolic_inst.A_outs\[9\]\[3\]
+ systolic_inst.B_outs\[9\]\[4\] VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__and4_1
XFILLER_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19632_ net119 _06639_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__nand2_1
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16844_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[10\] _04162_
+ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__a21bo_1
XFILLER_238_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19563_ _06552_ _06553_ _06575_ _06595_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__a211o_1
XFILLER_150_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16775_ _04057_ _04093_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__and2_1
X_13987_ deser_B.shift_reg\[21\] deser_B.shift_reg\[22\] net125 VGND VGND VPWR VPWR
+ _00813_ sky130_fd_sc_hd__mux2_1
XFILLER_234_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18514_ _05643_ _05644_ _05632_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__or3b_1
XFILLER_234_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15726_ _12751_ _12754_ _12777_ VGND VGND VPWR VPWR _12778_ sky130_fd_sc_hd__a21oi_1
XFILLER_46_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19494_ _06532_ _06534_ _06537_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_124_Left_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18445_ _05564_ _05566_ _05577_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__a21oi_1
X_15657_ net108 _12710_ _12711_ _12680_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_17_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14608_ _11750_ _11773_ _11763_ _11772_ VGND VGND VPWR VPWR _11774_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_222_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18376_ net105 systolic_inst.acc_wires\[9\]\[27\] net66 _05533_ VGND VGND VPWR VPWR
+ _01389_ sky130_fd_sc_hd__a22o_1
X_15588_ _12577_ _12643_ VGND VGND VPWR VPWR _12644_ sky130_fd_sc_hd__nor2_1
XFILLER_30_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17327_ _04546_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__or2_1
XFILLER_30_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14539_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[15\]\[2\]
+ VGND VGND VPWR VPWR _11715_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_135_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17258_ _04516_ _04517_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_96_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16209_ _03590_ _03591_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_133_Left_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17189_ systolic_inst.B_outs\[9\]\[3\] systolic_inst.B_outs\[5\]\[3\] net116 VGND
+ VGND VPWR VPWR _01277_ sky130_fd_sc_hd__mux2_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_241_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_241_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_200_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22910_ systolic_inst.B_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[6\] systolic_inst.A_outs\[1\]\[7\]
+ systolic_inst.B_outs\[1\]\[3\] VGND VGND VPWR VPWR _09589_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23890_ _10472_ _10475_ VGND VGND VPWR VPWR _10477_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_200_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22841_ systolic_inst.B_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[5\]
+ systolic_inst.B_outs\[1\]\[3\] VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__a22oi_1
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_142_Left_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_192_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25560_ systolic_inst.acc_wires\[1\]\[4\] C_out\[36\] net36 VGND VGND VPWR VPWR _02862_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22772_ _09424_ _09454_ VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__nand2_1
XFILLER_140_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24511_ C_out\[82\] _11302_ net81 ser_C.shift_reg\[82\] _10725_ VGND VGND VPWR VPWR
+ _02332_ sky130_fd_sc_hd__a221o_1
XFILLER_25_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21723_ _08521_ _08529_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__nand2_1
XFILLER_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25491_ _11223_ _11224_ systolic_inst.cycle_cnt\[19\] VGND VGND VPWR VPWR _02813_
+ sky130_fd_sc_hd__mux2_1
XFILLER_213_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24442_ net114 ser_C.shift_reg\[49\] VGND VGND VPWR VPWR _10691_ sky130_fd_sc_hd__and2_1
XFILLER_197_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27230_ clknet_leaf_276_clk _01028_ net138 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_185_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21654_ _08388_ _08422_ _08424_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__a21oi_1
X_20605_ _07463_ _07535_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27161_ clknet_leaf_297_clk _00959_ net138 VGND VGND VPWR VPWR systolic_inst.B_outs\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_24373_ C_out\[13\] net104 _10643_ ser_C.shift_reg\[13\] _10656_ VGND VGND VPWR VPWR
+ _02263_ sky130_fd_sc_hd__a221o_1
XFILLER_36_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21585_ _08350_ _08352_ _08394_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__and3_1
XFILLER_138_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26112_ deser_B.serial_word\[67\] deser_B.shift_reg\[67\] _00001_ VGND VGND VPWR
+ VPWR _03414_ sky130_fd_sc_hd__mux2_1
XFILLER_21_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23324_ _09945_ _09947_ _09950_ _09951_ VGND VGND VPWR VPWR _09953_ sky130_fd_sc_hd__a22o_1
XFILLER_138_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27092_ clknet_leaf_5_B_in_serial_clk _00890_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_20536_ systolic_inst.B_outs\[5\]\[5\] systolic_inst.A_outs\[5\]\[7\] VGND VGND VPWR
+ VPWR _07469_ sky130_fd_sc_hd__nand2_1
XFILLER_126_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_186_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26043_ systolic_inst.B_outs\[15\]\[7\] systolic_inst.B_outs\[11\]\[7\] net118 VGND
+ VGND VPWR VPWR _03345_ sky130_fd_sc_hd__mux2_1
X_23255_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[28\]
+ VGND VGND VPWR VPWR _09900_ sky130_fd_sc_hd__or2_1
X_20467_ systolic_inst.A_outs\[5\]\[3\] systolic_inst.A_outs\[5\]\[4\] systolic_inst.B_outs\[5\]\[6\]
+ systolic_inst.B_outs\[5\]\[7\] VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__and4b_1
XFILLER_181_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22206_ _08951_ _08947_ VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__nand2b_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23186_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[16\]
+ _09838_ VGND VGND VPWR VPWR _09842_ sky130_fd_sc_hd__a21oi_1
X_20398_ systolic_inst.A_outs\[5\]\[2\] systolic_inst.B_outs\[5\]\[6\] _07333_ VGND
+ VGND VPWR VPWR _07335_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_145_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22137_ _08864_ _08867_ _08884_ _08885_ VGND VGND VPWR VPWR _08886_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_145_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27994_ clknet_leaf_127_clk _01792_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_22068_ _08832_ _08836_ VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_141_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26945_ clknet_leaf_25_A_in_serial_clk _00743_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21019_ _07888_ _07891_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13910_ deser_A.serial_word\[71\] deser_A.shift_reg\[71\] net57 VGND VGND VPWR VPWR
+ _00736_ sky130_fd_sc_hd__mux2_1
X_29664_ clknet_leaf_10_B_in_serial_clk _03459_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_181_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26876_ clknet_leaf_13_A_in_serial_clk _00674_ net144 VGND VGND VPWR VPWR deser_A.serial_word\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14890_ _12005_ _12011_ VGND VGND VPWR VPWR _12013_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28615_ clknet_leaf_218_clk _02413_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[163\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_807 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13841_ deser_A.serial_word\[2\] deser_A.shift_reg\[2\] net58 VGND VGND VPWR VPWR
+ _00667_ sky130_fd_sc_hd__mux2_1
X_25827_ systolic_inst.acc_wires\[9\]\[15\] C_out\[303\] net15 VGND VGND VPWR VPWR
+ _03129_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29595_ clknet_leaf_14_B_in_serial_clk _03390_ net152 VGND VGND VPWR VPWR deser_B.serial_word\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28546_ clknet_leaf_164_clk _02344_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_204_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13772_ B_in\[79\] deser_B.word_buffer\[79\] net86 VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__mux2_1
X_16560_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[29\]
+ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__xor2_1
XFILLER_222_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25758_ systolic_inst.acc_wires\[7\]\[10\] C_out\[234\] net42 VGND VGND VPWR VPWR
+ _03060_ sky130_fd_sc_hd__mux2_1
XFILLER_204_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15511_ _12537_ _12568_ VGND VGND VPWR VPWR _12570_ sky130_fd_sc_hd__xnor2_1
X_24709_ C_out\[181\] net99 net79 ser_C.shift_reg\[181\] _10824_ VGND VGND VPWR VPWR
+ _02431_ sky130_fd_sc_hd__a221o_1
XFILLER_128_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28477_ clknet_leaf_106_clk _02275_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_16491_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[18\]
+ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__or2_1
XFILLER_215_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25689_ systolic_inst.acc_wires\[5\]\[5\] C_out\[165\] net16 VGND VGND VPWR VPWR
+ _02991_ sky130_fd_sc_hd__mux2_1
XFILLER_203_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18230_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[9\]\[6\]
+ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__nand2_1
XFILLER_31_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15442_ _12461_ _12478_ _12477_ VGND VGND VPWR VPWR _12503_ sky130_fd_sc_hd__a21bo_1
X_27428_ clknet_leaf_249_clk _01226_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_230_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18161_ systolic_inst.B_outs\[9\]\[5\] systolic_inst.B_outs\[9\]\[6\] systolic_inst.A_outs\[9\]\[7\]
+ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__nand3_1
XFILLER_230_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27359_ clknet_leaf_327_clk _01157_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15373_ net107 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[0\] _12438_
+ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__a21o_1
XFILLER_106_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17112_ _04395_ _04401_ _04402_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14324_ _11470_ _11472_ _11509_ VGND VGND VPWR VPWR _11510_ sky130_fd_sc_hd__o21ai_1
XFILLER_102_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18092_ _05243_ _05245_ _05281_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__nand3_1
XFILLER_144_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29029_ clknet_leaf_128_clk _02827_ net144 VGND VGND VPWR VPWR C_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_14255_ _11438_ _11440_ systolic_inst.B_outs\[15\]\[7\] VGND VGND VPWR VPWR _11442_
+ sky130_fd_sc_hd__a21oi_1
X_17043_ _04337_ _04339_ _04335_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_130_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap129 net130 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_12
X_13206_ deser_A.word_buffer\[44\] deser_A.serial_word\[44\] net127 VGND VGND VPWR
+ VPWR _00054_ sky130_fd_sc_hd__mux2_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14186_ _11354_ _11356_ _11374_ net107 VGND VGND VPWR VPWR _11376_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_91_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13137_ _11286_ _11287_ _11289_ VGND VGND VPWR VPWR _11290_ sky130_fd_sc_hd__or3_1
XFILLER_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18994_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[29\]
+ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__xor2_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17945_ _05109_ _05138_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__nand2b_1
XFILLER_152_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17876_ _05041_ _05070_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__or2_1
XFILLER_241_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19615_ systolic_inst.A_outs\[6\]\[3\] systolic_inst.A_outs\[5\]\[3\] net120 VGND
+ VGND VPWR VPWR _01525_ sky130_fd_sc_hd__mux2_1
XFILLER_4_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16827_ _04108_ _04110_ _04144_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__nand3_1
XFILLER_26_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19546_ _06573_ _06579_ _06580_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__a21oi_1
X_16758_ _04061_ _04078_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15709_ _12761_ _12760_ VGND VGND VPWR VPWR _12762_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_234_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_4_B_in_serial_clk clknet_2_2__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_4_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_19477_ _06515_ _06517_ _06513_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__a21bo_1
X_16689_ _04009_ _04010_ _03987_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_234_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18428_ _05561_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__or2_1
XFILLER_22_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18359_ _05514_ _05516_ _05519_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__a21oi_2
XFILLER_187_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21370_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[17\]
+ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__xor2_1
XFILLER_30_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20321_ _07255_ _07258_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23040_ systolic_inst.A_outs\[1\]\[6\] _11277_ _09686_ _09689_ _09714_ VGND VGND
+ VPWR VPWR _09715_ sky130_fd_sc_hd__o311a_1
X_20252_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[2\] _07193_ VGND
+ VGND VPWR VPWR _07195_ sky130_fd_sc_hd__a21o_1
XFILLER_200_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_181_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20183_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[25\]
+ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__xor2_2
XFILLER_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24991_ C_out\[322\] net102 net80 ser_C.shift_reg\[322\] _10965_ VGND VGND VPWR VPWR
+ _02572_ sky130_fd_sc_hd__a221o_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26730_ clknet_leaf_78_clk _00532_ net143 VGND VGND VPWR VPWR B_in\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23942_ systolic_inst.B_shift\[14\]\[3\] B_in\[19\] net59 VGND VGND VPWR VPWR _10500_
+ sky130_fd_sc_hd__mux2_1
X_23873_ _10446_ _10448_ _10460_ _10461_ _10454_ VGND VGND VPWR VPWR _10462_ sky130_fd_sc_hd__a311oi_4
X_26661_ clknet_leaf_2_B_in_serial_clk _00464_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_179_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28400_ clknet_leaf_319_clk _02198_ VGND VGND VPWR VPWR systolic_inst.A_shift\[16\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25612_ systolic_inst.acc_wires\[2\]\[24\] C_out\[88\] net51 VGND VGND VPWR VPWR
+ _02914_ sky130_fd_sc_hd__mux2_1
X_22824_ _09503_ _09504_ _09453_ _09455_ VGND VGND VPWR VPWR _09506_ sky130_fd_sc_hd__o211a_1
XFILLER_44_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29380_ clknet_leaf_247_clk _03178_ net145 VGND VGND VPWR VPWR C_out\[352\] sky130_fd_sc_hd__dfrtp_1
X_26592_ clknet_leaf_30_A_in_serial_clk _00395_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28331_ clknet_leaf_2_clk _02129_ VGND VGND VPWR VPWR systolic_inst.A_shift\[27\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25543_ systolic_inst.acc_wires\[0\]\[19\] C_out\[19\] net54 VGND VGND VPWR VPWR
+ _02845_ sky130_fd_sc_hd__mux2_1
X_22755_ _09427_ _09437_ VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__xor2_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21706_ net122 _08511_ _08512_ _08513_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__a31o_1
XFILLER_38_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25474_ _11212_ _11213_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__and2_1
X_28262_ clknet_leaf_48_clk _02060_ VGND VGND VPWR VPWR systolic_inst.B_shift\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_22686_ systolic_inst.B_outs\[0\]\[5\] systolic_inst.B_shift\[0\]\[5\] net121 VGND
+ VGND VPWR VPWR _01855_ sky130_fd_sc_hd__mux2_1
XFILLER_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24425_ C_out\[39\] _11302_ net81 ser_C.shift_reg\[39\] _10682_ VGND VGND VPWR VPWR
+ _02289_ sky130_fd_sc_hd__a221o_1
X_27213_ clknet_leaf_294_clk _01011_ net138 VGND VGND VPWR VPWR systolic_inst.A_outs\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_212_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21637_ _08441_ _08444_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28193_ clknet_leaf_129_clk _01991_ VGND VGND VPWR VPWR systolic_inst.B_shift\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_170_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24356_ net7 ser_C.shift_reg\[6\] VGND VGND VPWR VPWR _10648_ sky130_fd_sc_hd__and2_1
X_27144_ clknet_leaf_5_clk _00942_ VGND VGND VPWR VPWR systolic_inst.A_shift\[21\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_21568_ _08348_ _08377_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__nor2_1
XFILLER_166_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_185_Right_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23307_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[3\] _09935_ VGND
+ VGND VPWR VPWR _09937_ sky130_fd_sc_hd__and3_1
Xclkbuf_5_16__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_16__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_126_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27075_ clknet_leaf_26_B_in_serial_clk _00873_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20519_ _07451_ _07452_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__nor2_1
XFILLER_197_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24287_ systolic_inst.B_shift\[27\]\[7\] B_in\[95\] _00008_ VGND VGND VPWR VPWR _10617_
+ sky130_fd_sc_hd__mux2_1
X_21499_ systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[3\] VGND VGND VPWR
+ VPWR _08313_ sky130_fd_sc_hd__nand2_1
XFILLER_154_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14040_ deser_B.shift_reg\[74\] deser_B.shift_reg\[75\] deser_B.receiving VGND VGND
+ VPWR VPWR _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23238_ _09881_ _09883_ _09885_ VGND VGND VPWR VPWR _09886_ sky130_fd_sc_hd__or3_1
XFILLER_158_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26026_ systolic_inst.acc_wires\[15\]\[22\] ser_C.parallel_data\[502\] net37 VGND
+ VGND VPWR VPWR _03328_ sky130_fd_sc_hd__mux2_1
XFILLER_106_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23169_ net65 _09826_ _09827_ systolic_inst.acc_wires\[1\]\[14\] net109 VGND VGND
+ VPWR VPWR _01888_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_8_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27977_ clknet_leaf_169_clk _01775_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_164_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15991_ systolic_inst.A_outs\[12\]\[1\] systolic_inst.B_outs\[12\]\[2\] systolic_inst.B_outs\[12\]\[3\]
+ systolic_inst.A_outs\[12\]\[0\] VGND VGND VPWR VPWR _12990_ sky130_fd_sc_hd__a22oi_1
XFILLER_216_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17730_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[23\]
+ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__xor2_1
X_14942_ _12061_ _12063_ VGND VGND VPWR VPWR _12064_ sky130_fd_sc_hd__and2_1
X_26928_ clknet_leaf_5_A_in_serial_clk _00726_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29647_ clknet_leaf_1_B_in_serial_clk _03442_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_17661_ net105 systolic_inst.acc_wires\[10\]\[12\] _11712_ _04897_ VGND VGND VPWR
+ VPWR _01310_ sky130_fd_sc_hd__a22o_1
X_26859_ clknet_leaf_0_B_in_serial_clk _00661_ net134 VGND VGND VPWR VPWR deser_B.bit_idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14873_ _11264_ _11995_ VGND VGND VPWR VPWR _11996_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19400_ net119 _06447_ _06457_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16612_ _03935_ _03936_ _03926_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__a21o_1
X_13824_ net126 net3 VGND VGND VPWR VPWR _11321_ sky130_fd_sc_hd__nand2b_1
X_29578_ clknet_leaf_23_B_in_serial_clk _03373_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_17592_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[10\]\[3\]
+ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__nand2_1
Xclkbuf_2_0__f_A_in_serial_clk clknet_0_A_in_serial_clk VGND VGND VPWR VPWR clknet_2_0__leaf_A_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19331_ _06389_ _06390_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__xnor2_1
X_28529_ clknet_leaf_166_clk _02327_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_188_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16543_ _03893_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__inv_2
XFILLER_56_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13755_ B_in\[62\] deser_B.word_buffer\[62\] net87 VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__mux2_1
XFILLER_44_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19262_ _06323_ _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__nand2b_1
XFILLER_189_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16474_ _03834_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13686_ deser_B.word_buffer\[122\] deser_B.serial_word\[122\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18213_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__inv_2
XFILLER_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15425_ _12484_ _12485_ VGND VGND VPWR VPWR _12486_ sky130_fd_sc_hd__nor2_1
XFILLER_176_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19193_ _06182_ _06217_ _06219_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18144_ _05262_ _05300_ _05299_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__a21bo_1
X_15356_ systolic_inst.A_outs\[13\]\[0\] systolic_inst.A_outs\[12\]\[0\] net115 VGND
+ VGND VPWR VPWR _01074_ sky130_fd_sc_hd__mux2_1
XFILLER_141_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14307_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[5\] _11455_ _11454_
+ VGND VGND VPWR VPWR _11493_ sky130_fd_sc_hd__a31o_1
XFILLER_176_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18075_ systolic_inst.A_outs\[9\]\[5\] systolic_inst.B_outs\[9\]\[6\] _11263_ systolic_inst.A_outs\[9\]\[4\]
+ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__o2bb2a_1
X_15287_ _11712_ _12379_ _12380_ systolic_inst.acc_wires\[14\]\[20\] net107 VGND VGND
+ VPWR VPWR _01062_ sky130_fd_sc_hd__a32o_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_242_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17026_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[11\]\[8\]
+ _04327_ _04329_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_242_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14238_ _11425_ VGND VGND VPWR VPWR _11426_ sky130_fd_sc_hd__inv_2
XFILLER_171_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14169_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[3\]
+ systolic_inst.B_outs\[15\]\[1\] VGND VGND VPWR VPWR _11359_ sky130_fd_sc_hd__a22oi_1
XFILLER_98_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xload_slew132 net134 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_16
Xload_slew143 net144 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_16
X_18977_ _06070_ _06071_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__nand2_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17928_ _05120_ _05121_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17859_ _05054_ _05051_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_236_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_236_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20870_ _07735_ _07747_ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__and2_1
XFILLER_226_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19529_ _06565_ _06567_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__xor2_1
XFILLER_241_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22540_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[2\]\[11\]
+ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__nand2_1
XFILLER_179_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22471_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[2\]\[1\]
+ VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__and2_1
XFILLER_210_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24210_ _10590_ systolic_inst.A_shift\[20\]\[4\] net71 VGND VGND VPWR VPWR _02166_
+ sky130_fd_sc_hd__mux2_1
X_21422_ _08256_ _08258_ _08261_ _11713_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__a31o_1
X_25190_ net111 ser_C.shift_reg\[423\] VGND VGND VPWR VPWR _11065_ sky130_fd_sc_hd__and2_1
XFILLER_198_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24141_ systolic_inst.A_shift\[29\]\[2\] A_in\[106\] net59 VGND VGND VPWR VPWR _10572_
+ sky130_fd_sc_hd__mux2_1
XFILLER_175_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21353_ net63 _08202_ _08203_ systolic_inst.acc_wires\[4\]\[14\] _11258_ VGND VGND
+ VPWR VPWR _01696_ sky130_fd_sc_hd__a32o_1
XFILLER_175_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20304_ _07233_ _07243_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__nor2_1
X_24072_ _10553_ systolic_inst.B_shift\[15\]\[7\] net71 VGND VGND VPWR VPWR _02065_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21284_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[4\]\[5\]
+ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__nand2_1
XFILLER_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23023_ _09696_ _09697_ VGND VGND VPWR VPWR _09699_ sky130_fd_sc_hd__xor2_1
X_27900_ clknet_leaf_42_clk _01698_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20235_ systolic_inst.B_outs\[4\]\[4\] systolic_inst.B_outs\[0\]\[4\] net117 VGND
+ VGND VPWR VPWR _01598_ sky130_fd_sc_hd__mux2_1
XFILLER_116_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28880_ clknet_leaf_288_clk _02678_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[428\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_157_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27831_ clknet_leaf_142_clk _01629_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_20166_ net62 _07135_ _07136_ systolic_inst.acc_wires\[6\]\[22\] net106 VGND VGND
+ VPWR VPWR _01576_ sky130_fd_sc_hd__a32o_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27762_ clknet_leaf_211_clk _01560_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_20097_ _07076_ _07077_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__nor2_1
X_24974_ net111 ser_C.shift_reg\[315\] VGND VGND VPWR VPWR _10957_ sky130_fd_sc_hd__and2_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29501_ clknet_leaf_268_clk _03299_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[473\]
+ sky130_fd_sc_hd__dfrtp_1
X_26713_ clknet_leaf_26_B_in_serial_clk _00516_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_217_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23925_ _10495_ systolic_inst.B_shift\[18\]\[6\] net71 VGND VGND VPWR VPWR _01976_
+ sky130_fd_sc_hd__mux2_1
X_27693_ clknet_leaf_200_clk _01491_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29432_ clknet_leaf_336_clk _03230_ net131 VGND VGND VPWR VPWR C_out\[404\] sky130_fd_sc_hd__dfrtp_1
XFILLER_229_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26644_ clknet_leaf_14_B_in_serial_clk _00447_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_229_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23856_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[25\]
+ VGND VGND VPWR VPWR _10448_ sky130_fd_sc_hd__xor2_2
XFILLER_44_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22807_ systolic_inst.A_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[5\] VGND VGND VPWR
+ VPWR _09489_ sky130_fd_sc_hd__nand2_1
X_29363_ clknet_leaf_225_clk _03161_ net140 VGND VGND VPWR VPWR C_out\[335\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26575_ clknet_leaf_24_A_in_serial_clk _00378_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_23787_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[0\]\[13\]
+ _10385_ VGND VGND VPWR VPWR _10390_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20999_ _07805_ _07842_ _07841_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__a21bo_1
XFILLER_213_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28314_ clknet_leaf_9_clk _02112_ VGND VGND VPWR VPWR systolic_inst.A_shift\[29\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25526_ systolic_inst.acc_wires\[0\]\[2\] C_out\[2\] net33 VGND VGND VPWR VPWR _02828_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13540_ deser_A.shift_reg\[104\] deser_A.shift_reg\[105\] net129 VGND VGND VPWR VPWR
+ _00377_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22738_ _09403_ _09405_ _09404_ VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__a21bo_1
X_29294_ clknet_leaf_315_clk _03092_ net142 VGND VGND VPWR VPWR C_out\[266\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28245_ clknet_leaf_73_clk _02043_ VGND VGND VPWR VPWR systolic_inst.B_shift\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13471_ deser_A.shift_reg\[35\] deser_A.shift_reg\[36\] deser_A.receiving VGND VGND
+ VPWR VPWR _00308_ sky130_fd_sc_hd__mux2_1
X_25457_ _11200_ _11201_ systolic_inst.cycle_cnt\[8\] VGND VGND VPWR VPWR _02802_
+ sky130_fd_sc_hd__mux2_1
X_22669_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[31\]
+ VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15210_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[14\]\[10\]
+ VGND VGND VPWR VPWR _12314_ sky130_fd_sc_hd__nand2_1
X_24408_ net114 ser_C.shift_reg\[32\] VGND VGND VPWR VPWR _10674_ sky130_fd_sc_hd__and2_1
XFILLER_16_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28176_ clknet_leaf_75_clk _01974_ VGND VGND VPWR VPWR systolic_inst.B_shift\[18\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16190_ _03533_ _03535_ _03573_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__a21o_1
XFILLER_142_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25388_ _11163_ systolic_inst.A_shift\[2\]\[1\] net71 VGND VGND VPWR VPWR _02771_
+ sky130_fd_sc_hd__mux2_1
XFILLER_187_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15141_ _12174_ _12235_ VGND VGND VPWR VPWR _12256_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27127_ clknet_leaf_16_clk _00925_ VGND VGND VPWR VPWR systolic_inst.A_shift\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24339_ systolic_inst.A_shift\[8\]\[2\] net70 net83 systolic_inst.A_shift\[9\]\[2\]
+ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__a22o_1
XFILLER_177_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15072_ _12188_ _12189_ VGND VGND VPWR VPWR _12190_ sky130_fd_sc_hd__nand2_1
X_27058_ clknet_leaf_4_B_in_serial_clk _00856_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_141_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14023_ deser_B.shift_reg\[57\] deser_B.shift_reg\[58\] net125 VGND VGND VPWR VPWR
+ _00849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18900_ net63 _06005_ _06006_ systolic_inst.acc_wires\[8\]\[14\] net108 VGND VGND
+ VPWR VPWR _01440_ sky130_fd_sc_hd__a32o_1
XFILLER_84_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26009_ systolic_inst.acc_wires\[15\]\[5\] ser_C.parallel_data\[485\] net23 VGND
+ VGND VPWR VPWR _03311_ sky130_fd_sc_hd__mux2_1
X_19880_ _06822_ _06878_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__nand2_1
XFILLER_175_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18831_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[8\]\[5\]
+ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18762_ _05850_ _05852_ _05884_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__nor3_1
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15974_ systolic_inst.B_outs\[11\]\[7\] systolic_inst.B_outs\[7\]\[7\] net118 VGND
+ VGND VPWR VPWR _01153_ sky130_fd_sc_hd__mux2_1
XFILLER_212_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17713_ systolic_inst.acc_wires\[10\]\[16\] systolic_inst.acc_wires\[10\]\[17\] systolic_inst.acc_wires\[10\]\[18\]
+ systolic_inst.acc_wires\[10\]\[19\] systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__o41a_1
X_14925_ _12046_ _12045_ VGND VGND VPWR VPWR _12047_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_121_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18693_ _05817_ _05818_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_121_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _11712_ _04881_ _04882_ systolic_inst.acc_wires\[10\]\[10\] net105 VGND VGND
+ VPWR VPWR _01308_ sky130_fd_sc_hd__a32o_1
XFILLER_236_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14856_ _11948_ _11979_ VGND VGND VPWR VPWR _11980_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_82_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13807_ B_in\[114\] deser_B.word_buffer\[114\] net85 VGND VGND VPWR VPWR _00644_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_231_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17575_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[10\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_231_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_221_Right_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14787_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[2\] VGND VGND
+ VPWR VPWR _11913_ sky130_fd_sc_hd__and2_1
X_19314_ _06373_ _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__nand2_1
XFILLER_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16526_ _03871_ _03875_ _03877_ net61 VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__a31o_1
XFILLER_220_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13738_ B_in\[45\] deser_B.word_buffer\[45\] net84 VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__mux2_1
XFILLER_188_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19245_ _06306_ _06307_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_119_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16457_ _03819_ _03820_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__and2_1
X_13669_ deser_B.word_buffer\[105\] deser_B.serial_word\[105\] net123 VGND VGND VPWR
+ VPWR _00506_ sky130_fd_sc_hd__mux2_1
XFILLER_176_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15408_ systolic_inst.A_outs\[13\]\[4\] _12469_ VGND VGND VPWR VPWR _12470_ sky130_fd_sc_hd__nand2_1
X_19176_ _06236_ _06239_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16388_ net67 _03759_ _03761_ systolic_inst.acc_wires\[12\]\[3\] net108 VGND VGND
+ VPWR VPWR _01173_ sky130_fd_sc_hd__a32o_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18127_ _05249_ _05252_ _05284_ _05282_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_229_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15339_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[29\]
+ VGND VGND VPWR VPWR _12424_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_229_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18058_ _05247_ _05248_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_225_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17009_ _04309_ _04310_ _04308_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__a21bo_1
XFILLER_104_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20020_ _07011_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_176_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21971_ _08756_ _08755_ systolic_inst.acc_wires\[3\]\[15\] net106 VGND VGND VPWR
+ VPWR _01761_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_176_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23710_ _10317_ _10318_ _10316_ VGND VGND VPWR VPWR _10324_ sky130_fd_sc_hd__a21bo_1
XFILLER_55_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20922_ _07796_ _07797_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__nand2b_1
X_24690_ net112 ser_C.shift_reg\[173\] VGND VGND VPWR VPWR _10815_ sky130_fd_sc_hd__and2_1
XFILLER_187_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23641_ _10080_ _10230_ _10259_ VGND VGND VPWR VPWR _10261_ sky130_fd_sc_hd__or3_1
XFILLER_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20853_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[2\] _07728_ _07730_
+ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__a22oi_1
XFILLER_242_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23572_ systolic_inst.A_outs\[0\]\[5\] systolic_inst.B_outs\[0\]\[6\] _10193_ VGND
+ VGND VPWR VPWR _10194_ sky130_fd_sc_hd__a21oi_1
X_26360_ clknet_leaf_18_clk _00167_ net134 VGND VGND VPWR VPWR A_in\[28\] sky130_fd_sc_hd__dfrtp_1
X_20784_ _07683_ _07685_ _07688_ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__a21oi_2
XFILLER_167_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22523_ _09251_ _09250_ systolic_inst.acc_wires\[2\]\[8\] net109 VGND VGND VPWR VPWR
+ _01818_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_168_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25311_ ser_C.parallel_data\[482\] net102 net74 ser_C.shift_reg\[482\] _11125_ VGND
+ VGND VPWR VPWR _02732_ sky130_fd_sc_hd__a221o_1
XFILLER_210_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26291_ clknet_leaf_2_A_in_serial_clk _00099_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_214_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28030_ clknet_leaf_160_clk _01828_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22454_ _09124_ _09192_ VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__xnor2_1
X_25242_ net111 ser_C.shift_reg\[449\] VGND VGND VPWR VPWR _11091_ sky130_fd_sc_hd__and2_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21405_ _08239_ _08240_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__nor2_1
XFILLER_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25173_ C_out\[413\] net101 net73 ser_C.shift_reg\[413\] _11056_ VGND VGND VPWR VPWR
+ _02663_ sky130_fd_sc_hd__a221o_1
X_22385_ _09125_ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__inv_2
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24124_ _10563_ systolic_inst.A_shift\[29\]\[1\] net71 VGND VGND VPWR VPWR _02107_
+ sky130_fd_sc_hd__mux2_1
X_21336_ _08187_ _08188_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__nand2_1
XFILLER_136_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24055_ systolic_inst.B_shift\[4\]\[7\] B_in\[7\] _00008_ VGND VGND VPWR VPWR _10545_
+ sky130_fd_sc_hd__mux2_1
X_28932_ clknet_leaf_265_clk _02730_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21267_ _08129_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__inv_2
XFILLER_104_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23006_ _09681_ _09682_ VGND VGND VPWR VPWR _09683_ sky130_fd_sc_hd__nand2_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20218_ net68 _07179_ _07180_ systolic_inst.acc_wires\[6\]\[30\] net106 VGND VGND
+ VPWR VPWR _01584_ sky130_fd_sc_hd__a32o_1
XFILLER_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28863_ clknet_leaf_332_clk _02661_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[411\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21198_ _08041_ _08065_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_161_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27814_ clknet_leaf_140_clk _01612_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_104_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20149_ _07100_ _07121_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__nor2_1
X_28794_ clknet_leaf_233_clk _02592_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_237_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27745_ clknet_leaf_213_clk _01543_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24957_ C_out\[305\] net103 net76 ser_C.shift_reg\[305\] _10948_ VGND VGND VPWR VPWR
+ _02555_ sky130_fd_sc_hd__a221o_1
X_14710_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[27\]
+ VGND VGND VPWR VPWR _11861_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23908_ systolic_inst.B_shift\[17\]\[6\] B_in\[78\] _00008_ VGND VGND VPWR VPWR _10487_
+ sky130_fd_sc_hd__mux2_1
XFILLER_233_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27676_ clknet_leaf_200_clk _01474_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15690_ _12672_ _12678_ _12708_ _12741_ _12707_ VGND VGND VPWR VPWR _12744_ sky130_fd_sc_hd__a311oi_4
XFILLER_45_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24888_ net110 ser_C.shift_reg\[272\] VGND VGND VPWR VPWR _10914_ sky130_fd_sc_hd__and2_1
X_29415_ clknet_leaf_328_clk _03213_ net136 VGND VGND VPWR VPWR C_out\[387\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26627_ clknet_leaf_20_B_in_serial_clk _00430_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14641_ _11801_ _11802_ VGND VGND VPWR VPWR _11803_ sky130_fd_sc_hd__nand2_1
XFILLER_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23839_ _10430_ _10431_ _10432_ VGND VGND VPWR VPWR _10434_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_159_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29346_ clknet_leaf_224_clk _03144_ net140 VGND VGND VPWR VPWR C_out\[318\] sky130_fd_sc_hd__dfrtp_1
X_17360_ systolic_inst.A_outs\[10\]\[2\] systolic_inst.B_outs\[10\]\[5\] _04580_ _04579_
+ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__a31oi_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14572_ _11743_ VGND VGND VPWR VPWR _11744_ sky130_fd_sc_hd__inv_2
X_26558_ clknet_leaf_2_A_in_serial_clk _00361_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_198_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16311_ _03689_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__xnor2_1
X_25509_ _11233_ _11235_ systolic_inst.cycle_cnt\[26\] VGND VGND VPWR VPWR _02820_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_955 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13523_ deser_A.shift_reg\[87\] deser_A.shift_reg\[88\] net129 VGND VGND VPWR VPWR
+ _00360_ sky130_fd_sc_hd__mux2_1
X_29277_ clknet_leaf_188_clk _03075_ net148 VGND VGND VPWR VPWR C_out\[249\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17291_ _04548_ _04549_ _04537_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__or3b_1
XFILLER_203_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26489_ clknet_leaf_8_A_in_serial_clk _00292_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_207_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19030_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[1\]
+ systolic_inst.B_outs\[7\]\[0\] VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__a22o_1
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28228_ clknet_leaf_47_clk _02026_ VGND VGND VPWR VPWR systolic_inst.B_shift\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16242_ net115 _03623_ _03624_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__and3_1
XFILLER_13_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13454_ deser_A.shift_reg\[18\] deser_A.shift_reg\[19\] deser_A.receiving VGND VGND
+ VPWR VPWR _00291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28159_ clknet_leaf_107_clk _01957_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_16173_ _03517_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__nor2_1
X_13385_ A_in\[94\] deser_A.word_buffer\[94\] net95 VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__mux2_1
XFILLER_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15124_ _12238_ _12239_ VGND VGND VPWR VPWR _12240_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_895 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19932_ _06927_ _06928_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__xnor2_1
X_15055_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[7\] _12144_ _12109_
+ VGND VGND VPWR VPWR _12173_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_71_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14006_ deser_B.shift_reg\[40\] deser_B.shift_reg\[41\] deser_B.receiving VGND VGND
+ VPWR VPWR _00832_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_220_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19863_ systolic_inst.A_outs\[6\]\[3\] systolic_inst.A_outs\[6\]\[4\] systolic_inst.B_outs\[6\]\[6\]
+ systolic_inst.B_outs\[6\]\[7\] VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_220_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_220_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18814_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__inv_2
X_19794_ systolic_inst.A_outs\[6\]\[2\] systolic_inst.B_outs\[6\]\[6\] _11278_ systolic_inst.A_outs\[6\]\[1\]
+ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18745_ _05839_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__xnor2_1
X_15957_ _12969_ _12973_ _12974_ net61 VGND VGND VPWR VPWR _12976_ sky130_fd_sc_hd__a31o_1
XFILLER_23_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14908_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[7\]
+ VGND VGND VPWR VPWR _12030_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_69_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18676_ _05695_ _05800_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__nand2_1
XFILLER_236_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15888_ _12914_ _12916_ _12917_ VGND VGND VPWR VPWR _12918_ sky130_fd_sc_hd__or3_1
XFILLER_188_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_218_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17627_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[10\]\[8\]
+ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__xnor2_1
X_14839_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[5\]
+ systolic_inst.A_outs\[14\]\[6\] VGND VGND VPWR VPWR _11963_ sky130_fd_sc_hd__and4_1
XFILLER_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17558_ _04807_ _04808_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__nor2_1
XFILLER_189_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16509_ _03863_ _03864_ _03860_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17489_ _04741_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19228_ _06254_ _06256_ _06290_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__nand3_1
XFILLER_20_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_227_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19159_ _06186_ _06188_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__and2b_1
XFILLER_30_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22170_ systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[5\] systolic_inst.A_outs\[2\]\[6\]
+ systolic_inst.B_outs\[2\]\[0\] VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__a22oi_1
XFILLER_173_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21121_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[4\]\[4\] systolic_inst.A_outs\[4\]\[7\]
+ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__o21a_1
XFILLER_236_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21052_ systolic_inst.A_outs\[4\]\[4\] systolic_inst.B_outs\[4\]\[5\] systolic_inst.A_outs\[4\]\[7\]
+ systolic_inst.B_outs\[4\]\[1\] VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__a22o_1
XFILLER_8_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20003_ _06995_ _06997_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__nand2_1
XFILLER_8_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25860_ systolic_inst.acc_wires\[10\]\[16\] C_out\[336\] net12 VGND VGND VPWR VPWR
+ _03162_ sky130_fd_sc_hd__mux2_1
XFILLER_28_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24811_ C_out\[232\] net99 net79 ser_C.shift_reg\[232\] _10875_ VGND VGND VPWR VPWR
+ _02482_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_203_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25791_ systolic_inst.acc_wires\[8\]\[11\] C_out\[267\] net29 VGND VGND VPWR VPWR
+ _03093_ sky130_fd_sc_hd__mux2_1
XFILLER_228_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27530_ clknet_leaf_243_clk _01328_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_24742_ net112 ser_C.shift_reg\[199\] VGND VGND VPWR VPWR _10841_ sky130_fd_sc_hd__and2_1
XFILLER_227_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21954_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[3\]\[13\]
+ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_19_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27461_ clknet_leaf_195_clk _01259_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_76_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20905_ systolic_inst.B_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[4\] systolic_inst.B_outs\[4\]\[5\]
+ systolic_inst.A_outs\[4\]\[0\] VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__a22o_1
XFILLER_215_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21885_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[3\]\[3\]
+ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__nand2_1
X_24673_ C_out\[163\] net103 net76 ser_C.shift_reg\[163\] _10806_ VGND VGND VPWR VPWR
+ _02413_ sky130_fd_sc_hd__a221o_1
XFILLER_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29200_ clknet_leaf_142_clk _02998_ net149 VGND VGND VPWR VPWR C_out\[172\] sky130_fd_sc_hd__dfrtp_1
XFILLER_242_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26412_ clknet_leaf_29_clk _00219_ net133 VGND VGND VPWR VPWR A_in\[80\] sky130_fd_sc_hd__dfrtp_1
X_23624_ _10205_ _10208_ _10243_ VGND VGND VPWR VPWR _10245_ sky130_fd_sc_hd__or3_1
X_20836_ systolic_inst.B_outs\[3\]\[1\] systolic_inst.B_shift\[3\]\[1\] net120 VGND
+ VGND VPWR VPWR _01659_ sky130_fd_sc_hd__mux2_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27392_ clknet_leaf_338_clk _01190_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_39_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29131_ clknet_leaf_169_clk _02929_ net148 VGND VGND VPWR VPWR C_out\[103\] sky130_fd_sc_hd__dfrtp_1
X_26343_ clknet_leaf_63_clk _00150_ net144 VGND VGND VPWR VPWR A_in\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_211_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20767_ systolic_inst.acc_wires\[5\]\[20\] systolic_inst.acc_wires\[5\]\[21\] systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__o21a_1
X_23555_ _10134_ _10136_ _10175_ _10177_ VGND VGND VPWR VPWR _10178_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_154_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29062_ clknet_leaf_108_clk _02860_ net150 VGND VGND VPWR VPWR C_out\[34\] sky130_fd_sc_hd__dfrtp_1
X_22506_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[2\]\[6\]
+ VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__nand2_1
X_23486_ _10105_ _10108_ VGND VGND VPWR VPWR _10110_ sky130_fd_sc_hd__xnor2_1
X_26274_ clknet_leaf_20_A_in_serial_clk _00082_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20698_ _07591_ _07614_ _07604_ _07613_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_126_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28013_ clknet_leaf_112_clk _01811_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_182_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22437_ _09148_ _09152_ VGND VGND VPWR VPWR _09177_ sky130_fd_sc_hd__nor2_1
X_25225_ C_out\[439\] net101 net73 ser_C.shift_reg\[439\] _11082_ VGND VGND VPWR VPWR
+ _02689_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_28_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13170_ deser_A.word_buffer\[8\] deser_A.serial_word\[8\] net127 VGND VGND VPWR VPWR
+ _00018_ sky130_fd_sc_hd__mux2_1
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22368_ _09093_ _09109_ VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__xor2_1
X_25156_ net110 ser_C.shift_reg\[406\] VGND VGND VPWR VPWR _11048_ sky130_fd_sc_hd__and2_1
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24107_ systolic_inst.B_shift\[1\]\[2\] _11332_ net83 systolic_inst.B_shift\[5\]\[2\]
+ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__a22o_1
XFILLER_151_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21319_ _08165_ _08169_ _08172_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__a21o_1
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25087_ C_out\[370\] net98 net78 ser_C.shift_reg\[370\] _11013_ VGND VGND VPWR VPWR
+ _02620_ sky130_fd_sc_hd__a221o_1
X_22299_ _09004_ _09005_ _09007_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__o21a_1
XFILLER_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24038_ _10536_ systolic_inst.B_shift\[4\]\[6\] _11332_ VGND VGND VPWR VPWR _02048_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28915_ clknet_leaf_282_clk _02713_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_105_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28846_ clknet_leaf_334_clk _02644_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[394\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16860_ _04169_ _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__nand2_1
X_15811_ net61 _12851_ VGND VGND VPWR VPWR _12852_ sky130_fd_sc_hd__nor2_1
XFILLER_237_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28777_ clknet_leaf_229_clk _02575_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[325\]
+ sky130_fd_sc_hd__dfrtp_1
X_16791_ _04101_ _04109_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__or2_1
XFILLER_111_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25989_ systolic_inst.acc_wires\[14\]\[17\] ser_C.parallel_data\[465\] net25 VGND
+ VGND VPWR VPWR _03291_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_37_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18530_ _05658_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__nand2_1
XFILLER_111_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27728_ clknet_leaf_140_clk _01526_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_15742_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[14\] _12793_ net115
+ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _05585_ _05592_ _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__and3_1
XFILLER_93_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15673_ _12694_ _12696_ _12726_ VGND VGND VPWR VPWR _12727_ sky130_fd_sc_hd__a21o_1
X_27659_ clknet_leaf_302_clk _01457_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_193_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_193_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17412_ _04665_ _04666_ _04667_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__a21oi_1
X_14624_ _11786_ _11787_ VGND VGND VPWR VPWR _11788_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_64_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _05536_ _05539_ _05543_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__o31a_1
XFILLER_18_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17343_ _04572_ _04574_ _04573_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__o21bai_1
X_29329_ clknet_leaf_221_clk _03127_ net139 VGND VGND VPWR VPWR C_out\[301\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14555_ _11722_ _11723_ _11721_ VGND VGND VPWR VPWR _11729_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13506_ deser_A.shift_reg\[70\] deser_A.shift_reg\[71\] net129 VGND VGND VPWR VPWR
+ _00343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17274_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[5\]
+ systolic_inst.A_outs\[10\]\[6\] VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_12_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14486_ _11666_ _11665_ VGND VGND VPWR VPWR _11667_ sky130_fd_sc_hd__and2b_1
XFILLER_31_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19013_ systolic_inst.A_outs\[7\]\[2\] systolic_inst.A_outs\[6\]\[2\] net119 VGND
+ VGND VPWR VPWR _01460_ sky130_fd_sc_hd__mux2_1
X_16225_ _03564_ _03572_ _03571_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__a21bo_1
XFILLER_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13437_ deser_A.shift_reg\[1\] deser_A.shift_reg\[2\] deser_A.receiving VGND VGND
+ VPWR VPWR _00274_ sky130_fd_sc_hd__mux2_1
Xclkload205 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload205/Y sky130_fd_sc_hd__clkinv_2
Xclkload216 clknet_leaf_44_clk VGND VGND VPWR VPWR clkload216/Y sky130_fd_sc_hd__inv_6
Xclkload227 clknet_leaf_71_clk VGND VGND VPWR VPWR clkload227/Y sky130_fd_sc_hd__clkinv_2
Xclkload238 clknet_leaf_87_clk VGND VGND VPWR VPWR clkload238/X sky130_fd_sc_hd__clkbuf_4
Xclkload249 clknet_leaf_125_clk VGND VGND VPWR VPWR clkload249/Y sky130_fd_sc_hd__clkinv_2
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16156_ _13094_ _03500_ _03499_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__o21a_1
X_13368_ A_in\[77\] deser_A.word_buffer\[77\] net96 VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15107_ _12222_ _12223_ VGND VGND VPWR VPWR _12224_ sky130_fd_sc_hd__nor2_1
XFILLER_138_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16087_ net108 _13082_ VGND VGND VPWR VPWR _13083_ sky130_fd_sc_hd__nor2_1
X_13299_ A_in\[8\] deser_A.word_buffer\[8\] net93 VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__mux2_1
XFILLER_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19915_ _06854_ _06912_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15038_ _12118_ _12120_ _12156_ VGND VGND VPWR VPWR _12157_ sky130_fd_sc_hd__a21o_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19846_ _06820_ _06845_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19777_ net106 _06776_ _06777_ _06778_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__o31ai_1
X_16989_ _04296_ _04297_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__a21o_1
XFILLER_83_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18728_ _05801_ _05851_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__xor2_1
XFILLER_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18659_ _05734_ _05751_ _05750_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_184_clk clknet_5_26__leaf_clk VGND VGND VPWR VPWR clknet_leaf_184_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21670_ _08477_ _08478_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__nor2_1
XFILLER_197_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_190_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_190_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20621_ net116 _07548_ _07549_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_211_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23340_ _09947_ _09966_ _09967_ VGND VGND VPWR VPWR _09968_ sky130_fd_sc_hd__nand3b_2
X_20552_ _07483_ _07484_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__or2_1
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23271_ _09909_ _09912_ VGND VGND VPWR VPWR _09914_ sky130_fd_sc_hd__or2_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20483_ _07415_ _07416_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22222_ _08931_ _08967_ VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__or2_1
XFILLER_146_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25010_ net111 ser_C.shift_reg\[333\] VGND VGND VPWR VPWR _10975_ sky130_fd_sc_hd__and2_1
XFILLER_192_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_209_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22153_ _08898_ _08900_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[3\]
+ VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_209_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21104_ _07959_ _07974_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__xor2_1
X_22084_ systolic_inst.A_outs\[2\]\[6\] systolic_inst.A_outs\[1\]\[6\] net122 VGND
+ VGND VPWR VPWR _01784_ sky130_fd_sc_hd__mux2_1
X_26961_ clknet_leaf_27_A_in_serial_clk _00759_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_205_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28700_ clknet_leaf_188_clk _02498_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[248\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25912_ systolic_inst.acc_wires\[12\]\[4\] C_out\[388\] net21 VGND VGND VPWR VPWR
+ _03214_ sky130_fd_sc_hd__mux2_1
X_21035_ _07864_ _07866_ _07906_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__and3_1
X_29680_ clknet_leaf_106_clk _03475_ net151 VGND VGND VPWR VPWR ser_C.bit_idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_26892_ clknet_leaf_7_A_in_serial_clk _00690_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28631_ clknet_leaf_205_clk _02429_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[179\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_143_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_197_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25843_ systolic_inst.acc_wires\[9\]\[31\] C_out\[319\] net13 VGND VGND VPWR VPWR
+ _03145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28562_ clknet_leaf_168_clk _02360_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25774_ systolic_inst.acc_wires\[7\]\[26\] C_out\[250\] net44 VGND VGND VPWR VPWR
+ _03076_ sky130_fd_sc_hd__mux2_1
XFILLER_216_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22986_ _09628_ _09630_ _09629_ VGND VGND VPWR VPWR _09663_ sky130_fd_sc_hd__o21ba_1
XFILLER_227_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27513_ clknet_leaf_226_clk _01311_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_24725_ C_out\[189\] net99 net79 ser_C.shift_reg\[189\] _10832_ VGND VGND VPWR VPWR
+ _02439_ sky130_fd_sc_hd__a221o_1
XFILLER_83_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_175_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_175_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_216_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28493_ clknet_leaf_117_clk _02291_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_21937_ _08726_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27444_ clknet_leaf_242_clk _01242_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24656_ net7 ser_C.shift_reg\[156\] VGND VGND VPWR VPWR _10798_ sky130_fd_sc_hd__and2_1
XFILLER_231_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21868_ net122 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[3\]\[0\]
+ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__a21oi_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23607_ _10226_ _10227_ VGND VGND VPWR VPWR _10228_ sky130_fd_sc_hd__nand2_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20819_ _07716_ _07717_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__nand2_1
X_27375_ clknet_leaf_327_clk _01173_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_24587_ C_out\[120\] net100 net82 ser_C.shift_reg\[120\] _10763_ VGND VGND VPWR VPWR
+ _02370_ sky130_fd_sc_hd__a221o_1
XFILLER_208_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21799_ _08551_ _08603_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__and2b_1
XFILLER_169_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29114_ clknet_leaf_157_clk _02912_ net151 VGND VGND VPWR VPWR C_out\[86\] sky130_fd_sc_hd__dfrtp_1
XFILLER_168_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14340_ systolic_inst.B_outs\[15\]\[3\] systolic_inst.B_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[5\]
+ systolic_inst.A_outs\[15\]\[6\] VGND VGND VPWR VPWR _11525_ sky130_fd_sc_hd__and4_1
X_26326_ clknet_leaf_30_A_in_serial_clk _00134_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_23538_ _10080_ _10122_ _10160_ VGND VGND VPWR VPWR _10161_ sky130_fd_sc_hd__o21a_1
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29045_ clknet_leaf_101_clk _02843_ net150 VGND VGND VPWR VPWR C_out\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14271_ _11417_ _11456_ VGND VGND VPWR VPWR _11458_ sky130_fd_sc_hd__or2_1
X_26257_ clknet_leaf_4_A_in_serial_clk _00065_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_23469_ _10050_ _10052_ _10091_ _10093_ VGND VGND VPWR VPWR _10094_ sky130_fd_sc_hd__a211oi_2
XFILLER_109_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16010_ _13004_ _13007_ VGND VGND VPWR VPWR _13008_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25208_ net110 ser_C.shift_reg\[432\] VGND VGND VPWR VPWR _11074_ sky130_fd_sc_hd__and2_1
XFILLER_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13222_ deser_A.word_buffer\[60\] deser_A.serial_word\[60\] net128 VGND VGND VPWR
+ VPWR _00070_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26188_ ser_C.bit_idx\[5\] ser_C.bit_idx\[6\] _11250_ VGND VGND VPWR VPWR _11254_
+ sky130_fd_sc_hd__and3_1
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13153_ net1 deser_A.receiving VGND VGND VPWR VPWR _11304_ sky130_fd_sc_hd__nor2_1
X_25139_ C_out\[396\] net101 net73 ser_C.shift_reg\[396\] _11039_ VGND VGND VPWR VPWR
+ _02646_ sky130_fd_sc_hd__a221o_1
XFILLER_139_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17961_ _05147_ _05153_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19700_ _06675_ _06703_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__nand2_1
X_16912_ systolic_inst.A_outs\[11\]\[6\] _11262_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__or2_1
X_17892_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[4\] VGND VGND VPWR
+ VPWR _05087_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19631_ systolic_inst.A_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[1\]
+ systolic_inst.B_outs\[6\]\[0\] VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__a22o_1
X_16843_ net105 _04160_ _04161_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_105_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28829_ clknet_leaf_195_clk _02627_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[377\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1007 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19562_ _06574_ _06581_ _06586_ _06591_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_66_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16774_ _04057_ _04093_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__nor2_1
XFILLER_111_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13986_ deser_B.shift_reg\[20\] deser_B.shift_reg\[21\] net125 VGND VGND VPWR VPWR
+ _00812_ sky130_fd_sc_hd__mux2_1
XFILLER_46_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18513_ _05641_ _05642_ _05612_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_215_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15725_ _12775_ _12776_ VGND VGND VPWR VPWR _12777_ sky130_fd_sc_hd__or2_1
XFILLER_80_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19493_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[7\]\[12\]
+ _06534_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_166_clk clknet_5_31__leaf_clk VGND VGND VPWR VPWR clknet_leaf_166_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_234_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18444_ _05564_ _05566_ _05577_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__and3_1
XFILLER_221_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15656_ _12672_ _12678_ _12709_ VGND VGND VPWR VPWR _12711_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_199_Right_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14607_ _11756_ _11772_ VGND VGND VPWR VPWR _11773_ sky130_fd_sc_hd__nor2_1
X_18375_ _05531_ _05532_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__xnor2_1
X_15587_ _12616_ _12617_ _12618_ VGND VGND VPWR VPWR _12643_ sky130_fd_sc_hd__o21ba_1
XFILLER_57_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17326_ _04576_ _04582_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14538_ _11711_ net69 _11714_ systolic_inst.acc_wires\[15\]\[1\] net107 VGND VGND
+ VPWR VPWR _00979_ sky130_fd_sc_hd__a32o_1
XFILLER_175_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17257_ _04514_ _04515_ _04513_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__a21o_1
XFILLER_128_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14469_ systolic_inst.B_outs\[15\]\[6\] systolic_inst.A_outs\[15\]\[7\] VGND VGND
+ VPWR VPWR _11650_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_42_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16208_ _03517_ _03589_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_96_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17188_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.B_outs\[5\]\[2\] net116 VGND
+ VGND VPWR VPWR _01276_ sky130_fd_sc_hd__mux2_1
X_16139_ _03522_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__nor2_1
XFILLER_115_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_241_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19829_ _06825_ _06828_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__xnor2_1
XFILLER_233_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22840_ systolic_inst.B_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[4\]
+ systolic_inst.A_outs\[1\]\[5\] VGND VGND VPWR VPWR _09521_ sky130_fd_sc_hd__and4_1
XFILLER_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_157_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_157_clk
+ sky130_fd_sc_hd__clkbuf_8
X_22771_ _09449_ _09452_ VGND VGND VPWR VPWR _09454_ sky130_fd_sc_hd__xnor2_1
X_24510_ net112 ser_C.shift_reg\[83\] VGND VGND VPWR VPWR _10725_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21722_ _08526_ _08527_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_49_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25490_ _11222_ _11224_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__and2_1
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24441_ C_out\[47\] _11302_ net81 ser_C.shift_reg\[47\] _10690_ VGND VGND VPWR VPWR
+ _02297_ sky130_fd_sc_hd__a221o_1
X_21653_ _08452_ _08460_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__xnor2_1
XFILLER_220_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20604_ _07533_ _07534_ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__nor2_1
XFILLER_166_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27160_ clknet_leaf_297_clk _00958_ net138 VGND VGND VPWR VPWR systolic_inst.B_outs\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_24372_ net7 ser_C.shift_reg\[14\] VGND VGND VPWR VPWR _10656_ sky130_fd_sc_hd__and2_1
X_21584_ _08350_ _08352_ _08394_ VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__a21oi_1
XFILLER_178_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26111_ deser_B.serial_word\[66\] deser_B.shift_reg\[66\] _00001_ VGND VGND VPWR
+ VPWR _03413_ sky130_fd_sc_hd__mux2_1
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23323_ _09945_ _09947_ _09950_ _09951_ VGND VGND VPWR VPWR _09952_ sky130_fd_sc_hd__nand4_1
XFILLER_165_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20535_ _07466_ _07467_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__nor2_1
XFILLER_123_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27091_ clknet_leaf_5_B_in_serial_clk _00889_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26042_ systolic_inst.B_outs\[15\]\[6\] systolic_inst.B_outs\[11\]\[6\] net118 VGND
+ VGND VPWR VPWR _03344_ sky130_fd_sc_hd__mux2_1
X_23254_ _09883_ _09885_ _09897_ _09898_ _09891_ VGND VGND VPWR VPWR _09899_ sky130_fd_sc_hd__a311oi_4
XFILLER_197_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20466_ systolic_inst.B_outs\[5\]\[5\] systolic_inst.A_outs\[5\]\[5\] VGND VGND VPWR
+ VPWR _07401_ sky130_fd_sc_hd__nand2_1
XFILLER_146_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_207_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22205_ _11265_ _08950_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__xnor2_1
X_23185_ _09840_ VGND VGND VPWR VPWR _09841_ sky130_fd_sc_hd__inv_2
X_20397_ systolic_inst.A_outs\[5\]\[2\] systolic_inst.B_outs\[5\]\[6\] VGND VGND VPWR
+ VPWR _07334_ sky130_fd_sc_hd__nand2_1
XFILLER_134_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22136_ _08882_ _08883_ _08876_ VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_145_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27993_ clknet_leaf_123_clk _01791_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_160_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22067_ net65 _08837_ _08838_ systolic_inst.acc_wires\[3\]\[29\] net106 VGND VGND
+ VPWR VPWR _01775_ sky130_fd_sc_hd__a32o_1
X_26944_ clknet_leaf_20_A_in_serial_clk _00742_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21018_ _07850_ _07889_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29663_ clknet_leaf_10_B_in_serial_clk _03458_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_26875_ clknet_leaf_13_A_in_serial_clk _00673_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28614_ clknet_leaf_218_clk _02412_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[162\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_210_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13840_ deser_A.serial_word\[1\] deser_A.shift_reg\[1\] net58 VGND VGND VPWR VPWR
+ _00666_ sky130_fd_sc_hd__mux2_1
XFILLER_101_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25826_ systolic_inst.acc_wires\[9\]\[14\] C_out\[302\] net15 VGND VGND VPWR VPWR
+ _03128_ sky130_fd_sc_hd__mux2_1
X_29594_ clknet_leaf_13_B_in_serial_clk _03389_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28545_ clknet_leaf_164_clk _02343_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13771_ B_in\[78\] deser_B.word_buffer\[78\] net86 VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_148_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_148_clk
+ sky130_fd_sc_hd__clkbuf_8
X_25757_ systolic_inst.acc_wires\[7\]\[9\] C_out\[233\] net42 VGND VGND VPWR VPWR
+ _03059_ sky130_fd_sc_hd__mux2_1
X_22969_ _09609_ _09611_ _09646_ VGND VGND VPWR VPWR _09647_ sky130_fd_sc_hd__and3_1
XFILLER_128_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15510_ _12537_ _12568_ VGND VGND VPWR VPWR _12569_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24708_ net113 ser_C.shift_reg\[182\] VGND VGND VPWR VPWR _10824_ sky130_fd_sc_hd__and2_1
XFILLER_71_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28476_ clknet_leaf_107_clk _02274_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_188_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16490_ net67 _03848_ _03849_ systolic_inst.acc_wires\[12\]\[17\] net108 VGND VGND
+ VPWR VPWR _01187_ sky130_fd_sc_hd__a32o_1
X_25688_ systolic_inst.acc_wires\[5\]\[4\] C_out\[164\] net16 VGND VGND VPWR VPWR
+ _02990_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15441_ _12482_ _12500_ VGND VGND VPWR VPWR _12502_ sky130_fd_sc_hd__xnor2_1
X_27427_ clknet_leaf_249_clk _01225_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_175_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24639_ C_out\[146\] net104 net76 ser_C.shift_reg\[146\] _10789_ VGND VGND VPWR VPWR
+ _02396_ sky130_fd_sc_hd__a221o_1
XFILLER_230_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18160_ systolic_inst.B_outs\[9\]\[5\] systolic_inst.A_outs\[9\]\[7\] _05324_ _05323_
+ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__a31o_1
X_27358_ clknet_leaf_322_clk _01156_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_15372_ net116 systolic_inst.B_outs\[13\]\[0\] systolic_inst.A_outs\[13\]\[0\] VGND
+ VGND VPWR VPWR _12438_ sky130_fd_sc_hd__and3_1
XFILLER_180_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17111_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__inv_2
X_26309_ clknet_leaf_24_A_in_serial_clk _00117_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_14323_ _11506_ _11507_ VGND VGND VPWR VPWR _11509_ sky130_fd_sc_hd__xor2_1
XFILLER_183_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18091_ _05220_ _05280_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_320_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_320_clk
+ sky130_fd_sc_hd__clkbuf_8
X_27289_ clknet_leaf_319_clk _01087_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_59_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29028_ clknet_leaf_128_clk _02826_ net144 VGND VGND VPWR VPWR C_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_17042_ _04342_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__nand2_1
X_14254_ systolic_inst.B_outs\[15\]\[7\] _11438_ _11440_ VGND VGND VPWR VPWR _11441_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_130_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap119 systolic_inst.ce_local VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_130_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13205_ deser_A.word_buffer\[43\] deser_A.serial_word\[43\] net127 VGND VGND VPWR
+ VPWR _00053_ sky130_fd_sc_hd__mux2_1
XFILLER_136_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14185_ _11354_ _11356_ _11374_ VGND VGND VPWR VPWR _11375_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_91_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13136_ systolic_inst.cycle_cnt\[1\] systolic_inst.cycle_cnt\[2\] systolic_inst.cycle_cnt\[3\]
+ VGND VGND VPWR VPWR _11289_ sky130_fd_sc_hd__o21a_1
XFILLER_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18993_ net108 systolic_inst.acc_wires\[8\]\[28\] net66 _06085_ VGND VGND VPWR VPWR
+ _01454_ sky130_fd_sc_hd__a22o_1
XFILLER_61_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17944_ _05135_ _05136_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__xnor2_1
XFILLER_238_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17875_ _05041_ _05070_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__nand2_1
XFILLER_239_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19614_ systolic_inst.A_outs\[6\]\[2\] systolic_inst.A_outs\[5\]\[2\] net120 VGND
+ VGND VPWR VPWR _01524_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16826_ _04108_ _04110_ _04144_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__a21o_1
XFILLER_24_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19545_ _06580_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__inv_2
XFILLER_59_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16757_ _04075_ _04076_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__xor2_1
XFILLER_94_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13969_ deser_B.shift_reg\[3\] deser_B.shift_reg\[4\] net125 VGND VGND VPWR VPWR
+ _00795_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_139_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15708_ _12715_ _12729_ _12727_ VGND VGND VPWR VPWR _12761_ sky130_fd_sc_hd__o21a_1
XFILLER_206_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19476_ _06520_ _06521_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__nand2_1
X_16688_ _03987_ _04009_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_234_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_234_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15639_ _12693_ _12692_ VGND VGND VPWR VPWR _12694_ sky130_fd_sc_hd__nand2b_1
X_18427_ systolic_inst.B_outs\[8\]\[0\] systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[1\]
+ systolic_inst.A_outs\[8\]\[2\] VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__and4_1
XFILLER_94_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18358_ _05517_ _05518_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__or2_1
XFILLER_175_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17309_ _04564_ _04565_ systolic_inst.B_outs\[10\]\[7\] VGND VGND VPWR VPWR _04567_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18289_ _05454_ _05459_ _05458_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__a21o_1
XFILLER_147_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_311_clk clknet_5_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_311_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20320_ _07258_ _07255_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__nand2b_1
XFILLER_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20251_ systolic_inst.A_outs\[5\]\[0\] systolic_inst.B_outs\[5\]\[2\] _07193_ VGND
+ VGND VPWR VPWR _07194_ sky130_fd_sc_hd__nand3_1
XFILLER_190_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_181_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20182_ net106 systolic_inst.acc_wires\[6\]\[24\] net62 _07150_ VGND VGND VPWR VPWR
+ _01578_ sky130_fd_sc_hd__a22o_1
XFILLER_142_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24990_ net111 ser_C.shift_reg\[323\] VGND VGND VPWR VPWR _10965_ sky130_fd_sc_hd__and2_1
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_235_Right_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23941_ _10499_ systolic_inst.B_shift\[10\]\[2\] _11332_ VGND VGND VPWR VPWR _01988_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26660_ clknet_leaf_2_B_in_serial_clk _00463_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_23872_ systolic_inst.acc_wires\[0\]\[26\] systolic_inst.acc_wires\[0\]\[27\] systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _10461_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_179_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25611_ systolic_inst.acc_wires\[2\]\[23\] C_out\[87\] net52 VGND VGND VPWR VPWR
+ _02913_ sky130_fd_sc_hd__mux2_1
X_22823_ _09453_ _09455_ _09503_ _09504_ VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__a211oi_1
X_26591_ clknet_leaf_30_A_in_serial_clk _00394_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28330_ clknet_leaf_2_clk _02128_ VGND VGND VPWR VPWR systolic_inst.A_shift\[27\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25542_ systolic_inst.acc_wires\[0\]\[18\] C_out\[18\] net54 VGND VGND VPWR VPWR
+ _02844_ sky130_fd_sc_hd__mux2_1
XFILLER_198_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22754_ _09427_ _09437_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__nor2_1
XFILLER_241_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21705_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[9\] VGND
+ VGND VPWR VPWR _08513_ sky130_fd_sc_hd__and2_1
X_28261_ clknet_leaf_57_clk _02059_ VGND VGND VPWR VPWR systolic_inst.B_shift\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25473_ systolic_inst.cycle_cnt\[12\] _11306_ _11206_ systolic_inst.cycle_cnt\[13\]
+ VGND VGND VPWR VPWR _11213_ sky130_fd_sc_hd__a31o_1
XFILLER_129_1377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22685_ systolic_inst.B_outs\[0\]\[4\] systolic_inst.B_shift\[0\]\[4\] net121 VGND
+ VGND VPWR VPWR _01854_ sky130_fd_sc_hd__mux2_1
XFILLER_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27212_ clknet_leaf_292_clk _01010_ net139 VGND VGND VPWR VPWR systolic_inst.A_outs\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_24424_ net114 ser_C.shift_reg\[40\] VGND VGND VPWR VPWR _10682_ sky130_fd_sc_hd__and2_1
XFILLER_139_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21636_ _08444_ _08441_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__and2b_1
X_28192_ clknet_leaf_129_clk _01990_ VGND VGND VPWR VPWR systolic_inst.B_shift\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_170_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27143_ clknet_leaf_7_clk _00941_ VGND VGND VPWR VPWR systolic_inst.A_shift\[21\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24355_ C_out\[4\] net104 _10643_ ser_C.shift_reg\[4\] _10647_ VGND VGND VPWR VPWR
+ _02254_ sky130_fd_sc_hd__a221o_1
XFILLER_165_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21567_ _08348_ _08377_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__and2_1
XFILLER_139_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_302_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_302_clk
+ sky130_fd_sc_hd__clkbuf_8
X_23306_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[3\] VGND VGND VPWR
+ VPWR _09936_ sky130_fd_sc_hd__nand2_1
XFILLER_60_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27074_ clknet_leaf_11_B_in_serial_clk _00872_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_20518_ _07449_ _07450_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__and2b_1
XFILLER_193_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21498_ _08310_ _08311_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__or2_1
X_24286_ _10616_ systolic_inst.B_shift\[23\]\[6\] net72 VGND VGND VPWR VPWR _02216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26025_ systolic_inst.acc_wires\[15\]\[21\] ser_C.parallel_data\[501\] net37 VGND
+ VGND VPWR VPWR _03327_ sky130_fd_sc_hd__mux2_1
X_23237_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[25\]
+ VGND VGND VPWR VPWR _09885_ sky130_fd_sc_hd__xor2_2
X_20449_ _07382_ _07383_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23168_ _09822_ _09825_ VGND VGND VPWR VPWR _09827_ sky130_fd_sc_hd__or2_1
XFILLER_162_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22119_ _08855_ _08857_ _08868_ VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__and3_1
X_27976_ clknet_leaf_172_clk _01774_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_23099_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[1\]\[5\]
+ VGND VGND VPWR VPWR _09767_ sky130_fd_sc_hd__nand2_1
X_15990_ net115 _12987_ _12988_ _12989_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__a31o_1
XFILLER_212_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14941_ _12059_ _12060_ VGND VGND VPWR VPWR _12063_ sky130_fd_sc_hd__nand2_1
XFILLER_88_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26927_ clknet_leaf_5_A_in_serial_clk _00725_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_202_Right_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17660_ _04895_ _04896_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__nor2_1
X_26858_ clknet_leaf_0_B_in_serial_clk _00660_ net134 VGND VGND VPWR VPWR deser_B.bit_idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_29646_ clknet_leaf_33_B_in_serial_clk _03441_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_14872_ _11993_ _11994_ VGND VGND VPWR VPWR _11995_ sky130_fd_sc_hd__nand2_1
XFILLER_236_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16611_ _03926_ _03935_ _03936_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__nand3_1
X_13823_ deser_B.bit_idx\[1\] _11319_ VGND VGND VPWR VPWR _11320_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_123_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25809_ systolic_inst.acc_wires\[8\]\[29\] C_out\[285\] net27 VGND VGND VPWR VPWR
+ _03111_ sky130_fd_sc_hd__mux2_1
XFILLER_217_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29577_ clknet_leaf_23_B_in_serial_clk _03372_ net137 VGND VGND VPWR VPWR deser_B.serial_word\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17591_ _11712_ _04835_ _04837_ systolic_inst.acc_wires\[10\]\[2\] net107 VGND VGND
+ VPWR VPWR _01300_ sky130_fd_sc_hd__a32o_1
X_26789_ clknet_leaf_69_clk _00591_ net153 VGND VGND VPWR VPWR B_in\[61\] sky130_fd_sc_hd__dfrtp_1
XFILLER_235_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28528_ clknet_leaf_166_clk _02326_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19330_ _06390_ _06389_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__and2b_1
XFILLER_141_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16542_ _03891_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__and2_1
XFILLER_204_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13754_ B_in\[61\] deser_B.word_buffer\[61\] net87 VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__mux2_1
XFILLER_1_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19261_ _06281_ _06289_ _06288_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__a21bo_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28459_ clknet_leaf_124_clk _02257_ net144 VGND VGND VPWR VPWR ser_C.shift_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_16473_ _03826_ _03831_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13685_ deser_B.word_buffer\[121\] deser_B.serial_word\[121\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18212_ _05384_ _05388_ _05391_ _05392_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__o211a_1
XFILLER_176_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15424_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[4\]
+ systolic_inst.A_outs\[13\]\[5\] VGND VGND VPWR VPWR _12485_ sky130_fd_sc_hd__and4_1
XFILLER_54_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19192_ _06247_ _06255_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18143_ _05329_ _05330_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__nand2_1
X_15355_ _12437_ _12436_ systolic_inst.acc_wires\[14\]\[31\] net107 VGND VGND VPWR
+ VPWR _01073_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_184_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ _11487_ _11491_ VGND VGND VPWR VPWR _11492_ sky130_fd_sc_hd__xnor2_1
X_18074_ systolic_inst.A_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[5\] systolic_inst.B_outs\[9\]\[6\]
+ systolic_inst.B_outs\[9\]\[7\] VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__and4b_1
XFILLER_157_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15286_ _12375_ _12377_ _12378_ VGND VGND VPWR VPWR _12380_ sky130_fd_sc_hd__or3_1
XFILLER_32_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_242_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17025_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[11\]\[9\]
+ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__xor2_1
XFILLER_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14237_ _11395_ _11423_ _11424_ VGND VGND VPWR VPWR _11425_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_242_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14168_ net118 _11356_ _11357_ _11358_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__a31o_1
XFILLER_28_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13119_ systolic_inst.B_outs\[10\]\[7\] VGND VGND VPWR VPWR _11275_ sky130_fd_sc_hd__inv_2
XFILLER_140_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14099_ net133 net59 VGND VGND VPWR VPWR _11333_ sky130_fd_sc_hd__and2_4
X_18976_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[26\]
+ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__nand2_1
XFILLER_26_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17927_ systolic_inst.A_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[4\]
+ systolic_inst.B_outs\[9\]\[3\] VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_33_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17858_ _05052_ _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_236_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_236_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16809_ _04057_ _04127_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__nor2_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17789_ systolic_inst.A_outs\[9\]\[4\] systolic_inst.A_outs\[8\]\[4\] net117 VGND
+ VGND VPWR VPWR _01334_ sky130_fd_sc_hd__mux2_1
XFILLER_241_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19528_ _06557_ _06559_ _06566_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_46_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_22__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_5_22__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_241_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19459_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[7\]\[9\]
+ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__xor2_1
XFILLER_50_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22470_ net122 _09205_ _09206_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__a21oi_1
XFILLER_195_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_187_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21421_ _08256_ _08258_ _08261_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__a21oi_2
XFILLER_202_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21352_ _08199_ _08201_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__or2_1
XFILLER_120_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24140_ _10571_ systolic_inst.A_shift\[28\]\[1\] net70 VGND VGND VPWR VPWR _02115_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20303_ _07241_ _07242_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__or2_1
XFILLER_198_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24071_ systolic_inst.B_shift\[19\]\[7\] B_in\[31\] _00008_ VGND VGND VPWR VPWR _10553_
+ sky130_fd_sc_hd__mux2_1
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21283_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[4\]\[5\]
+ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__and2_1
XFILLER_144_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23022_ _09696_ _09697_ VGND VGND VPWR VPWR _09698_ sky130_fd_sc_hd__nand2b_1
X_20234_ systolic_inst.B_outs\[4\]\[3\] systolic_inst.B_outs\[0\]\[3\] net117 VGND
+ VGND VPWR VPWR _01597_ sky130_fd_sc_hd__mux2_1
XFILLER_144_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27830_ clknet_leaf_141_clk _01628_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20165_ _07132_ _07133_ _07134_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__or3_1
XFILLER_58_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27761_ clknet_leaf_212_clk _01559_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20096_ _07073_ _07074_ _07075_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__a21oi_1
X_24973_ C_out\[313\] net103 net76 ser_C.shift_reg\[313\] _10956_ VGND VGND VPWR VPWR
+ _02563_ sky130_fd_sc_hd__a221o_1
XFILLER_170_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26712_ clknet_leaf_26_B_in_serial_clk _00515_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_29500_ clknet_leaf_268_clk _03298_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[472\]
+ sky130_fd_sc_hd__dfrtp_1
X_23924_ systolic_inst.B_shift\[22\]\[6\] B_in\[86\] net59 VGND VGND VPWR VPWR _10495_
+ sky130_fd_sc_hd__mux2_1
X_27692_ clknet_leaf_200_clk _01490_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29431_ clknet_leaf_337_clk _03229_ net131 VGND VGND VPWR VPWR C_out\[403\] sky130_fd_sc_hd__dfrtp_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26643_ clknet_leaf_14_B_in_serial_clk _00446_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_23855_ _10447_ _10446_ systolic_inst.acc_wires\[0\]\[24\] _11258_ VGND VGND VPWR
+ VPWR _01954_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22806_ systolic_inst.B_outs\[1\]\[3\] systolic_inst.A_outs\[1\]\[4\] VGND VGND VPWR
+ VPWR _09488_ sky130_fd_sc_hd__nand2_1
X_29362_ clknet_leaf_226_clk _03160_ net140 VGND VGND VPWR VPWR C_out\[334\] sky130_fd_sc_hd__dfrtp_1
XFILLER_226_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26574_ clknet_leaf_25_A_in_serial_clk _00377_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_23786_ _10387_ _10388_ VGND VGND VPWR VPWR _10389_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_172_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20998_ _07871_ _07870_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[7\]
+ net108 VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_214_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28313_ clknet_leaf_8_clk _02111_ VGND VGND VPWR VPWR systolic_inst.A_shift\[29\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_25525_ systolic_inst.acc_wires\[0\]\[1\] C_out\[1\] net32 VGND VGND VPWR VPWR _02827_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22737_ _09421_ _09420_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[4\]
+ _11258_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__a2bb2o_1
X_29293_ clknet_leaf_314_clk _03091_ net142 VGND VGND VPWR VPWR C_out\[265\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28244_ clknet_leaf_77_clk _02042_ VGND VGND VPWR VPWR systolic_inst.B_shift\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25456_ _11198_ _11201_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__and2_1
X_13470_ deser_A.shift_reg\[34\] deser_A.shift_reg\[35\] deser_A.receiving VGND VGND
+ VPWR VPWR _00307_ sky130_fd_sc_hd__mux2_1
XFILLER_231_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22668_ net65 _09373_ _09374_ systolic_inst.acc_wires\[2\]\[30\] net109 VGND VGND
+ VPWR VPWR _01840_ sky130_fd_sc_hd__a32o_1
XFILLER_185_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24407_ C_out\[30\] _11302_ net81 ser_C.shift_reg\[30\] _10673_ VGND VGND VPWR VPWR
+ _02280_ sky130_fd_sc_hd__a221o_1
XFILLER_142_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21619_ _08412_ _08428_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__xnor2_1
X_28175_ clknet_leaf_75_clk _01973_ VGND VGND VPWR VPWR systolic_inst.B_shift\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25387_ systolic_inst.A_shift\[3\]\[1\] A_in\[17\] net59 VGND VGND VPWR VPWR _11163_
+ sky130_fd_sc_hd__mux2_1
X_22599_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[20\]
+ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__xor2_1
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15140_ _12177_ _12240_ _12238_ VGND VGND VPWR VPWR _12255_ sky130_fd_sc_hd__a21oi_1
X_27126_ clknet_leaf_17_clk _00924_ VGND VGND VPWR VPWR systolic_inst.A_shift\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24338_ systolic_inst.A_shift\[8\]\[1\] net70 net83 systolic_inst.A_shift\[9\]\[1\]
+ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__a22o_1
X_27057_ clknet_leaf_1_B_in_serial_clk _00855_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_15071_ _12153_ _12155_ _12187_ VGND VGND VPWR VPWR _12189_ sky130_fd_sc_hd__nand3_1
X_24269_ systolic_inst.B_shift\[17\]\[4\] net72 _11333_ B_in\[108\] VGND VGND VPWR
+ VPWR _02206_ sky130_fd_sc_hd__a22o_1
XFILLER_142_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14022_ deser_B.shift_reg\[56\] deser_B.shift_reg\[57\] net125 VGND VGND VPWR VPWR
+ _00848_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26008_ systolic_inst.acc_wires\[15\]\[4\] ser_C.parallel_data\[484\] net23 VGND
+ VGND VPWR VPWR _03310_ sky130_fd_sc_hd__mux2_1
XFILLER_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18830_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[8\]\[5\]
+ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15973_ systolic_inst.B_outs\[11\]\[6\] systolic_inst.B_outs\[7\]\[6\] net119 VGND
+ VGND VPWR VPWR _01152_ sky130_fd_sc_hd__mux2_1
X_18761_ _05850_ _05852_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__o21a_1
X_27959_ clknet_leaf_170_clk _01757_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _04919_ _04940_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__nor2_1
X_14924_ systolic_inst.A_outs\[14\]\[2\] systolic_inst.B_outs\[14\]\[5\] _12009_ _12008_
+ VGND VGND VPWR VPWR _12046_ sky130_fd_sc_hd__a31oi_1
XFILLER_62_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18692_ _05777_ _05779_ _05816_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_121_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29629_ clknet_leaf_9_B_in_serial_clk _03424_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_14855_ _11973_ _11977_ VGND VGND VPWR VPWR _11979_ sky130_fd_sc_hd__xor2_1
X_17643_ _04878_ _04880_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13806_ B_in\[113\] deser_B.word_buffer\[113\] net88 VGND VGND VPWR VPWR _00643_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17574_ net105 systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] _04816_
+ _04823_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__a22o_1
X_14786_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[3\] _11912_ net118
+ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_231_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_231_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19313_ _06237_ _06372_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__nand2_2
XFILLER_147_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16525_ _03871_ _03875_ _03877_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__a21oi_1
X_13737_ B_in\[44\] deser_B.word_buffer\[44\] net84 VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__mux2_1
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_143_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19244_ _06238_ _06305_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_119_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16456_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[12\]\[13\]
+ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__nand2_1
XFILLER_32_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13668_ deser_B.word_buffer\[104\] deser_B.serial_word\[104\] net123 VGND VGND VPWR
+ VPWR _00505_ sky130_fd_sc_hd__mux2_1
XFILLER_177_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15407_ systolic_inst.B_outs\[13\]\[0\] systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[3\]
+ VGND VGND VPWR VPWR _12469_ sky130_fd_sc_hd__and3_1
XFILLER_176_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19175_ _06239_ _06236_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_26_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16387_ _03760_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__inv_2
X_13599_ deser_B.word_buffer\[35\] deser_B.serial_word\[35\] net123 VGND VGND VPWR
+ VPWR _00436_ sky130_fd_sc_hd__mux2_1
XFILLER_185_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18126_ _05313_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_229_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15338_ net107 systolic_inst.acc_wires\[14\]\[28\] _11712_ _12423_ VGND VGND VPWR
+ VPWR _01070_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_229_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18057_ _05186_ _05211_ _05210_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__a21boi_2
X_15269_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[18\]
+ VGND VGND VPWR VPWR _12365_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_225_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17008_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[11\]\[6\]
+ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__or2_1
XFILLER_99_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18959_ _06048_ _06052_ _06055_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__a21o_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21970_ _08748_ _08751_ _08754_ net60 VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_176_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20921_ _07793_ _07794_ _07795_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__o21bai_1
XFILLER_187_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23640_ _10080_ _10230_ _10259_ VGND VGND VPWR VPWR _10260_ sky130_fd_sc_hd__o21a_1
XFILLER_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1087 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20852_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[2\] _07728_ _07730_
+ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__and4_1
XFILLER_148_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23571_ _10154_ _10192_ VGND VGND VPWR VPWR _10193_ sky130_fd_sc_hd__nor2_1
XFILLER_81_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20783_ _07686_ _07687_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__or2_1
XFILLER_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
X_25310_ net111 ser_C.shift_reg\[483\] VGND VGND VPWR VPWR _11125_ sky130_fd_sc_hd__and2_1
X_22522_ _09248_ _09249_ net65 VGND VGND VPWR VPWR _09251_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26290_ clknet_leaf_2_A_in_serial_clk _00098_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_214_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25241_ ser_C.parallel_data\[447\] net102 net74 ser_C.shift_reg\[447\] _11090_ VGND
+ VGND VPWR VPWR _02697_ sky130_fd_sc_hd__a221o_1
XFILLER_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22453_ _09190_ _09191_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__nor2_1
XFILLER_148_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21404_ systolic_inst.acc_wires\[4\]\[20\] systolic_inst.acc_wires\[4\]\[21\] systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__o21a_1
XFILLER_136_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25172_ net110 ser_C.shift_reg\[414\] VGND VGND VPWR VPWR _11056_ sky130_fd_sc_hd__and2_1
X_22384_ _09123_ _09124_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__nand2_1
XFILLER_159_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24123_ systolic_inst.A_shift\[30\]\[1\] A_in\[113\] net59 VGND VGND VPWR VPWR _10563_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21335_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[4\]\[12\]
+ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__nand2_1
XFILLER_11_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24054_ _10544_ systolic_inst.B_shift\[0\]\[6\] _11332_ VGND VGND VPWR VPWR _02056_
+ sky130_fd_sc_hd__mux2_1
X_28931_ clknet_leaf_265_clk _02729_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[479\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21266_ _08119_ _08122_ _08126_ _08127_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__o211a_1
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23005_ _09614_ _09619_ _09648_ _09647_ VGND VGND VPWR VPWR _09682_ sky130_fd_sc_hd__a31o_1
XFILLER_173_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20217_ _07175_ _07178_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__or2_1
XFILLER_104_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21197_ _08063_ _08064_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__xnor2_1
X_28862_ clknet_leaf_332_clk _02660_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[410\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20148_ _07101_ _07106_ _07111_ _07115_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__or4_1
X_27813_ clknet_leaf_140_clk _01611_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_28793_ clknet_leaf_233_clk _02591_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[341\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20079_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[6\]\[9\]
+ _07057_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__a21oi_1
X_27744_ clknet_leaf_212_clk _01542_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24956_ net111 ser_C.shift_reg\[306\] VGND VGND VPWR VPWR _10948_ sky130_fd_sc_hd__and2_1
XFILLER_44_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23907_ _10486_ systolic_inst.B_shift\[13\]\[5\] net72 VGND VGND VPWR VPWR _01967_
+ sky130_fd_sc_hd__mux2_1
X_27675_ clknet_leaf_141_clk _01473_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_57_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24887_ C_out\[270\] net103 net75 ser_C.shift_reg\[270\] _10913_ VGND VGND VPWR VPWR
+ _02520_ sky130_fd_sc_hd__a221o_1
XFILLER_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26626_ clknet_leaf_23_B_in_serial_clk _00429_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14640_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[16\]
+ VGND VGND VPWR VPWR _11802_ sky130_fd_sc_hd__xnor2_1
X_29414_ clknet_leaf_328_clk _03212_ net136 VGND VGND VPWR VPWR C_out\[386\] sky130_fd_sc_hd__dfrtp_1
X_23838_ _10431_ _10432_ _10430_ VGND VGND VPWR VPWR _10433_ sky130_fd_sc_hd__o21ai_1
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29345_ clknet_leaf_224_clk _03143_ net147 VGND VGND VPWR VPWR C_out\[317\] sky130_fd_sc_hd__dfrtp_1
X_14571_ _11739_ _11740_ _11741_ VGND VGND VPWR VPWR _11743_ sky130_fd_sc_hd__and3_1
XFILLER_72_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26557_ clknet_leaf_2_A_in_serial_clk _00360_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_199_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23769_ _10357_ _10373_ VGND VGND VPWR VPWR _10374_ sky130_fd_sc_hd__nor2_1
XFILLER_198_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_clk clknet_5_19__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16310_ systolic_inst.A_outs\[12\]\[6\] _11260_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_101_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25508_ _00008_ _11233_ VGND VGND VPWR VPWR _11235_ sky130_fd_sc_hd__nor2_1
XFILLER_198_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13522_ deser_A.shift_reg\[86\] deser_A.shift_reg\[87\] net129 VGND VGND VPWR VPWR
+ _00359_ sky130_fd_sc_hd__mux2_1
XFILLER_242_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29276_ clknet_leaf_188_clk _03074_ net146 VGND VGND VPWR VPWR C_out\[248\] sky130_fd_sc_hd__dfrtp_1
X_17290_ _04546_ _04547_ _04519_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a21oi_1
X_26488_ clknet_leaf_8_A_in_serial_clk _00291_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28227_ clknet_leaf_124_clk _02025_ VGND VGND VPWR VPWR systolic_inst.B_shift\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16241_ _03548_ _03552_ _03583_ _03584_ _03621_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__a311o_2
X_25439_ _11279_ _11188_ _11189_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__and3_1
X_13453_ deser_A.shift_reg\[17\] deser_A.shift_reg\[18\] deser_A.receiving VGND VGND
+ VPWR VPWR _00290_ sky130_fd_sc_hd__mux2_1
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28158_ clknet_leaf_106_clk _01956_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16172_ _03523_ _03525_ _03522_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__o21ba_1
XFILLER_51_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13384_ A_in\[93\] deser_A.word_buffer\[93\] net95 VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27109_ clknet_leaf_26_B_in_serial_clk _00907_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_15123_ _12211_ _12214_ _12237_ VGND VGND VPWR VPWR _12239_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28089_ clknet_leaf_116_clk _01887_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_177_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19931_ systolic_inst.B_outs\[6\]\[5\] systolic_inst.A_outs\[6\]\[7\] VGND VGND VPWR
+ VPWR _06928_ sky130_fd_sc_hd__nand2_1
X_15054_ net118 _12170_ _12171_ _12172_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_71_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14005_ deser_B.shift_reg\[39\] deser_B.shift_reg\[40\] deser_B.receiving VGND VGND
+ VPWR VPWR _00831_ sky130_fd_sc_hd__mux2_1
XFILLER_141_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_220_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19862_ systolic_inst.B_outs\[6\]\[5\] systolic_inst.A_outs\[6\]\[5\] VGND VGND VPWR
+ VPWR _06861_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_220_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_220_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18813_ _05922_ _05925_ _05929_ _05930_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__o211a_1
X_19793_ systolic_inst.A_outs\[6\]\[1\] systolic_inst.A_outs\[6\]\[2\] systolic_inst.B_outs\[6\]\[6\]
+ systolic_inst.B_outs\[6\]\[7\] VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__and4b_1
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18744_ _05866_ _05867_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__nor2_1
X_15956_ _12969_ _12973_ _12974_ VGND VGND VPWR VPWR _12975_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14907_ _12001_ _12003_ _12002_ VGND VGND VPWR VPWR _12029_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_69_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15887_ systolic_inst.acc_wires\[13\]\[16\] systolic_inst.acc_wires\[13\]\[17\] systolic_inst.acc_wires\[13\]\[18\]
+ systolic_inst.acc_wires\[13\]\[19\] systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12917_ sky130_fd_sc_hd__o41a_1
X_18675_ _05695_ _05800_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__or2_1
XFILLER_184_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17626_ _04863_ _04864_ _04862_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_218_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14838_ systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[5\] systolic_inst.A_outs\[14\]\[6\]
+ systolic_inst.B_outs\[14\]\[0\] VGND VGND VPWR VPWR _11962_ sky130_fd_sc_hd__a22oi_1
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14769_ _11895_ _11896_ VGND VGND VPWR VPWR _11897_ sky130_fd_sc_hd__nand2_1
X_17557_ _04805_ _04806_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_28_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_177_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16508_ _03860_ _03863_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__or3_1
XFILLER_225_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17488_ _04739_ _04740_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__nand2_1
XFILLER_177_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19227_ _06254_ _06256_ _06290_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16439_ _03801_ _03802_ _03803_ net61 VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__a31o_1
XFILLER_34_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19158_ _06207_ _06223_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18109_ _05263_ _05265_ _05264_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__o21ba_1
XFILLER_69_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19089_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[5\] _06154_ _06155_
+ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__o2bb2a_1
X_21120_ _07989_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__inv_2
XFILLER_236_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21051_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.A_outs\[4\]\[7\] VGND VGND VPWR
+ VPWR _07923_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_58_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20002_ _06949_ _06972_ _06973_ _06996_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__o211ai_2
XFILLER_115_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24810_ net113 ser_C.shift_reg\[233\] VGND VGND VPWR VPWR _10875_ sky130_fd_sc_hd__and2_1
XFILLER_80_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25790_ systolic_inst.acc_wires\[8\]\[10\] C_out\[266\] net22 VGND VGND VPWR VPWR
+ _03092_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_203_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24741_ C_out\[197\] net97 net77 ser_C.shift_reg\[197\] _10840_ VGND VGND VPWR VPWR
+ _02447_ sky130_fd_sc_hd__a221o_1
XFILLER_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21953_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[3\]\[13\]
+ VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__or2_1
XFILLER_82_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_195_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27460_ clknet_leaf_238_clk _01258_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_20904_ systolic_inst.A_outs\[4\]\[0\] systolic_inst.B_outs\[4\]\[1\] systolic_inst.A_outs\[4\]\[4\]
+ systolic_inst.B_outs\[4\]\[5\] VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_195_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24672_ net110 ser_C.shift_reg\[164\] VGND VGND VPWR VPWR _10806_ sky130_fd_sc_hd__and2_1
XFILLER_242_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21884_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[3\]\[3\]
+ VGND VGND VPWR VPWR _08682_ sky130_fd_sc_hd__and2_1
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26411_ clknet_leaf_5_clk _00218_ net131 VGND VGND VPWR VPWR A_in\[79\] sky130_fd_sc_hd__dfrtp_1
X_23623_ _10205_ _10208_ _10243_ VGND VGND VPWR VPWR _10244_ sky130_fd_sc_hd__o21ai_2
XFILLER_36_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20835_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_shift\[3\]\[0\] net120 VGND
+ VGND VPWR VPWR _01658_ sky130_fd_sc_hd__mux2_1
X_27391_ clknet_leaf_337_clk _01189_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_clk clknet_5_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
X_29130_ clknet_leaf_172_clk _02928_ net148 VGND VGND VPWR VPWR C_out\[102\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26342_ clknet_leaf_60_clk _00149_ net144 VGND VGND VPWR VPWR A_in\[10\] sky130_fd_sc_hd__dfrtp_1
X_23554_ _10172_ _10174_ _10109_ _10111_ VGND VGND VPWR VPWR _10177_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_154_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20766_ _07671_ _07672_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_154_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29061_ clknet_leaf_108_clk _02859_ net150 VGND VGND VPWR VPWR C_out\[33\] sky130_fd_sc_hd__dfrtp_1
X_22505_ net65 _09234_ _09236_ systolic_inst.acc_wires\[2\]\[5\] net109 VGND VGND
+ VPWR VPWR _01815_ sky130_fd_sc_hd__a32o_1
XFILLER_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26273_ clknet_leaf_21_A_in_serial_clk _00081_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23485_ _10105_ _10106_ _10107_ VGND VGND VPWR VPWR _10109_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_150_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20697_ _07597_ _07613_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__nor2_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28012_ clknet_leaf_152_clk _01810_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_206_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25224_ net110 ser_C.shift_reg\[440\] VGND VGND VPWR VPWR _11082_ sky130_fd_sc_hd__and2_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22436_ _09174_ _09175_ VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__and2b_1
XFILLER_149_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25155_ C_out\[404\] net101 net73 ser_C.shift_reg\[404\] _11047_ VGND VGND VPWR VPWR
+ _02654_ sky130_fd_sc_hd__a221o_1
X_22367_ _09107_ _09108_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__nand2_1
X_24106_ systolic_inst.B_shift\[1\]\[1\] _11332_ net83 systolic_inst.B_shift\[5\]\[1\]
+ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__a22o_1
XFILLER_151_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21318_ _08165_ _08169_ _08172_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__nand3_1
XFILLER_174_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25086_ net113 ser_C.shift_reg\[371\] VGND VGND VPWR VPWR _11013_ sky130_fd_sc_hd__and2_1
X_22298_ _09024_ _09041_ VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__xor2_1
XFILLER_105_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24037_ systolic_inst.B_shift\[8\]\[6\] B_in\[38\] _00008_ VGND VGND VPWR VPWR _10536_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28914_ clknet_leaf_282_clk _02712_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_148_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21249_ _08113_ _08114_ net117 VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__o21ai_1
XFILLER_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28845_ clknet_leaf_334_clk _02643_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[393\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15810_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[13\]\[8\]
+ _12847_ VGND VGND VPWR VPWR _12851_ sky130_fd_sc_hd__and3_1
X_16790_ _04101_ _04109_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__nand2_1
X_25988_ systolic_inst.acc_wires\[14\]\[16\] ser_C.parallel_data\[464\] net25 VGND
+ VGND VPWR VPWR _03290_ sky130_fd_sc_hd__mux2_1
X_28776_ clknet_leaf_229_clk _02574_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[324\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_237_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15741_ _12789_ _12791_ VGND VGND VPWR VPWR _12793_ sky130_fd_sc_hd__xor2_1
X_27727_ clknet_leaf_215_clk _01525_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_24939_ C_out\[296\] net102 net76 ser_C.shift_reg\[296\] _10939_ VGND VGND VPWR VPWR
+ _02546_ sky130_fd_sc_hd__a221o_1
XFILLER_219_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _12687_ _12725_ VGND VGND VPWR VPWR _12726_ sky130_fd_sc_hd__xnor2_1
X_18460_ _05589_ _05590_ _05572_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_103_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27658_ clknet_leaf_302_clk _01456_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[15\]\[14\]
+ VGND VGND VPWR VPWR _11787_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _04632_ _04635_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__nor2_1
X_26609_ clknet_leaf_15_B_in_serial_clk _00412_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_18391_ systolic_inst.acc_wires\[9\]\[28\] systolic_inst.acc_wires\[9\]\[29\] systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_64_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27589_ clknet_leaf_223_clk _01387_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_25_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_14_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_950 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17342_ systolic_inst.B_outs\[10\]\[7\] _04564_ _04565_ VGND VGND VPWR VPWR _04599_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_18_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14554_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[15\]\[4\]
+ VGND VGND VPWR VPWR _11728_ sky130_fd_sc_hd__or2_1
X_29328_ clknet_leaf_221_clk _03126_ net139 VGND VGND VPWR VPWR C_out\[300\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13505_ deser_A.shift_reg\[69\] deser_A.shift_reg\[70\] net129 VGND VGND VPWR VPWR
+ _00342_ sky130_fd_sc_hd__mux2_1
XFILLER_159_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17273_ systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[5\] systolic_inst.A_outs\[10\]\[6\]
+ systolic_inst.B_outs\[10\]\[0\] VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__a22oi_1
X_29259_ clknet_leaf_196_clk _03057_ net146 VGND VGND VPWR VPWR C_out\[231\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _11622_ _11634_ _11632_ VGND VGND VPWR VPWR _11666_ sky130_fd_sc_hd__o21a_1
XFILLER_202_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19012_ systolic_inst.A_outs\[7\]\[1\] systolic_inst.A_outs\[6\]\[1\] net119 VGND
+ VGND VPWR VPWR _01459_ sky130_fd_sc_hd__mux2_1
X_16224_ _03605_ _03606_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13436_ _00002_ _11310_ _11318_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__and3b_1
Xclkload206 clknet_leaf_36_clk VGND VGND VPWR VPWR clkload206/Y sky130_fd_sc_hd__inv_6
XFILLER_173_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload217 clknet_leaf_49_clk VGND VGND VPWR VPWR clkload217/Y sky130_fd_sc_hd__clkinv_8
Xclkload228 clknet_leaf_72_clk VGND VGND VPWR VPWR clkload228/X sky130_fd_sc_hd__clkbuf_8
Xclkload239 clknet_leaf_89_clk VGND VGND VPWR VPWR clkload239/X sky130_fd_sc_hd__clkbuf_4
X_16155_ _03521_ _03538_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__xor2_1
X_13367_ A_in\[76\] deser_A.word_buffer\[76\] net96 VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__mux2_1
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15106_ _12220_ _12221_ VGND VGND VPWR VPWR _12223_ sky130_fd_sc_hd__and2b_1
XFILLER_127_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16086_ _13054_ _13079_ _13080_ VGND VGND VPWR VPWR _13082_ sky130_fd_sc_hd__nor3_1
X_13298_ A_in\[7\] deser_A.word_buffer\[7\] net93 VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__mux2_1
X_19914_ _06909_ _06910_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__xnor2_1
X_15037_ _12146_ _12154_ VGND VGND VPWR VPWR _12156_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19845_ _06842_ _06843_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19776_ net106 systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[7\] VGND
+ VGND VPWR VPWR _06778_ sky130_fd_sc_hd__nand2_1
X_16988_ _04291_ _04292_ _04290_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18727_ _05801_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__and2b_1
XFILLER_110_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15939_ _12959_ _12960_ VGND VGND VPWR VPWR _12961_ sky130_fd_sc_hd__nand2_1
XFILLER_97_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18658_ _05766_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__xor2_1
Xwire47 net49 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_8
XFILLER_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire58 _00002_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_12
X_17609_ _04850_ _04851_ _04852_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__a21o_1
XFILLER_91_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18589_ _05664_ _05679_ _05678_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__o21a_1
XFILLER_33_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_190_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20620_ net116 systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[5\]\[0\]
+ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_211_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20551_ _07430_ _07482_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__nor2_1
XFILLER_193_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23270_ _09909_ _09912_ VGND VGND VPWR VPWR _09913_ sky130_fd_sc_hd__nand2_1
XFILLER_158_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20482_ _07416_ _07415_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__nand2b_1
XFILLER_20_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22221_ _08959_ _08965_ VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22152_ systolic_inst.A_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\]
+ systolic_inst.A_outs\[2\]\[1\] VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__a22o_1
XFILLER_173_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21103_ _07971_ _07972_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__xor2_1
XFILLER_156_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22083_ systolic_inst.A_outs\[2\]\[5\] systolic_inst.A_outs\[1\]\[5\] net122 VGND
+ VGND VPWR VPWR _01783_ sky130_fd_sc_hd__mux2_1
XFILLER_160_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26960_ clknet_leaf_27_A_in_serial_clk _00758_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_236_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_205_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25911_ systolic_inst.acc_wires\[12\]\[3\] C_out\[387\] net21 VGND VGND VPWR VPWR
+ _03213_ sky130_fd_sc_hd__mux2_1
X_21034_ _07864_ _07866_ _07906_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__a21oi_2
X_26891_ clknet_leaf_8_A_in_serial_clk _00689_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28630_ clknet_leaf_204_clk _02428_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_143_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25842_ systolic_inst.acc_wires\[9\]\[30\] C_out\[318\] net13 VGND VGND VPWR VPWR
+ _03144_ sky130_fd_sc_hd__mux2_1
XFILLER_75_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28561_ clknet_leaf_167_clk _02359_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_170_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25773_ systolic_inst.acc_wires\[7\]\[25\] C_out\[249\] net44 VGND VGND VPWR VPWR
+ _03075_ sky130_fd_sc_hd__mux2_1
X_22985_ _09659_ _09660_ VGND VGND VPWR VPWR _09662_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24724_ net113 ser_C.shift_reg\[190\] VGND VGND VPWR VPWR _10832_ sky130_fd_sc_hd__and2_1
XFILLER_28_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27512_ clknet_leaf_231_clk _01310_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_28492_ clknet_leaf_116_clk _02290_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_21936_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[3\]\[11\]
+ VGND VGND VPWR VPWR _08726_ sky130_fd_sc_hd__nand2_1
XFILLER_227_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_216_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27443_ clknet_leaf_242_clk _01241_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24655_ C_out\[154\] net104 _10643_ ser_C.shift_reg\[154\] _10797_ VGND VGND VPWR
+ VPWR _02404_ sky130_fd_sc_hd__a221o_1
XFILLER_70_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21867_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[3\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__a21o_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23606_ _10186_ _10225_ VGND VGND VPWR VPWR _10227_ sky130_fd_sc_hd__nand2_1
XFILLER_230_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20818_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[30\]
+ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_152_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27374_ clknet_leaf_327_clk _01172_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24586_ net114 ser_C.shift_reg\[121\] VGND VGND VPWR VPWR _10763_ sky130_fd_sc_hd__and2_1
XFILLER_169_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21798_ _08600_ _08601_ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29113_ clknet_leaf_157_clk _02911_ net150 VGND VGND VPWR VPWR C_out\[85\] sky130_fd_sc_hd__dfrtp_1
XFILLER_208_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26325_ clknet_leaf_30_A_in_serial_clk _00133_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_169_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23537_ _10120_ _10159_ VGND VGND VPWR VPWR _10160_ sky130_fd_sc_hd__xnor2_1
X_20749_ net106 systolic_inst.acc_wires\[5\]\[19\] net68 _07658_ VGND VGND VPWR VPWR
+ _01637_ sky130_fd_sc_hd__a22o_1
XFILLER_211_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29044_ clknet_leaf_100_clk _02842_ net152 VGND VGND VPWR VPWR C_out\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14270_ _11417_ _11456_ VGND VGND VPWR VPWR _11457_ sky130_fd_sc_hd__nand2_1
X_26256_ clknet_leaf_3_A_in_serial_clk _00064_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_23468_ _10089_ _10090_ _10072_ VGND VGND VPWR VPWR _10093_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25207_ C_out\[430\] net101 net73 ser_C.shift_reg\[430\] _11073_ VGND VGND VPWR VPWR
+ _02680_ sky130_fd_sc_hd__a221o_1
X_13221_ deser_A.word_buffer\[59\] deser_A.serial_word\[59\] net128 VGND VGND VPWR
+ VPWR _00069_ sky130_fd_sc_hd__mux2_1
XFILLER_109_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22419_ _09128_ _09131_ _09158_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__o21ai_1
X_26187_ _11252_ _11253_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__nor2_1
X_23399_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.A_outs\[0\]\[7\] VGND VGND VPWR
+ VPWR _10025_ sky130_fd_sc_hd__and2_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13152_ _11301_ _11303_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__nand2_1
XFILLER_178_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25138_ net110 ser_C.shift_reg\[397\] VGND VGND VPWR VPWR _11039_ sky130_fd_sc_hd__and2_1
XFILLER_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25069_ C_out\[361\] net97 net77 ser_C.shift_reg\[361\] _11004_ VGND VGND VPWR VPWR
+ _02611_ sky130_fd_sc_hd__a221o_1
X_17960_ _05148_ _05151_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__xnor2_1
XFILLER_215_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_219_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16911_ systolic_inst.B_outs\[11\]\[6\] systolic_inst.A_outs\[11\]\[7\] VGND VGND
+ VPWR VPWR _04227_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_109_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17891_ _05084_ _05085_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__or2_1
X_19630_ systolic_inst.B_outs\[6\]\[0\] systolic_inst.A_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[1\]
+ systolic_inst.A_outs\[6\]\[1\] VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__and4_1
XFILLER_215_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28828_ clknet_leaf_195_clk _02626_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[376\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16842_ _04158_ _04159_ _04157_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_6_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19561_ net62 _06593_ _06594_ systolic_inst.acc_wires\[7\]\[23\] net105 VGND VGND
+ VPWR VPWR _01513_ sky130_fd_sc_hd__a32o_1
XFILLER_150_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13985_ deser_B.shift_reg\[19\] deser_B.shift_reg\[20\] net125 VGND VGND VPWR VPWR
+ _00811_ sky130_fd_sc_hd__mux2_1
X_28759_ clknet_leaf_218_clk _02557_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[307\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16773_ _04063_ _04065_ _04062_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__o21ba_1
XFILLER_168_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_3__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_5_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_18512_ _05612_ _05641_ _05642_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_215_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ _12687_ _12774_ VGND VGND VPWR VPWR _12776_ sky130_fd_sc_hd__and2_1
XFILLER_46_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ _06530_ _06534_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__nand2_1
XFILLER_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_222_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18443_ _05570_ _05575_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_17_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15655_ _12672_ _12678_ _12709_ VGND VGND VPWR VPWR _12710_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_17_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14606_ _11762_ _11767_ _11768_ VGND VGND VPWR VPWR _11772_ sky130_fd_sc_hd__nand3_1
X_18374_ _05525_ _05529_ _05526_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_1_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15586_ net107 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[9\] _12641_
+ _12642_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__a22o_1
XFILLER_222_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14537_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[15\]\[0\]
+ _11708_ _11709_ VGND VGND VPWR VPWR _11714_ sky130_fd_sc_hd__a22o_1
X_17325_ _04576_ _04582_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__nor2_1
XFILLER_239_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14468_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[12\] _11649_ net118
+ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__mux2_1
X_17256_ _04513_ _04514_ _04515_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_42_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16207_ _03517_ _03589_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__nor2_1
X_13419_ net1 net130 deser_A.bit_idx\[0\] VGND VGND VPWR VPWR _11308_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_96_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17187_ systolic_inst.B_outs\[9\]\[1\] systolic_inst.B_outs\[5\]\[1\] net116 VGND
+ VGND VPWR VPWR _01275_ sky130_fd_sc_hd__mux2_1
X_14399_ _11580_ _11581_ _11582_ VGND VGND VPWR VPWR _11583_ sky130_fd_sc_hd__o21a_1
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16138_ systolic_inst.B_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[5\]
+ systolic_inst.B_outs\[12\]\[3\] VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__a22oi_1
XPHY_EDGE_ROW_216_Right_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16069_ systolic_inst.B_outs\[12\]\[3\] systolic_inst.A_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\]
+ systolic_inst.A_outs\[12\]\[2\] VGND VGND VPWR VPWR _13065_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_55_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_29_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_B_in_serial_clk B_in_serial_clk VGND VGND VPWR VPWR clknet_0_B_in_serial_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_51_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19828_ _06826_ _06827_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19759_ _06757_ _06760_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_192_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22770_ _09452_ _09449_ VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__nand2b_1
XFILLER_83_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21721_ _08527_ _08526_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_49_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24440_ net114 ser_C.shift_reg\[48\] VGND VGND VPWR VPWR _10690_ sky130_fd_sc_hd__and2_1
X_21652_ _08452_ _08460_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__nand2_1
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20603_ _07531_ _07532_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__and2b_1
X_24371_ C_out\[12\] net104 _10643_ ser_C.shift_reg\[12\] _10655_ VGND VGND VPWR VPWR
+ _02262_ sky130_fd_sc_hd__a221o_1
XFILLER_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21583_ _08363_ _08393_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26110_ deser_B.serial_word\[65\] deser_B.shift_reg\[65\] _00001_ VGND VGND VPWR
+ VPWR _03412_ sky130_fd_sc_hd__mux2_1
XFILLER_178_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23322_ _09948_ _09949_ _09931_ VGND VGND VPWR VPWR _09951_ sky130_fd_sc_hd__a21bo_1
X_27090_ clknet_leaf_5_B_in_serial_clk _00888_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_20534_ systolic_inst.A_outs\[5\]\[5\] systolic_inst.B_outs\[5\]\[6\] systolic_inst.A_outs\[5\]\[6\]
+ systolic_inst.B_outs\[5\]\[7\] VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__and4b_1
XFILLER_137_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26041_ systolic_inst.B_outs\[15\]\[5\] systolic_inst.B_outs\[11\]\[5\] net118 VGND
+ VGND VPWR VPWR _03343_ sky130_fd_sc_hd__mux2_1
X_23253_ systolic_inst.acc_wires\[1\]\[26\] systolic_inst.acc_wires\[1\]\[27\] systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09898_ sky130_fd_sc_hd__o21a_1
XFILLER_181_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20465_ _07364_ _07399_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__xor2_1
XFILLER_10_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22204_ _08948_ _08949_ VGND VGND VPWR VPWR _08950_ sky130_fd_sc_hd__nand2_1
X_23184_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[1\]\[17\]
+ VGND VGND VPWR VPWR _09840_ sky130_fd_sc_hd__xor2_2
XFILLER_180_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20396_ systolic_inst.A_outs\[5\]\[1\] systolic_inst.B_outs\[5\]\[7\] VGND VGND VPWR
+ VPWR _07333_ sky130_fd_sc_hd__and2b_1
XFILLER_84_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22135_ _08876_ _08882_ _08883_ VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_145_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27992_ clknet_leaf_122_clk _01790_ net153 VGND VGND VPWR VPWR systolic_inst.B_outs\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_145_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22066_ _08829_ _08832_ _08836_ VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__or3_1
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26943_ clknet_leaf_20_A_in_serial_clk _00741_ net131 VGND VGND VPWR VPWR deser_A.serial_word\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21017_ systolic_inst.A_outs\[4\]\[1\] _07852_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__nor2_1
XFILLER_212_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29662_ clknet_leaf_10_B_in_serial_clk _03457_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26874_ clknet_leaf_14_A_in_serial_clk _00672_ net143 VGND VGND VPWR VPWR deser_A.serial_word\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_28613_ clknet_leaf_40_clk _02411_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[161\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25825_ systolic_inst.acc_wires\[9\]\[13\] C_out\[301\] net15 VGND VGND VPWR VPWR
+ _03127_ sky130_fd_sc_hd__mux2_1
X_29593_ clknet_leaf_13_B_in_serial_clk _03388_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28544_ clknet_leaf_164_clk _02342_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13770_ B_in\[77\] deser_B.word_buffer\[77\] net88 VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__mux2_1
X_25756_ systolic_inst.acc_wires\[7\]\[8\] C_out\[232\] net42 VGND VGND VPWR VPWR
+ _03058_ sky130_fd_sc_hd__mux2_1
X_22968_ _09586_ _09645_ VGND VGND VPWR VPWR _09646_ sky130_fd_sc_hd__xnor2_1
XFILLER_210_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21919_ _08706_ _08709_ _08710_ net60 VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__a31o_1
X_24707_ C_out\[180\] net99 net79 ser_C.shift_reg\[180\] _10823_ VGND VGND VPWR VPWR
+ _02430_ sky130_fd_sc_hd__a221o_1
XFILLER_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28475_ clknet_leaf_106_clk _02273_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25687_ systolic_inst.acc_wires\[5\]\[3\] C_out\[163\] net16 VGND VGND VPWR VPWR
+ _02989_ sky130_fd_sc_hd__mux2_1
X_22899_ _09552_ _09578_ VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__xnor2_1
XFILLER_231_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15440_ _12482_ _12500_ VGND VGND VPWR VPWR _12501_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_175_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24638_ net7 ser_C.shift_reg\[147\] VGND VGND VPWR VPWR _10789_ sky130_fd_sc_hd__and2_1
XFILLER_128_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27426_ clknet_leaf_249_clk _01224_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_230_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15371_ systolic_inst.B_outs\[12\]\[7\] systolic_inst.B_outs\[8\]\[7\] net115 VGND
+ VGND VPWR VPWR _01089_ sky130_fd_sc_hd__mux2_1
XFILLER_230_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24569_ C_out\[111\] net100 net80 ser_C.shift_reg\[111\] _10754_ VGND VGND VPWR VPWR
+ _02361_ sky130_fd_sc_hd__a221o_1
X_27357_ clknet_leaf_323_clk _01155_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17110_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[21\]
+ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__xnor2_2
X_14322_ _11506_ _11507_ VGND VGND VPWR VPWR _11508_ sky130_fd_sc_hd__or2_1
XFILLER_141_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26308_ clknet_leaf_24_A_in_serial_clk _00116_ net134 VGND VGND VPWR VPWR deser_A.word_buffer\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_18090_ _05278_ _05279_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nor2_1
XFILLER_184_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27288_ clknet_leaf_319_clk _01086_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_134_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17041_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[11\]\[11\]
+ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__nand2_1
XFILLER_239_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29027_ clknet_leaf_92_clk _02825_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14253_ _11439_ VGND VGND VPWR VPWR _11440_ sky130_fd_sc_hd__inv_2
X_26239_ clknet_leaf_16_A_in_serial_clk _00047_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_171_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13204_ deser_A.word_buffer\[42\] deser_A.serial_word\[42\] net127 VGND VGND VPWR
+ VPWR _00052_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14184_ _11371_ _11372_ VGND VGND VPWR VPWR _11374_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_91_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13135_ systolic_inst.cycle_cnt\[19\] systolic_inst.cycle_cnt\[18\] systolic_inst.cycle_cnt\[17\]
+ systolic_inst.cycle_cnt\[16\] VGND VGND VPWR VPWR _11288_ sky130_fd_sc_hd__or4_1
XFILLER_140_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18992_ _06081_ _06084_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__xor2_1
XFILLER_98_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17943_ _05136_ _05135_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__nand2b_1
XFILLER_215_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17874_ _05067_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19613_ systolic_inst.A_outs\[6\]\[1\] systolic_inst.A_outs\[5\]\[1\] net120 VGND
+ VGND VPWR VPWR _01523_ sky130_fd_sc_hd__mux2_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16825_ _04134_ _04142_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_89_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19544_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[21\]
+ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__xnor2_2
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16756_ _04076_ _04075_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__and2b_1
X_13968_ deser_B.shift_reg\[2\] deser_B.shift_reg\[3\] net125 VGND VGND VPWR VPWR
+ _00794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15707_ _12716_ _12759_ VGND VGND VPWR VPWR _12760_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19475_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[7\]\[11\]
+ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__nand2_1
XFILLER_207_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16687_ _04007_ _04008_ _03978_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__a21o_1
X_13899_ deser_A.serial_word\[60\] deser_A.shift_reg\[60\] _00002_ VGND VGND VPWR
+ VPWR _00725_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_234_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_234_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18426_ systolic_inst.B_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[1\] systolic_inst.A_outs\[8\]\[2\]
+ systolic_inst.B_outs\[8\]\[0\] VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__a22oi_1
XFILLER_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15638_ _12651_ _12653_ _12652_ VGND VGND VPWR VPWR _12693_ sky130_fd_sc_hd__o21ba_1
XFILLER_107_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18357_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[24\]
+ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__and2_1
XFILLER_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15569_ systolic_inst.A_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[5\] _12589_ _12588_
+ VGND VGND VPWR VPWR _12626_ sky130_fd_sc_hd__a31oi_1
XFILLER_222_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17308_ systolic_inst.B_outs\[10\]\[7\] _04564_ _04565_ VGND VGND VPWR VPWR _04566_
+ sky130_fd_sc_hd__and3_1
XFILLER_174_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18288_ _05447_ _05452_ _05451_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__o21a_1
XFILLER_119_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17239_ _04498_ _04499_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__nand2_1
XFILLER_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20250_ _07185_ _07191_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_181_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20181_ _07148_ _07149_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__nor2_1
XFILLER_170_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23940_ systolic_inst.B_shift\[14\]\[2\] B_in\[18\] net59 VGND VGND VPWR VPWR _10499_
+ sky130_fd_sc_hd__mux2_1
XFILLER_233_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23871_ _10453_ _10457_ VGND VGND VPWR VPWR _10460_ sky130_fd_sc_hd__nor2_1
XFILLER_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25610_ systolic_inst.acc_wires\[2\]\[22\] C_out\[86\] net52 VGND VGND VPWR VPWR
+ _02912_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22822_ _09500_ _09501_ _09502_ VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_179_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26590_ clknet_leaf_30_A_in_serial_clk _00393_ net132 VGND VGND VPWR VPWR deser_A.shift_reg\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_64_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25541_ systolic_inst.acc_wires\[0\]\[17\] C_out\[17\] net54 VGND VGND VPWR VPWR
+ _02843_ sky130_fd_sc_hd__mux2_1
XFILLER_25_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22753_ _09435_ _09436_ VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__or2_1
XFILLER_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21704_ _08473_ _08477_ _08510_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__o21ai_1
X_28260_ clknet_leaf_57_clk _02058_ VGND VGND VPWR VPWR systolic_inst.B_shift\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25472_ _00008_ _11211_ VGND VGND VPWR VPWR _11212_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22684_ systolic_inst.B_outs\[0\]\[3\] systolic_inst.B_shift\[0\]\[3\] net121 VGND
+ VGND VPWR VPWR _01853_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24423_ C_out\[38\] _11302_ net81 ser_C.shift_reg\[38\] _10681_ VGND VGND VPWR VPWR
+ _02288_ sky130_fd_sc_hd__a221o_1
XFILLER_200_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27211_ clknet_leaf_247_clk _01009_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_21635_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] _08443_ VGND
+ VGND VPWR VPWR _08444_ sky130_fd_sc_hd__a21o_1
X_28191_ clknet_leaf_129_clk _01989_ VGND VGND VPWR VPWR systolic_inst.B_shift\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27142_ clknet_leaf_13_clk _00940_ VGND VGND VPWR VPWR systolic_inst.A_shift\[21\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24354_ net7 ser_C.shift_reg\[5\] VGND VGND VPWR VPWR _10647_ sky130_fd_sc_hd__and2_1
X_21566_ _08373_ _08376_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__xor2_1
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23305_ _09929_ _09934_ VGND VGND VPWR VPWR _09935_ sky130_fd_sc_hd__xnor2_1
X_27073_ clknet_leaf_10_B_in_serial_clk _00871_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_20517_ _07450_ _07449_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__and2b_1
X_24285_ systolic_inst.B_shift\[27\]\[6\] B_in\[94\] _00008_ VGND VGND VPWR VPWR _10616_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21497_ systolic_inst.A_outs\[3\]\[0\] systolic_inst.A_outs\[3\]\[1\] systolic_inst.B_outs\[3\]\[2\]
+ systolic_inst.B_outs\[3\]\[3\] VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__and4_1
XFILLER_193_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26024_ systolic_inst.acc_wires\[15\]\[20\] ser_C.parallel_data\[500\] net23 VGND
+ VGND VPWR VPWR _03326_ sky130_fd_sc_hd__mux2_1
X_23236_ _09884_ _09883_ systolic_inst.acc_wires\[1\]\[24\] net109 VGND VGND VPWR
+ VPWR _01898_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20448_ _07383_ _07382_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__nand2b_1
XFILLER_180_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23167_ _09822_ _09825_ VGND VGND VPWR VPWR _09826_ sky130_fd_sc_hd__nand2_1
XFILLER_106_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20379_ _07250_ _07251_ _07282_ _07281_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22118_ _08861_ _08866_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23098_ net64 _09764_ _09766_ systolic_inst.acc_wires\[1\]\[4\] _11258_ VGND VGND
+ VPWR VPWR _01878_ sky130_fd_sc_hd__a32o_1
X_27975_ clknet_leaf_172_clk _01773_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22049_ _08815_ _08819_ _08821_ net60 VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__a31o_1
X_14940_ _12061_ VGND VGND VPWR VPWR _12062_ sky130_fd_sc_hd__inv_2
X_26926_ clknet_leaf_5_A_in_serial_clk _00724_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29645_ clknet_leaf_32_B_in_serial_clk _03440_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_236_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26857_ clknet_leaf_0_B_in_serial_clk _00659_ net134 VGND VGND VPWR VPWR deser_B.bit_idx\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14871_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[6\]
+ systolic_inst.A_outs\[14\]\[7\] VGND VGND VPWR VPWR _11994_ sky130_fd_sc_hd__nand4_1
XFILLER_76_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16610_ systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[2\] systolic_inst.A_outs\[11\]\[3\]
+ systolic_inst.B_outs\[11\]\[0\] VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__a22o_1
XFILLER_217_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13822_ net126 deser_B.bit_idx\[0\] _11319_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_123_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25808_ systolic_inst.acc_wires\[8\]\[28\] C_out\[284\] net27 VGND VGND VPWR VPWR
+ _03110_ sky130_fd_sc_hd__mux2_1
X_29576_ clknet_leaf_22_B_in_serial_clk _03371_ net137 VGND VGND VPWR VPWR deser_B.serial_word\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17590_ _04836_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__inv_2
X_26788_ clknet_leaf_69_clk _00590_ net135 VGND VGND VPWR VPWR B_in\[60\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28527_ clknet_leaf_166_clk _02325_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_204_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13753_ B_in\[60\] deser_B.word_buffer\[60\] net89 VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__mux2_1
XFILLER_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16541_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[26\]
+ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__nand2_1
X_25739_ systolic_inst.acc_wires\[6\]\[23\] C_out\[215\] net46 VGND VGND VPWR VPWR
+ _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_189_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19260_ _06321_ _06322_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__nand2_1
XFILLER_56_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28458_ clknet_leaf_123_clk _02256_ net144 VGND VGND VPWR VPWR ser_C.shift_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13684_ deser_B.word_buffer\[120\] deser_B.serial_word\[120\] deser_B.serial_word_ready
+ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__mux2_1
X_16472_ _03833_ _03832_ systolic_inst.acc_wires\[12\]\[15\] net108 VGND VGND VPWR
+ VPWR _01185_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18211_ _05391_ _05392_ _05384_ _05388_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__a211o_1
X_15423_ systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[4\] systolic_inst.A_outs\[13\]\[5\]
+ systolic_inst.B_outs\[13\]\[0\] VGND VGND VPWR VPWR _12484_ sky130_fd_sc_hd__a22oi_1
X_27409_ clknet_leaf_226_clk _01207_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_19191_ _06247_ _06255_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__nand2_1
XFILLER_54_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28389_ clknet_leaf_34_clk _02187_ VGND VGND VPWR VPWR systolic_inst.A_shift\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15354_ _12430_ _12434_ _12435_ net61 VGND VGND VPWR VPWR _12437_ sky130_fd_sc_hd__a31o_1
X_18142_ _05262_ _05328_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__or2_1
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14305_ _11488_ _11489_ VGND VGND VPWR VPWR _11491_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_93_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15285_ _12377_ _12378_ _12375_ VGND VGND VPWR VPWR _12379_ sky130_fd_sc_hd__o21ai_2
X_18073_ systolic_inst.B_outs\[9\]\[5\] systolic_inst.A_outs\[9\]\[6\] VGND VGND VPWR
+ VPWR _05263_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_242_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14236_ _11421_ _11422_ _11410_ VGND VGND VPWR VPWR _11424_ sky130_fd_sc_hd__o21bai_1
X_17024_ _04328_ _04327_ systolic_inst.acc_wires\[11\]\[8\] net105 VGND VGND VPWR
+ VPWR _01242_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_242_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14167_ net107 systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[3\] VGND
+ VGND VPWR VPWR _11358_ sky130_fd_sc_hd__and2_1
XFILLER_140_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13118_ systolic_inst.B_outs\[3\]\[7\] VGND VGND VPWR VPWR _11274_ sky130_fd_sc_hd__inv_2
X_14098_ net151 _11306_ VGND VGND VPWR VPWR _11332_ sky130_fd_sc_hd__nand2_8
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18975_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[26\]
+ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_223_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xload_slew145 net147 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_16
X_17926_ systolic_inst.B_outs\[9\]\[3\] systolic_inst.A_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\]
+ systolic_inst.A_outs\[9\]\[4\] VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__and4_1
XFILLER_230_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17857_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[4\]
+ systolic_inst.A_outs\[9\]\[5\] VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__and4_1
XFILLER_239_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_236_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16808_ _04097_ _04098_ _04099_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_236_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17788_ systolic_inst.A_outs\[9\]\[3\] systolic_inst.A_outs\[8\]\[3\] net117 VGND
+ VGND VPWR VPWR _01333_ sky130_fd_sc_hd__mux2_1
XFILLER_81_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19527_ systolic_inst.acc_wires\[7\]\[16\] systolic_inst.acc_wires\[7\]\[17\] systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__o21a_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16739_ _04055_ _04058_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__xnor2_1
XFILLER_235_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19458_ net105 systolic_inst.acc_wires\[7\]\[8\] net62 _06506_ VGND VGND VPWR VPWR
+ _01498_ sky130_fd_sc_hd__a22o_1
XFILLER_22_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18409_ systolic_inst.A_outs\[8\]\[6\] systolic_inst.A_shift\[16\]\[6\] net115 VGND
+ VGND VPWR VPWR _01400_ sky130_fd_sc_hd__mux2_1
XFILLER_222_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19389_ _06445_ _06446_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_187_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21420_ _08259_ _08260_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__or2_1
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_296_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_296_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21351_ _08199_ _08201_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__nand2_1
XFILLER_11_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20302_ _07239_ _07240_ _07234_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24070_ _10552_ systolic_inst.B_shift\[15\]\[6\] net71 VGND VGND VPWR VPWR _02064_
+ sky130_fd_sc_hd__mux2_1
XFILLER_163_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21282_ net63 _08140_ _08142_ systolic_inst.acc_wires\[4\]\[4\] net108 VGND VGND
+ VPWR VPWR _01686_ sky130_fd_sc_hd__a32o_1
X_23021_ _09627_ _09665_ _09664_ VGND VGND VPWR VPWR _09697_ sky130_fd_sc_hd__a21bo_1
X_20233_ systolic_inst.B_outs\[4\]\[2\] systolic_inst.B_outs\[0\]\[2\] net117 VGND
+ VGND VPWR VPWR _01596_ sky130_fd_sc_hd__mux2_1
XFILLER_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20164_ _07133_ _07134_ _07132_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__o21ai_1
XFILLER_226_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_139_Left_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27760_ clknet_leaf_212_clk _01558_ net147 VGND VGND VPWR VPWR systolic_inst.acc_wires\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20095_ _07073_ _07074_ _07075_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__and3_1
X_24972_ net111 ser_C.shift_reg\[314\] VGND VGND VPWR VPWR _10956_ sky130_fd_sc_hd__and2_1
XFILLER_131_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26711_ clknet_leaf_3_B_in_serial_clk _00514_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_23923_ _10494_ systolic_inst.B_shift\[18\]\[5\] net71 VGND VGND VPWR VPWR _01975_
+ sky130_fd_sc_hd__mux2_1
X_27691_ clknet_leaf_184_clk _01489_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_44_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_220_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_220_clk
+ sky130_fd_sc_hd__clkbuf_8
X_29430_ clknet_leaf_337_clk _03228_ net131 VGND VGND VPWR VPWR C_out\[402\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23854_ _10440_ _10442_ _10445_ _11713_ VGND VGND VPWR VPWR _10447_ sky130_fd_sc_hd__a31o_1
X_26642_ clknet_leaf_14_B_in_serial_clk _00445_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_211_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22805_ _09451_ _09486_ VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__xnor2_1
X_29361_ clknet_leaf_231_clk _03159_ net140 VGND VGND VPWR VPWR C_out\[333\] sky130_fd_sc_hd__dfrtp_1
X_23785_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[0\]\[14\]
+ VGND VGND VPWR VPWR _10388_ sky130_fd_sc_hd__nand2_1
X_26573_ clknet_leaf_25_A_in_serial_clk _00376_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_20997_ _07828_ _07831_ _07869_ net117 VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__o31ai_1
XFILLER_41_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28312_ clknet_leaf_348_clk _02110_ VGND VGND VPWR VPWR systolic_inst.A_shift\[29\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_22736_ _09401_ _09418_ _09419_ _11258_ VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_172_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25524_ systolic_inst.acc_wires\[0\]\[0\] C_out\[0\] net32 VGND VGND VPWR VPWR _02826_
+ sky130_fd_sc_hd__mux2_1
XFILLER_214_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29292_ clknet_leaf_315_clk _03090_ net142 VGND VGND VPWR VPWR C_out\[264\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_148_Left_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25455_ _00008_ _11200_ VGND VGND VPWR VPWR _11201_ sky130_fd_sc_hd__nor2_1
X_28243_ clknet_leaf_49_clk _02041_ VGND VGND VPWR VPWR systolic_inst.B_shift\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22667_ _09369_ _09372_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__or2_1
XFILLER_201_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24406_ net114 ser_C.shift_reg\[31\] VGND VGND VPWR VPWR _10673_ sky130_fd_sc_hd__and2_1
XFILLER_181_1380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21618_ _08390_ _08425_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__xor2_1
XFILLER_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28174_ clknet_leaf_75_clk _01972_ VGND VGND VPWR VPWR systolic_inst.B_shift\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25386_ _11162_ systolic_inst.A_shift\[2\]\[0\] net71 VGND VGND VPWR VPWR _02770_
+ sky130_fd_sc_hd__mux2_1
X_22598_ net109 systolic_inst.acc_wires\[2\]\[19\] net65 _09315_ VGND VGND VPWR VPWR
+ _01829_ sky130_fd_sc_hd__a22o_1
XFILLER_224_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_287_clk clknet_5_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_287_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27125_ clknet_leaf_19_clk _00923_ VGND VGND VPWR VPWR systolic_inst.A_shift\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_24337_ systolic_inst.A_shift\[8\]\[0\] net70 net83 systolic_inst.A_shift\[9\]\[0\]
+ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__a22o_1
XFILLER_194_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21549_ _08354_ _08359_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__xor2_1
XFILLER_138_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27056_ clknet_leaf_1_B_in_serial_clk _00854_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_15070_ _12153_ _12155_ _12187_ VGND VGND VPWR VPWR _12188_ sky130_fd_sc_hd__a21o_1
X_24268_ systolic_inst.B_shift\[17\]\[3\] net72 _11333_ B_in\[107\] VGND VGND VPWR
+ VPWR _02205_ sky130_fd_sc_hd__a22o_1
X_14021_ deser_B.shift_reg\[55\] deser_B.shift_reg\[56\] net125 VGND VGND VPWR VPWR
+ _00847_ sky130_fd_sc_hd__mux2_1
X_26007_ systolic_inst.acc_wires\[15\]\[3\] ser_C.parallel_data\[483\] net23 VGND
+ VGND VPWR VPWR _03309_ sky130_fd_sc_hd__mux2_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23219_ _09868_ _09869_ _09867_ VGND VGND VPWR VPWR _09870_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_112_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24199_ systolic_inst.B_shift\[22\]\[6\] net71 _11333_ B_in\[118\] VGND VGND VPWR
+ VPWR _02160_ sky130_fd_sc_hd__a22o_1
XFILLER_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18760_ _05834_ _05883_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__xnor2_1
X_27958_ clknet_leaf_170_clk _01756_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ systolic_inst.B_outs\[11\]\[5\] systolic_inst.B_outs\[7\]\[5\] net119 VGND
+ VGND VPWR VPWR _01151_ sky130_fd_sc_hd__mux2_1
XFILLER_96_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17711_ _04920_ _04925_ _04930_ _04934_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__or4_1
XFILLER_209_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14923_ _12041_ _12044_ VGND VGND VPWR VPWR _12045_ sky130_fd_sc_hd__xnor2_1
X_26909_ clknet_leaf_11_A_in_serial_clk _00707_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_18691_ _05777_ _05779_ _05816_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_86_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27889_ clknet_leaf_309_clk _01687_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_236_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_211_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_211_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29628_ clknet_leaf_9_B_in_serial_clk _03423_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_208_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17642_ _04878_ _04880_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__nand2_1
XFILLER_1_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14854_ _11973_ _11974_ _11976_ VGND VGND VPWR VPWR _11978_ sky130_fd_sc_hd__or3_1
XFILLER_208_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13805_ B_in\[112\] deser_B.word_buffer\[112\] net88 VGND VGND VPWR VPWR _00642_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29559_ clknet_leaf_14_B_in_serial_clk _03354_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17573_ net118 _04812_ _04822_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__and3_1
XFILLER_21_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14785_ _11909_ _11910_ VGND VGND VPWR VPWR _11912_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_231_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_231_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19312_ _06237_ _06372_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__or2_1
XFILLER_147_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16524_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__inv_2
XFILLER_1_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13736_ B_in\[43\] deser_B.word_buffer\[43\] net84 VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19243_ _06238_ _06305_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__nor2_1
XFILLER_91_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16455_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[12\]\[13\]
+ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__or2_1
XFILLER_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13667_ deser_B.word_buffer\[103\] deser_B.serial_word\[103\] net123 VGND VGND VPWR
+ VPWR _00504_ sky130_fd_sc_hd__mux2_1
XFILLER_32_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15406_ systolic_inst.B_outs\[13\]\[1\] systolic_inst.A_outs\[13\]\[3\] systolic_inst.A_outs\[13\]\[4\]
+ systolic_inst.B_outs\[13\]\[0\] VGND VGND VPWR VPWR _12468_ sky130_fd_sc_hd__a22o_1
X_19174_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] _06238_ VGND
+ VGND VPWR VPWR _06239_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_26_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13598_ deser_B.word_buffer\[34\] deser_B.serial_word\[34\] net124 VGND VGND VPWR
+ VPWR _00435_ sky130_fd_sc_hd__mux2_1
X_16386_ _03751_ _03754_ _03756_ _03758_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_26_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_278_clk clknet_5_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_278_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18125_ _05311_ _05312_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__and2_1
XFILLER_145_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15337_ _12419_ _12422_ VGND VGND VPWR VPWR _12423_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_229_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1 _10481_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18056_ _05245_ _05246_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__nand2_1
XFILLER_144_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15268_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[18\]
+ VGND VGND VPWR VPWR _12364_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_10_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_225_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17007_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[6\] systolic_inst.acc_wires\[11\]\[6\]
+ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__nand2_1
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14219_ _11405_ _11406_ VGND VGND VPWR VPWR _11407_ sky130_fd_sc_hd__or2_1
X_15199_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[14\]\[8\]
+ VGND VGND VPWR VPWR _12305_ sky130_fd_sc_hd__and2_1
XFILLER_154_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18958_ _06048_ _06052_ _06055_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__nand3_1
XFILLER_140_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17909_ _05101_ _05102_ _05071_ _05074_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_176_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18889_ _05984_ _05987_ _05990_ _05995_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__a211o_1
XFILLER_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_176_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_202_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_202_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_176_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20920_ _07793_ _07794_ _07795_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__nor3b_1
XFILLER_39_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20851_ _07729_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__inv_2
XFILLER_187_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23570_ systolic_inst.B_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[7\]
+ VGND VGND VPWR VPWR _10192_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20782_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[24\]
+ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__and2_1
XFILLER_211_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22521_ _09248_ _09249_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__and2_1
XFILLER_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25240_ net111 ser_C.shift_reg\[448\] VGND VGND VPWR VPWR _11090_ sky130_fd_sc_hd__and2_1
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22452_ _09188_ _09189_ VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__and2b_1
XFILLER_50_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21403_ _08244_ _08245_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_269_clk clknet_5_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_269_clk
+ sky130_fd_sc_hd__clkbuf_8
X_25171_ C_out\[412\] net101 net73 ser_C.shift_reg\[412\] _11055_ VGND VGND VPWR VPWR
+ _02662_ sky130_fd_sc_hd__a221o_1
X_22383_ _08984_ _09122_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__nand2_1
XFILLER_148_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24122_ _10562_ systolic_inst.A_shift\[29\]\[0\] net71 VGND VGND VPWR VPWR _02106_
+ sky130_fd_sc_hd__mux2_1
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21334_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[4\]\[12\]
+ VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__or2_1
XFILLER_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24053_ systolic_inst.B_shift\[4\]\[6\] B_in\[6\] _00008_ VGND VGND VPWR VPWR _10544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28930_ clknet_leaf_265_clk _02728_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[478\]
+ sky130_fd_sc_hd__dfrtp_1
X_21265_ _08126_ _08127_ _08119_ _08122_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__a211o_1
XFILLER_237_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23004_ _09678_ _09680_ VGND VGND VPWR VPWR _09681_ sky130_fd_sc_hd__nand2_1
XFILLER_137_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20216_ _07175_ _07178_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__nand2_1
XFILLER_143_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28861_ clknet_leaf_332_clk _02659_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[409\]
+ sky130_fd_sc_hd__dfrtp_1
X_21196_ _08031_ _08034_ _08032_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_161_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27812_ clknet_leaf_140_clk _01610_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_235_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20147_ _07118_ _07119_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_161_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28792_ clknet_leaf_233_clk _02590_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_213_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27743_ clknet_leaf_213_clk _01541_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20078_ _07059_ _07060_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__and2_1
XFILLER_131_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24955_ C_out\[304\] net103 net76 ser_C.shift_reg\[304\] _10947_ VGND VGND VPWR VPWR
+ _02554_ sky130_fd_sc_hd__a221o_1
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23906_ systolic_inst.B_shift\[17\]\[5\] B_in\[77\] _00008_ VGND VGND VPWR VPWR _10486_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27674_ clknet_leaf_147_clk _01472_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_2_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24886_ net110 ser_C.shift_reg\[271\] VGND VGND VPWR VPWR _10913_ sky130_fd_sc_hd__and2_1
XFILLER_218_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29413_ clknet_leaf_327_clk _03211_ net136 VGND VGND VPWR VPWR C_out\[385\] sky130_fd_sc_hd__dfrtp_1
X_26625_ clknet_leaf_23_B_in_serial_clk _00428_ net137 VGND VGND VPWR VPWR deser_B.word_buffer\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23837_ _10424_ _10425_ VGND VGND VPWR VPWR _10432_ sky130_fd_sc_hd__and2b_1
XFILLER_57_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29344_ clknet_leaf_213_clk _03142_ net149 VGND VGND VPWR VPWR C_out\[316\] sky130_fd_sc_hd__dfrtp_1
X_14570_ _11739_ _11740_ _11741_ VGND VGND VPWR VPWR _11742_ sky130_fd_sc_hd__a21o_1
XFILLER_54_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23768_ _10363_ _10368_ _10369_ VGND VGND VPWR VPWR _10373_ sky130_fd_sc_hd__nand3_1
X_26556_ clknet_leaf_27_A_in_serial_clk _00359_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_220_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25507_ _11233_ _11234_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__nor2_1
XFILLER_198_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13521_ deser_A.shift_reg\[85\] deser_A.shift_reg\[86\] net129 VGND VGND VPWR VPWR
+ _00358_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22719_ systolic_inst.A_outs\[1\]\[0\] systolic_inst.A_outs\[1\]\[1\] systolic_inst.B_outs\[1\]\[3\]
+ systolic_inst.B_outs\[1\]\[4\] VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__nand4_1
X_29275_ clknet_leaf_188_clk _03073_ net146 VGND VGND VPWR VPWR C_out\[247\] sky130_fd_sc_hd__dfrtp_1
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23699_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[0\]\[0\]
+ _10311_ _10312_ VGND VGND VPWR VPWR _10315_ sky130_fd_sc_hd__a22o_1
X_26487_ clknet_leaf_8_A_in_serial_clk _00290_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_242_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28226_ clknet_leaf_97_clk _02024_ VGND VGND VPWR VPWR systolic_inst.B_shift\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13452_ deser_A.shift_reg\[16\] deser_A.shift_reg\[17\] deser_A.receiving VGND VGND
+ VPWR VPWR _00289_ sky130_fd_sc_hd__mux2_1
X_16240_ _03548_ _03584_ _03621_ _03622_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__o211ai_1
X_25438_ _11257_ _11258_ _11186_ VGND VGND VPWR VPWR _11189_ sky130_fd_sc_hd__or3_1
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28157_ clknet_leaf_107_clk _01955_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_25369_ systolic_inst.B_shift\[18\]\[0\] B_in\[48\] _00008_ VGND VGND VPWR VPWR _11154_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16171_ _03514_ _03520_ _03519_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__a21o_1
X_13383_ A_in\[92\] deser_A.word_buffer\[92\] net92 VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__mux2_1
XFILLER_127_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27108_ clknet_leaf_2_B_in_serial_clk _00906_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15122_ _12211_ _12214_ _12237_ VGND VGND VPWR VPWR _12238_ sky130_fd_sc_hd__a21oi_1
XFILLER_103_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28088_ clknet_leaf_117_clk _01886_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19930_ _06925_ _06926_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__nor2_1
X_15053_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[11\] VGND
+ VGND VPWR VPWR _12172_ sky130_fd_sc_hd__and2_1
X_27039_ clknet_leaf_14_B_in_serial_clk _00837_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14004_ deser_B.shift_reg\[38\] deser_B.shift_reg\[39\] deser_B.receiving VGND VGND
+ VPWR VPWR _00830_ sky130_fd_sc_hd__mux2_1
X_19861_ _06825_ _06859_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_220_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18812_ _05929_ _05930_ _05922_ _05925_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__a211o_1
X_19792_ systolic_inst.A_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[5\] VGND VGND VPWR
+ VPWR _06793_ sky130_fd_sc_hd__nand2_1
XFILLER_122_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18743_ _05864_ _05865_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nor2_1
X_15955_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[31\]
+ VGND VGND VPWR VPWR _12974_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14906_ systolic_inst.B_outs\[14\]\[7\] _11993_ _11994_ VGND VGND VPWR VPWR _12028_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_188_1342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18674_ systolic_inst.A_outs\[8\]\[6\] _05768_ _05769_ _05735_ VGND VGND VPWR VPWR
+ _05800_ sky130_fd_sc_hd__o2bb2a_1
X_15886_ _12894_ _12915_ VGND VGND VPWR VPWR _12916_ sky130_fd_sc_hd__nor2_1
XFILLER_110_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17625_ _11712_ _04865_ _04866_ systolic_inst.acc_wires\[10\]\[7\] net105 VGND VGND
+ VPWR VPWR _01305_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_218_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14837_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[3\] _11945_ _11944_
+ VGND VGND VPWR VPWR _11961_ sky130_fd_sc_hd__a31o_1
XFILLER_188_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_218_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17556_ _04806_ _04805_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_28_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14768_ systolic_inst.A_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[2\] VGND VGND
+ VPWR VPWR _11896_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16507_ systolic_inst.acc_wires\[12\]\[16\] systolic_inst.acc_wires\[12\]\[17\] systolic_inst.acc_wires\[12\]\[18\]
+ systolic_inst.acc_wires\[12\]\[19\] systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__o41a_1
XFILLER_71_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13719_ B_in\[26\] deser_B.word_buffer\[26\] net85 VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__mux2_1
XFILLER_204_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17487_ _04601_ _04738_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__nand2_2
X_14699_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[15\]\[25\]
+ VGND VGND VPWR VPWR _11852_ sky130_fd_sc_hd__xor2_2
XFILLER_225_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19226_ _06281_ _06289_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__xnor2_1
X_16438_ _03801_ _03802_ _03803_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_15_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19157_ _06184_ _06220_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__xor2_1
X_16369_ _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__inv_2
XFILLER_121_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18108_ _05295_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__xnor2_1
X_19088_ _06154_ _06155_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[5\]
+ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__and4bb_1
XFILLER_195_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18039_ _05228_ _05229_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21050_ _07920_ _07921_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20001_ _06944_ _06972_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__or2_1
XFILLER_87_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_203_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_199_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21952_ net68 _08739_ _08740_ systolic_inst.acc_wires\[3\]\[12\] net106 VGND VGND
+ VPWR VPWR _01758_ sky130_fd_sc_hd__a32o_1
X_24740_ net112 ser_C.shift_reg\[198\] VGND VGND VPWR VPWR _10840_ sky130_fd_sc_hd__and2_1
XFILLER_28_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ _07750_ _07777_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_195_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24671_ C_out\[162\] net103 net76 ser_C.shift_reg\[162\] _10805_ VGND VGND VPWR VPWR
+ _02412_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21883_ net68 _08679_ _08681_ systolic_inst.acc_wires\[3\]\[2\] net106 VGND VGND
+ VPWR VPWR _01748_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_195_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23622_ _10241_ _10242_ VGND VGND VPWR VPWR _10243_ sky130_fd_sc_hd__and2_1
X_26410_ clknet_leaf_4_clk _00217_ net131 VGND VGND VPWR VPWR A_in\[78\] sky130_fd_sc_hd__dfrtp_1
X_20834_ systolic_inst.A_outs\[4\]\[7\] systolic_inst.A_shift\[8\]\[7\] net121 VGND
+ VGND VPWR VPWR _01657_ sky130_fd_sc_hd__mux2_1
X_27390_ clknet_leaf_337_clk _01188_ net131 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23553_ _10109_ _10111_ _10172_ _10174_ VGND VGND VPWR VPWR _10176_ sky130_fd_sc_hd__a211o_1
X_26341_ clknet_leaf_59_clk _00148_ net144 VGND VGND VPWR VPWR A_in\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20765_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[22\]
+ VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_154_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22504_ _09235_ VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__inv_2
XFILLER_168_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29060_ clknet_leaf_108_clk _02858_ net150 VGND VGND VPWR VPWR C_out\[32\] sky130_fd_sc_hd__dfrtp_1
XFILLER_211_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26272_ clknet_leaf_21_A_in_serial_clk _00080_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_210_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23484_ _10106_ _10107_ VGND VGND VPWR VPWR _10108_ sky130_fd_sc_hd__nor2_1
XFILLER_161_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20696_ _07603_ _07608_ _07609_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_150_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28011_ clknet_leaf_149_clk _01809_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_202_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25223_ C_out\[438\] net101 net73 ser_C.shift_reg\[438\] _11081_ VGND VGND VPWR VPWR
+ _02688_ sky130_fd_sc_hd__a221o_1
X_22435_ _09142_ _09145_ _09173_ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__or3_1
XFILLER_195_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25154_ net110 ser_C.shift_reg\[405\] VGND VGND VPWR VPWR _11047_ sky130_fd_sc_hd__and2_1
XFILLER_100_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22366_ _09069_ _09071_ _09106_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__nand3_1
XFILLER_191_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24105_ systolic_inst.B_shift\[1\]\[0\] _11332_ net83 systolic_inst.B_shift\[5\]\[0\]
+ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__a22o_1
X_21317_ _08170_ _08171_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__nand2_1
XFILLER_124_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25085_ C_out\[369\] net98 net78 ser_C.shift_reg\[369\] _11012_ VGND VGND VPWR VPWR
+ _02619_ sky130_fd_sc_hd__a221o_1
X_22297_ _09039_ _09040_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__nand2_1
XFILLER_2_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24036_ _10535_ systolic_inst.B_shift\[4\]\[5\] net72 VGND VGND VPWR VPWR _02047_
+ sky130_fd_sc_hd__mux2_1
X_28913_ clknet_leaf_284_clk _02711_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[461\]
+ sky130_fd_sc_hd__dfrtp_1
X_21248_ _08100_ _08101_ _08073_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__mux2_1
XFILLER_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28844_ clknet_leaf_333_clk _02642_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[392\]
+ sky130_fd_sc_hd__dfrtp_1
X_21179_ _07997_ _08014_ _08013_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__o21ba_1
XFILLER_120_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28775_ clknet_leaf_251_clk _02573_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[323\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25987_ systolic_inst.acc_wires\[14\]\[15\] ser_C.parallel_data\[463\] net26 VGND
+ VGND VPWR VPWR _03289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27726_ clknet_leaf_215_clk _01524_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_15740_ _12789_ _12791_ VGND VGND VPWR VPWR _12792_ sky130_fd_sc_hd__nand2_1
XFILLER_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24938_ net111 ser_C.shift_reg\[297\] VGND VGND VPWR VPWR _10939_ sky130_fd_sc_hd__and2_1
XFILLER_234_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _12722_ _12723_ VGND VGND VPWR VPWR _12725_ sky130_fd_sc_hd__xnor2_1
X_27657_ clknet_leaf_301_clk _01455_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_24869_ C_out\[261\] net101 net73 ser_C.shift_reg\[261\] _10904_ VGND VGND VPWR VPWR
+ _02511_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_103_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _04627_ _04629_ _04664_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__nand3_1
X_26608_ clknet_leaf_15_B_in_serial_clk _00411_ net152 VGND VGND VPWR VPWR deser_B.word_buffer\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14622_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[15\]\[14\]
+ VGND VGND VPWR VPWR _11786_ sky130_fd_sc_hd__or2_1
X_18390_ net105 systolic_inst.acc_wires\[9\]\[29\] net66 _05545_ VGND VGND VPWR VPWR
+ _01391_ sky130_fd_sc_hd__a22o_1
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27588_ clknet_leaf_216_clk _01386_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17341_ _04533_ _04569_ _04568_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__a21bo_1
X_29327_ clknet_leaf_221_clk _03125_ net139 VGND VGND VPWR VPWR C_out\[299\] sky130_fd_sc_hd__dfrtp_1
XFILLER_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14553_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[4\] systolic_inst.acc_wires\[15\]\[4\]
+ VGND VGND VPWR VPWR _11727_ sky130_fd_sc_hd__nand2_1
XFILLER_42_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26539_ clknet_leaf_21_A_in_serial_clk _00342_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13504_ deser_A.shift_reg\[68\] deser_A.shift_reg\[69\] net129 VGND VGND VPWR VPWR
+ _00341_ sky130_fd_sc_hd__mux2_1
X_29258_ clknet_leaf_196_clk _03056_ net146 VGND VGND VPWR VPWR C_out\[230\] sky130_fd_sc_hd__dfrtp_1
X_17272_ _04513_ _04515_ _04514_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_12_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14484_ _11622_ _11664_ VGND VGND VPWR VPWR _11665_ sky130_fd_sc_hd__xor2_1
XFILLER_186_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19011_ systolic_inst.A_outs\[7\]\[0\] systolic_inst.A_outs\[6\]\[0\] net119 VGND
+ VGND VPWR VPWR _01458_ sky130_fd_sc_hd__mux2_1
X_28209_ clknet_leaf_98_clk _02007_ VGND VGND VPWR VPWR systolic_inst.B_shift\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16223_ _03596_ _03604_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__or2_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13435_ deser_A.bit_idx\[5\] _11316_ deser_A.bit_idx\[6\] VGND VGND VPWR VPWR _11318_
+ sky130_fd_sc_hd__a21o_1
X_29189_ clknet_leaf_307_clk _02987_ net141 VGND VGND VPWR VPWR C_out\[161\] sky130_fd_sc_hd__dfrtp_1
XFILLER_228_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload207 clknet_leaf_37_clk VGND VGND VPWR VPWR clkload207/Y sky130_fd_sc_hd__inv_8
Xclkload218 clknet_leaf_50_clk VGND VGND VPWR VPWR clkload218/Y sky130_fd_sc_hd__clkinv_8
XFILLER_139_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload229 clknet_leaf_73_clk VGND VGND VPWR VPWR clkload229/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16154_ _03521_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__or2_1
X_13366_ A_in\[75\] deser_A.word_buffer\[75\] net94 VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__mux2_1
XFILLER_170_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15105_ _12221_ _12220_ VGND VGND VPWR VPWR _12222_ sky130_fd_sc_hd__and2b_1
X_13297_ A_in\[6\] deser_A.word_buffer\[6\] net94 VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__mux2_1
X_16085_ _13079_ _13080_ _13054_ VGND VGND VPWR VPWR _13081_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19913_ _06910_ _06909_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__and2b_1
X_15036_ _12146_ _12154_ VGND VGND VPWR VPWR _12155_ sky130_fd_sc_hd__nand2_1
XFILLER_64_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19844_ _06843_ _06842_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__nand2b_1
XFILLER_116_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19775_ _06736_ _06739_ _06775_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_53_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16987_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[11\]\[3\]
+ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__or2_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18726_ _05848_ _05849_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__xnor2_1
XFILLER_225_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15938_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[28\]
+ VGND VGND VPWR VPWR _12960_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18657_ _05781_ _05782_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__xor2_1
X_15869_ _12899_ _12901_ VGND VGND VPWR VPWR _12902_ sky130_fd_sc_hd__xnor2_1
Xwire37 net39 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_8
XFILLER_240_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17608_ _04845_ _04846_ _04844_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__a21bo_1
XFILLER_24_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18588_ _05699_ _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__xor2_1
XFILLER_240_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17539_ _04758_ _04760_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__nor3_1
XFILLER_71_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20550_ _07430_ _07482_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__and2_1
XFILLER_225_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19209_ _06244_ _06246_ _06243_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20481_ _07377_ _07378_ _07380_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__o21a_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22220_ _08959_ _08965_ VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__nor2_1
XFILLER_160_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22151_ systolic_inst.A_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[3\] systolic_inst.B_outs\[2\]\[4\]
+ systolic_inst.A_outs\[2\]\[1\] VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_209_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_209_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21102_ _07971_ _07972_ VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__and2b_1
XFILLER_156_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22082_ systolic_inst.A_outs\[2\]\[4\] systolic_inst.A_outs\[1\]\[4\] net122 VGND
+ VGND VPWR VPWR _01782_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_205_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25910_ systolic_inst.acc_wires\[12\]\[2\] C_out\[386\] net21 VGND VGND VPWR VPWR
+ _03212_ sky130_fd_sc_hd__mux2_1
XFILLER_59_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21033_ _07872_ _07904_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__xor2_1
XFILLER_160_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26890_ clknet_leaf_6_A_in_serial_clk _00688_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25841_ systolic_inst.acc_wires\[9\]\[29\] C_out\[317\] net12 VGND VGND VPWR VPWR
+ _03143_ sky130_fd_sc_hd__mux2_1
XFILLER_234_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_197_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28560_ clknet_leaf_168_clk _02358_ net148 VGND VGND VPWR VPWR ser_C.shift_reg\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22984_ systolic_inst.B_outs\[1\]\[5\] systolic_inst.A_outs\[1\]\[7\] _09659_ VGND
+ VGND VPWR VPWR _09661_ sky130_fd_sc_hd__and3_1
X_25772_ systolic_inst.acc_wires\[7\]\[24\] C_out\[248\] net44 VGND VGND VPWR VPWR
+ _03074_ sky130_fd_sc_hd__mux2_1
XFILLER_234_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_18_A_in_serial_clk clknet_2_3__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_18_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_227_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27511_ clknet_leaf_231_clk _01309_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_24723_ C_out\[188\] net99 net79 ser_C.shift_reg\[188\] _10831_ VGND VGND VPWR VPWR
+ _02438_ sky130_fd_sc_hd__a221o_1
X_28491_ clknet_leaf_116_clk _02289_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_21935_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[3\]\[11\]
+ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__or2_1
XFILLER_43_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27442_ clknet_leaf_243_clk _01240_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_242_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21866_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] _08660_
+ _08667_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__a22o_1
X_24654_ net7 ser_C.shift_reg\[155\] VGND VGND VPWR VPWR _10797_ sky130_fd_sc_hd__and2_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20817_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[30\]
+ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__nand2_1
X_23605_ _10186_ _10225_ VGND VGND VPWR VPWR _10226_ sky130_fd_sc_hd__or2_1
XFILLER_242_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27373_ clknet_leaf_327_clk _01171_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24585_ C_out\[119\] net100 net82 ser_C.shift_reg\[119\] _10762_ VGND VGND VPWR VPWR
+ _02369_ sky130_fd_sc_hd__a221o_1
XFILLER_208_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21797_ _08601_ _08600_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__and2b_1
XFILLER_230_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29112_ clknet_leaf_158_clk _02910_ net150 VGND VGND VPWR VPWR C_out\[84\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26324_ clknet_leaf_30_A_in_serial_clk _00132_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_184_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20748_ _07656_ _07657_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__xnor2_1
X_23536_ systolic_inst.A_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[7\] VGND VGND VPWR
+ VPWR _10159_ sky130_fd_sc_hd__nand2b_1
XFILLER_208_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29043_ clknet_leaf_99_clk _02841_ net152 VGND VGND VPWR VPWR C_out\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23467_ _10072_ _10089_ _10090_ VGND VGND VPWR VPWR _10092_ sky130_fd_sc_hd__nand3_1
XFILLER_17_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26255_ clknet_leaf_4_A_in_serial_clk _00063_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_183_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20679_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[5\]\[8\]
+ _07595_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__and3_1
XFILLER_137_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13220_ deser_A.word_buffer\[58\] deser_A.serial_word\[58\] net128 VGND VGND VPWR
+ VPWR _00068_ sky130_fd_sc_hd__mux2_1
X_22418_ _09130_ _09156_ VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__xnor2_1
X_25206_ net110 ser_C.shift_reg\[431\] VGND VGND VPWR VPWR _11073_ sky130_fd_sc_hd__and2_1
XFILLER_195_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26186_ ser_C.bit_idx\[5\] _11250_ _11303_ VGND VGND VPWR VPWR _11253_ sky130_fd_sc_hd__o21ai_1
X_23398_ _09998_ _10001_ _09999_ VGND VGND VPWR VPWR _10024_ sky130_fd_sc_hd__o21ba_1
XFILLER_178_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13151_ net7 net10 VGND VGND VPWR VPWR _11303_ sky130_fd_sc_hd__nand2b_1
XFILLER_192_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22349_ _08985_ _09090_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__or2_1
XFILLER_152_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25137_ C_out\[395\] net101 net73 ser_C.shift_reg\[395\] _11038_ VGND VGND VPWR VPWR
+ _02645_ sky130_fd_sc_hd__a221o_1
XFILLER_128_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25068_ net112 ser_C.shift_reg\[362\] VGND VGND VPWR VPWR _11004_ sky130_fd_sc_hd__and2_1
XFILLER_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_215_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24019_ systolic_inst.B_shift\[6\]\[2\] _11332_ net83 systolic_inst.B_shift\[10\]\[2\]
+ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__a22o_1
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16910_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[12\] _04226_ net119
+ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17890_ _05053_ _05083_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__nor2_1
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28827_ clknet_leaf_238_clk _02625_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[375\]
+ sky130_fd_sc_hd__dfrtp_1
X_16841_ _04157_ _04158_ _04159_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__and3_1
XFILLER_238_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19560_ _06585_ _06589_ _06592_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__a21o_1
XFILLER_65_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28758_ clknet_leaf_219_clk _02556_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[306\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16772_ _04054_ _04060_ _04059_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a21o_1
X_13984_ deser_B.shift_reg\[18\] deser_B.shift_reg\[19\] net125 VGND VGND VPWR VPWR
+ _00810_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18511_ _05635_ _05636_ _05640_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__a21o_1
XFILLER_185_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27709_ clknet_leaf_194_clk _01507_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_15723_ _12687_ _12774_ VGND VGND VPWR VPWR _12775_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_215_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19491_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[7\]\[12\]
+ _06532_ _06534_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__a211o_1
XFILLER_20_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28689_ clknet_leaf_191_clk _02487_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[237\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18442_ _05570_ _05575_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__nand2_1
X_15654_ _12707_ _12708_ VGND VGND VPWR VPWR _12709_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_17_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ net105 systolic_inst.acc_wires\[15\]\[11\] net69 _11771_ VGND VGND VPWR VPWR
+ _00989_ sky130_fd_sc_hd__a22o_1
X_18373_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[27\]
+ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15585_ _12605_ _12608_ _12640_ net115 VGND VGND VPWR VPWR _12642_ sky130_fd_sc_hd__o31a_1
XFILLER_226_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17324_ _04544_ _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__xnor2_1
XFILLER_222_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14536_ net107 systolic_inst.load_acc VGND VGND VPWR VPWR _11713_ sky130_fd_sc_hd__or2_4
XFILLER_105_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_239_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_230_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17255_ systolic_inst.A_outs\[10\]\[2\] systolic_inst.B_outs\[10\]\[3\] systolic_inst.B_outs\[10\]\[4\]
+ systolic_inst.A_outs\[10\]\[1\] VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__a22o_1
XFILLER_30_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14467_ _11647_ _11648_ VGND VGND VPWR VPWR _11649_ sky130_fd_sc_hd__nor2_1
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16206_ _03560_ _03561_ _03562_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__o21ba_1
XFILLER_70_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13418_ A_in\[127\] deser_A.word_buffer\[127\] net92 VGND VGND VPWR VPWR _00266_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17186_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[5\]\[0\] net116 VGND
+ VGND VPWR VPWR _01274_ sky130_fd_sc_hd__mux2_1
X_14398_ _11508_ _11510_ _11547_ _11548_ VGND VGND VPWR VPWR _11582_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_180_Right_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16137_ systolic_inst.B_outs\[12\]\[3\] systolic_inst.B_outs\[12\]\[4\] systolic_inst.A_outs\[12\]\[4\]
+ systolic_inst.A_outs\[12\]\[5\] VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__and4_1
XFILLER_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13349_ A_in\[58\] deser_A.word_buffer\[58\] net91 VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16068_ systolic_inst.A_outs\[12\]\[2\] systolic_inst.B_outs\[12\]\[3\] systolic_inst.A_outs\[12\]\[3\]
+ systolic_inst.B_outs\[12\]\[4\] VGND VGND VPWR VPWR _13064_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_55_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15019_ _12137_ _12138_ VGND VGND VPWR VPWR _12139_ sky130_fd_sc_hd__nor2_1
XFILLER_116_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19827_ systolic_inst.B_outs\[6\]\[3\] systolic_inst.B_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[5\]
+ systolic_inst.A_outs\[6\]\[6\] VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_200_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19758_ _06726_ _06758_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__xnor2_1
XFILLER_238_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_192_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18709_ _05694_ _05832_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_192_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19689_ systolic_inst.A_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[5\] VGND VGND VPWR
+ VPWR _06693_ sky130_fd_sc_hd__nand2_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21720_ _08490_ _08492_ _08491_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__o21ba_1
XFILLER_80_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21651_ _08457_ _08458_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_111_Left_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20602_ _07532_ _07531_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__and2b_1
XFILLER_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24370_ net7 ser_C.shift_reg\[13\] VGND VGND VPWR VPWR _10655_ sky130_fd_sc_hd__and2_1
XFILLER_127_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21582_ _08380_ _08392_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23321_ _09931_ _09948_ _09949_ VGND VGND VPWR VPWR _09950_ sky130_fd_sc_hd__nand3b_1
XFILLER_177_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20533_ systolic_inst.B_outs\[5\]\[6\] systolic_inst.A_outs\[5\]\[6\] _11276_ systolic_inst.A_outs\[5\]\[5\]
+ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23252_ _09890_ _09894_ VGND VGND VPWR VPWR _09897_ sky130_fd_sc_hd__nor2_1
XFILLER_193_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26040_ systolic_inst.B_outs\[15\]\[4\] systolic_inst.B_outs\[11\]\[4\] net118 VGND
+ VGND VPWR VPWR _03342_ sky130_fd_sc_hd__mux2_1
X_20464_ systolic_inst.A_outs\[5\]\[6\] _07398_ _07397_ VGND VGND VPWR VPWR _07399_
+ sky130_fd_sc_hd__a21bo_1
X_22203_ systolic_inst.B_outs\[2\]\[0\] systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[6\]
+ systolic_inst.A_outs\[2\]\[7\] VGND VGND VPWR VPWR _08949_ sky130_fd_sc_hd__nand4_1
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23183_ net109 systolic_inst.acc_wires\[1\]\[16\] _09837_ _09839_ VGND VGND VPWR
+ VPWR _01890_ sky130_fd_sc_hd__a22o_1
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20395_ _07331_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__inv_2
X_22134_ _08862_ _08880_ _08881_ VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__or3_1
XFILLER_134_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27991_ clknet_leaf_121_clk _01789_ net152 VGND VGND VPWR VPWR systolic_inst.B_outs\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_145_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_120_Left_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22065_ _08829_ _08832_ _08836_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__o21ai_1
X_26942_ clknet_leaf_19_A_in_serial_clk _00740_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21016_ systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[7\] VGND VGND VPWR
+ VPWR _07889_ sky130_fd_sc_hd__and2b_1
XFILLER_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29661_ clknet_leaf_10_B_in_serial_clk _03456_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_26873_ clknet_leaf_15_A_in_serial_clk _00671_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28612_ clknet_leaf_40_clk _02410_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[160\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25824_ systolic_inst.acc_wires\[9\]\[12\] C_out\[300\] net15 VGND VGND VPWR VPWR
+ _03126_ sky130_fd_sc_hd__mux2_1
X_29592_ clknet_leaf_13_B_in_serial_clk _03387_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28543_ clknet_leaf_164_clk _02341_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_25755_ systolic_inst.acc_wires\[7\]\[7\] C_out\[231\] net42 VGND VGND VPWR VPWR
+ _03057_ sky130_fd_sc_hd__mux2_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22967_ _09643_ _09644_ VGND VGND VPWR VPWR _09645_ sky130_fd_sc_hd__nor2_1
XFILLER_55_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24706_ net113 ser_C.shift_reg\[181\] VGND VGND VPWR VPWR _10823_ sky130_fd_sc_hd__and2_1
X_28474_ clknet_leaf_103_clk _02272_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_21918_ _08706_ _08709_ _08710_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25686_ systolic_inst.acc_wires\[5\]\[2\] C_out\[162\] net16 VGND VGND VPWR VPWR
+ _02988_ sky130_fd_sc_hd__mux2_1
X_22898_ _09575_ _09576_ VGND VGND VPWR VPWR _09578_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27425_ clknet_leaf_249_clk _01223_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_231_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_175_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24637_ C_out\[145\] net103 net76 ser_C.shift_reg\[145\] _10788_ VGND VGND VPWR VPWR
+ _02395_ sky130_fd_sc_hd__a221o_1
X_21849_ _08649_ _08650_ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_175_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27356_ clknet_leaf_323_clk _01154_ net136 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15370_ systolic_inst.B_outs\[12\]\[6\] systolic_inst.B_outs\[8\]\[6\] net115 VGND
+ VGND VPWR VPWR _01088_ sky130_fd_sc_hd__mux2_1
X_24568_ net113 ser_C.shift_reg\[112\] VGND VGND VPWR VPWR _10754_ sky130_fd_sc_hd__and2_1
XFILLER_145_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14321_ _11436_ _11467_ _11466_ VGND VGND VPWR VPWR _11507_ sky130_fd_sc_hd__a21oi_1
X_26307_ clknet_leaf_25_A_in_serial_clk _00115_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23519_ _10140_ _10141_ net121 VGND VGND VPWR VPWR _10143_ sky130_fd_sc_hd__o21ai_1
XFILLER_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27287_ clknet_leaf_320_clk _01085_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_24499_ C_out\[76\] net100 net80 ser_C.shift_reg\[76\] _10719_ VGND VGND VPWR VPWR
+ _02326_ sky130_fd_sc_hd__a221o_1
XFILLER_139_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29026_ clknet_leaf_92_clk _02824_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[11\]\[11\]
+ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__or2_1
X_14252_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[5\]
+ systolic_inst.A_outs\[15\]\[6\] VGND VGND VPWR VPWR _11439_ sky130_fd_sc_hd__and4_1
X_26238_ clknet_leaf_16_A_in_serial_clk _00046_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13203_ deser_A.word_buffer\[41\] deser_A.serial_word\[41\] net127 VGND VGND VPWR
+ VPWR _00051_ sky130_fd_sc_hd__mux2_1
XFILLER_137_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26169_ deser_B.serial_word\[124\] deser_B.shift_reg\[124\] net56 VGND VGND VPWR
+ VPWR _03471_ sky130_fd_sc_hd__mux2_1
X_14183_ _11371_ _11372_ VGND VGND VPWR VPWR _11373_ sky130_fd_sc_hd__nand2_1
XFILLER_174_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13134_ systolic_inst.cycle_cnt\[27\] systolic_inst.cycle_cnt\[26\] systolic_inst.cycle_cnt\[25\]
+ systolic_inst.cycle_cnt\[24\] VGND VGND VPWR VPWR _11287_ sky130_fd_sc_hd__or4_1
XFILLER_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18991_ _06082_ _06083_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__nand2_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_240_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17942_ _05084_ _05085_ _05098_ _05097_ _05065_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__o32a_1
XFILLER_139_1199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17873_ _05058_ _05066_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_128_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19612_ systolic_inst.A_outs\[6\]\[0\] systolic_inst.A_outs\[5\]\[0\] net120 VGND
+ VGND VPWR VPWR _01522_ sky130_fd_sc_hd__mux2_1
X_16824_ _04134_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__nand2_1
XFILLER_152_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19543_ net62 _06578_ _06579_ systolic_inst.acc_wires\[7\]\[20\] net105 VGND VGND
+ VPWR VPWR _01510_ sky130_fd_sc_hd__a32o_1
XFILLER_24_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16755_ _04001_ _04036_ _04038_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__a21oi_1
X_13967_ deser_B.shift_reg\[1\] deser_B.shift_reg\[2\] net125 VGND VGND VPWR VPWR
+ _00793_ sky130_fd_sc_hd__mux2_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_238_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15706_ _12756_ _12757_ VGND VGND VPWR VPWR _12759_ sky130_fd_sc_hd__xor2_1
X_19474_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[7\]\[11\]
+ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__or2_1
XFILLER_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16686_ _03978_ _04007_ _04008_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__nand3_1
XFILLER_34_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13898_ deser_A.serial_word\[59\] deser_A.shift_reg\[59\] _00002_ VGND VGND VPWR
+ VPWR _00724_ sky130_fd_sc_hd__mux2_1
XFILLER_55_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_234_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18425_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[2\] VGND
+ VGND VPWR VPWR _05560_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_234_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15637_ _12688_ _12691_ VGND VGND VPWR VPWR _12692_ sky130_fd_sc_hd__xor2_1
XFILLER_181_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18356_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[24\]
+ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_44_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _12621_ _12624_ VGND VGND VPWR VPWR _12625_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17307_ systolic_inst.B_outs\[10\]\[0\] systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[6\]
+ systolic_inst.A_outs\[10\]\[7\] VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__nand4_1
X_14519_ systolic_inst.row_loop\[3\].col_loop\[3\].pe_i.prod_reg\[14\] _11698_ net118
+ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__mux2_1
XFILLER_147_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18287_ _05456_ _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__nand2_1
XFILLER_30_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15499_ _12551_ _12557_ VGND VGND VPWR VPWR _12558_ sky130_fd_sc_hd__nor2_1
XFILLER_175_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17238_ _04479_ _04481_ _04497_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__or3b_1
XFILLER_31_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_185_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17169_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[30\]
+ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__or2_1
XFILLER_157_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_181_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20180_ _07142_ _07144_ _07147_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__a21oi_2
XFILLER_89_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_181_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23870_ _11258_ systolic_inst.acc_wires\[0\]\[27\] net64 _10459_ VGND VGND VPWR VPWR
+ _01957_ sky130_fd_sc_hd__a22o_1
XFILLER_57_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22821_ _09500_ _09501_ _09502_ VGND VGND VPWR VPWR _09503_ sky130_fd_sc_hd__and3_1
XFILLER_38_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25540_ systolic_inst.acc_wires\[0\]\[16\] C_out\[16\] net54 VGND VGND VPWR VPWR
+ _02842_ sky130_fd_sc_hd__mux2_1
XFILLER_53_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22752_ _09433_ _09434_ _09428_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21703_ _08473_ _08477_ _08510_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_138_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25471_ systolic_inst.ce_local _11210_ VGND VGND VPWR VPWR _11211_ sky130_fd_sc_hd__and2_1
X_22683_ systolic_inst.B_outs\[0\]\[2\] systolic_inst.B_shift\[0\]\[2\] net121 VGND
+ VGND VPWR VPWR _01852_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27210_ clknet_leaf_246_clk _01008_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24422_ net114 ser_C.shift_reg\[39\] VGND VGND VPWR VPWR _10681_ sky130_fd_sc_hd__and2_1
X_21634_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[7\]
+ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__o21ai_2
X_28190_ clknet_leaf_130_clk _01988_ VGND VGND VPWR VPWR systolic_inst.B_shift\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27141_ clknet_leaf_6_clk _00939_ VGND VGND VPWR VPWR systolic_inst.A_shift\[21\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21565_ _08374_ _08375_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__nor2_1
X_24353_ C_out\[3\] net104 _10643_ ser_C.shift_reg\[3\] _10646_ VGND VGND VPWR VPWR
+ _02253_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_170_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23304_ _09932_ _09933_ VGND VGND VPWR VPWR _09934_ sky130_fd_sc_hd__and2b_1
X_20516_ _07396_ _07414_ _07413_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__o21a_1
XFILLER_138_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27072_ clknet_leaf_10_B_in_serial_clk _00870_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_24284_ _10615_ systolic_inst.B_shift\[23\]\[5\] net72 VGND VGND VPWR VPWR _02215_
+ sky130_fd_sc_hd__mux2_1
X_21496_ systolic_inst.A_outs\[3\]\[1\] systolic_inst.B_outs\[3\]\[2\] systolic_inst.B_outs\[3\]\[3\]
+ systolic_inst.A_outs\[3\]\[0\] VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__a22oi_1
XFILLER_14_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23235_ _09877_ _09879_ _09882_ _11713_ VGND VGND VPWR VPWR _09884_ sky130_fd_sc_hd__a31o_1
XFILLER_153_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26023_ systolic_inst.acc_wires\[15\]\[19\] ser_C.parallel_data\[499\] net23 VGND
+ VGND VPWR VPWR _03325_ sky130_fd_sc_hd__mux2_1
X_20447_ _07327_ _07345_ _07344_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__o21a_1
XFILLER_140_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23166_ _09817_ _09824_ VGND VGND VPWR VPWR _09825_ sky130_fd_sc_hd__nand2_1
Xclkload390 clknet_leaf_11_B_in_serial_clk VGND VGND VPWR VPWR clkload390/Y sky130_fd_sc_hd__bufinv_16
X_20378_ _07314_ _07315_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__nand2b_1
XFILLER_134_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22117_ _08861_ _08866_ VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__nand2_1
XFILLER_171_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27974_ clknet_leaf_174_clk _01772_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_23097_ _09765_ VGND VGND VPWR VPWR _09766_ sky130_fd_sc_hd__inv_2
XFILLER_216_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22048_ _08815_ _08819_ _08821_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__a21oi_1
X_26925_ clknet_leaf_5_A_in_serial_clk _00723_ net132 VGND VGND VPWR VPWR deser_A.serial_word\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29644_ clknet_leaf_32_B_in_serial_clk _03439_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26856_ clknet_leaf_0_B_in_serial_clk _00658_ net134 VGND VGND VPWR VPWR deser_B.bit_idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14870_ systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[6\] systolic_inst.A_outs\[14\]\[7\]
+ systolic_inst.B_outs\[14\]\[0\] VGND VGND VPWR VPWR _11993_ sky130_fd_sc_hd__a22o_1
X_13821_ net3 net126 deser_B.bit_idx\[0\] VGND VGND VPWR VPWR _11319_ sky130_fd_sc_hd__o21a_1
XFILLER_21_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25807_ systolic_inst.acc_wires\[8\]\[27\] C_out\[283\] net28 VGND VGND VPWR VPWR
+ _03109_ sky130_fd_sc_hd__mux2_1
XFILLER_235_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29575_ clknet_leaf_22_B_in_serial_clk _03370_ net137 VGND VGND VPWR VPWR deser_B.serial_word\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26787_ clknet_leaf_62_clk _00589_ net144 VGND VGND VPWR VPWR B_in\[59\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23999_ systolic_inst.B_shift\[9\]\[3\] B_in\[11\] _00008_ VGND VGND VPWR VPWR _10525_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28526_ clknet_leaf_161_clk _02324_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_16540_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[26\]
+ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__or2_1
XFILLER_56_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25738_ systolic_inst.acc_wires\[6\]\[22\] C_out\[214\] net46 VGND VGND VPWR VPWR
+ _03040_ sky130_fd_sc_hd__mux2_1
X_13752_ B_in\[59\] deser_B.word_buffer\[59\] net85 VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__mux2_1
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28457_ clknet_leaf_127_clk _02255_ net144 VGND VGND VPWR VPWR ser_C.shift_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_16471_ _03825_ _03828_ _03831_ net61 VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__a31o_1
XFILLER_232_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13683_ deser_B.word_buffer\[119\] deser_B.serial_word\[119\] net124 VGND VGND VPWR
+ VPWR _00520_ sky130_fd_sc_hd__mux2_1
X_25669_ systolic_inst.acc_wires\[4\]\[17\] C_out\[145\] net16 VGND VGND VPWR VPWR
+ _02971_ sky130_fd_sc_hd__mux2_1
XFILLER_43_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18210_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[9\]\[3\]
+ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15422_ _12463_ _12465_ _12464_ VGND VGND VPWR VPWR _12483_ sky130_fd_sc_hd__a21bo_1
X_27408_ clknet_leaf_227_clk _01206_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_203_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19190_ _06252_ _06253_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_1151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28388_ clknet_leaf_31_clk _02186_ VGND VGND VPWR VPWR systolic_inst.A_shift\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1064 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18141_ _05262_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__nand2_1
X_27339_ clknet_leaf_285_clk _01137_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_15353_ _12430_ _12434_ _12435_ VGND VGND VPWR VPWR _12436_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14304_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[6\] _11488_ VGND
+ VGND VPWR VPWR _11490_ sky130_fd_sc_hd__and3_1
X_18072_ _05191_ _05261_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__xnor2_4
XFILLER_172_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15284_ systolic_inst.acc_wires\[14\]\[16\] systolic_inst.acc_wires\[14\]\[17\] systolic_inst.acc_wires\[14\]\[18\]
+ systolic_inst.acc_wires\[14\]\[19\] systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _12378_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_93_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29009_ clknet_leaf_104_clk _02807_ net151 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_17023_ _04325_ _04326_ net69 VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_242_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_216_Left_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14235_ _11421_ _11422_ _11410_ VGND VGND VPWR VPWR _11423_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_242_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_242_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14166_ _11345_ _11355_ VGND VGND VPWR VPWR _11357_ sky130_fd_sc_hd__nand2_1
XFILLER_217_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13117_ systolic_inst.B_outs\[15\]\[7\] VGND VGND VPWR VPWR _11273_ sky130_fd_sc_hd__inv_2
X_14097_ deser_B.receiving deser_B.shift_reg\[1\] deser_B.shift_reg\[0\] _11305_ _11331_
+ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__a221o_1
X_18974_ net66 _06068_ _06069_ systolic_inst.acc_wires\[8\]\[25\] net108 VGND VGND
+ VPWR VPWR _01451_ sky130_fd_sc_hd__a32o_1
XFILLER_98_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_223_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew146 net147 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_16
XFILLER_112_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17925_ systolic_inst.B_outs\[9\]\[2\] systolic_inst.A_outs\[9\]\[5\] VGND VGND VPWR
+ VPWR _05119_ sky130_fd_sc_hd__nand2_1
XFILLER_65_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17856_ systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[4\] systolic_inst.A_outs\[9\]\[5\]
+ systolic_inst.B_outs\[9\]\[0\] VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__a22oi_1
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16807_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[9\] _04125_
+ _04126_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_236_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_225_Left_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_236_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17787_ systolic_inst.A_outs\[9\]\[2\] systolic_inst.A_outs\[8\]\[2\] net117 VGND
+ VGND VPWR VPWR _01332_ sky130_fd_sc_hd__mux2_1
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14999_ _12116_ _12117_ VGND VGND VPWR VPWR _12119_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19526_ _06563_ _06564_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__nand2_1
XFILLER_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16738_ _04058_ _04055_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__and2b_1
XFILLER_223_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19457_ _06501_ _06505_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16669_ _03991_ _03988_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__and2b_1
XFILLER_222_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18408_ systolic_inst.A_outs\[8\]\[5\] systolic_inst.A_shift\[16\]\[5\] net115 VGND
+ VGND VPWR VPWR _01399_ sky130_fd_sc_hd__mux2_1
X_19388_ _06446_ _06445_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__nand2b_1
XFILLER_50_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18339_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[9\]\[22\]
+ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__or2_1
XFILLER_72_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_187_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21350_ _08195_ _08200_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_234_Left_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20301_ _07234_ _07239_ _07240_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__and3_1
XFILLER_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21281_ _08141_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__inv_2
XFILLER_163_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23020_ _09694_ _09695_ VGND VGND VPWR VPWR _09696_ sky130_fd_sc_hd__nand2_1
X_20232_ systolic_inst.B_outs\[4\]\[1\] systolic_inst.B_outs\[0\]\[1\] net117 VGND
+ VGND VPWR VPWR _01595_ sky130_fd_sc_hd__mux2_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20163_ _07125_ _07126_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__nor2_1
XFILLER_103_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20094_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[6\]\[12\]
+ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__xnor2_1
X_24971_ C_out\[312\] net103 net76 ser_C.shift_reg\[312\] _10955_ VGND VGND VPWR VPWR
+ _02562_ sky130_fd_sc_hd__a221o_1
XFILLER_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26710_ clknet_leaf_10_B_in_serial_clk _00513_ net144 VGND VGND VPWR VPWR deser_B.word_buffer\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_23922_ systolic_inst.B_shift\[22\]\[5\] B_in\[85\] net59 VGND VGND VPWR VPWR _10494_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27690_ clknet_leaf_184_clk _01488_ net146 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26641_ clknet_leaf_14_B_in_serial_clk _00444_ net152 VGND VGND VPWR VPWR deser_B.word_buffer\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23853_ _10440_ _10442_ _10445_ VGND VGND VPWR VPWR _10446_ sky130_fd_sc_hd__a21oi_2
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22804_ _09478_ _09484_ VGND VGND VPWR VPWR _09486_ sky130_fd_sc_hd__xor2_1
XFILLER_84_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29360_ clknet_leaf_231_clk _03158_ net140 VGND VGND VPWR VPWR C_out\[332\] sky130_fd_sc_hd__dfrtp_1
X_26572_ clknet_leaf_23_A_in_serial_clk _00375_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_23784_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[0\]\[14\]
+ VGND VGND VPWR VPWR _10387_ sky130_fd_sc_hd__or2_1
X_20996_ _07828_ _07831_ _07869_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__o21a_1
XFILLER_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28311_ clknet_leaf_346_clk _02109_ VGND VGND VPWR VPWR systolic_inst.A_shift\[29\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25523_ _11244_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__inv_2
XFILLER_225_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22735_ _09418_ _09419_ _09401_ VGND VGND VPWR VPWR _09420_ sky130_fd_sc_hd__a21oi_1
XFILLER_197_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29291_ clknet_leaf_315_clk _03089_ net142 VGND VGND VPWR VPWR C_out\[263\] sky130_fd_sc_hd__dfrtp_1
XFILLER_198_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28242_ clknet_leaf_134_clk _02040_ VGND VGND VPWR VPWR systolic_inst.B_shift\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25454_ systolic_inst.ce_local _11199_ VGND VGND VPWR VPWR _11200_ sky130_fd_sc_hd__and2_1
XFILLER_13_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22666_ _09369_ _09372_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__nand2_1
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24405_ C_out\[29\] _11302_ net81 ser_C.shift_reg\[29\] _10672_ VGND VGND VPWR VPWR
+ _02279_ sky130_fd_sc_hd__a221o_1
X_28173_ clknet_leaf_78_clk _01971_ VGND VGND VPWR VPWR systolic_inst.B_shift\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21617_ _08390_ _08425_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__and2_1
XFILLER_181_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25385_ systolic_inst.A_shift\[3\]\[0\] A_in\[16\] net59 VGND VGND VPWR VPWR _11162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22597_ _09313_ _09314_ VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27124_ clknet_leaf_20_clk _00922_ VGND VGND VPWR VPWR systolic_inst.A_shift\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24336_ _10641_ systolic_inst.A_shift\[9\]\[7\] net70 VGND VGND VPWR VPWR _02241_
+ sky130_fd_sc_hd__mux2_1
X_21548_ _08354_ _08359_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__nand2b_1
XFILLER_217_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27055_ clknet_leaf_2_B_in_serial_clk _00853_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24267_ systolic_inst.B_shift\[17\]\[2\] net72 _11333_ B_in\[106\] VGND VGND VPWR
+ VPWR _02204_ sky130_fd_sc_hd__a22o_1
X_21479_ systolic_inst.B_outs\[2\]\[7\] systolic_inst.B_shift\[2\]\[7\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__mux2_1
XFILLER_153_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14020_ deser_B.shift_reg\[54\] deser_B.shift_reg\[55\] net125 VGND VGND VPWR VPWR
+ _00846_ sky130_fd_sc_hd__mux2_1
X_26006_ systolic_inst.acc_wires\[15\]\[2\] ser_C.parallel_data\[482\] net23 VGND
+ VGND VPWR VPWR _03308_ sky130_fd_sc_hd__mux2_1
X_23218_ _09860_ _09861_ VGND VGND VPWR VPWR _09869_ sky130_fd_sc_hd__nor2_1
XFILLER_181_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24198_ systolic_inst.B_shift\[22\]\[5\] net71 _11333_ B_in\[117\] VGND VGND VPWR
+ VPWR _02159_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_112_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23149_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[12\] systolic_inst.acc_wires\[1\]\[12\]
+ VGND VGND VPWR VPWR _09810_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27957_ clknet_leaf_169_clk _01755_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15971_ systolic_inst.B_outs\[11\]\[4\] systolic_inst.B_outs\[7\]\[4\] net119 VGND
+ VGND VPWR VPWR _01150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ _04937_ _04938_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__and2_1
X_14922_ _12042_ _12043_ VGND VGND VPWR VPWR _12044_ sky130_fd_sc_hd__nor2_1
X_26908_ clknet_leaf_17_A_in_serial_clk _00706_ net143 VGND VGND VPWR VPWR deser_A.serial_word\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18690_ _05806_ _05814_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_86_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27888_ clknet_leaf_309_clk _01686_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17641_ _04873_ _04879_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__nand2_1
X_29627_ clknet_leaf_9_B_in_serial_clk _03422_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_26839_ clknet_leaf_83_clk _00641_ net144 VGND VGND VPWR VPWR B_in\[111\] sky130_fd_sc_hd__dfrtp_1
X_14853_ _11974_ _11976_ VGND VGND VPWR VPWR _11977_ sky130_fd_sc_hd__nor2_1
XFILLER_236_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ B_in\[111\] deser_B.word_buffer\[111\] net88 VGND VGND VPWR VPWR _00641_
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29558_ clknet_leaf_16_B_in_serial_clk _03353_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_17572_ _04818_ _04821_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14784_ _11909_ _11910_ VGND VGND VPWR VPWR _11911_ sky130_fd_sc_hd__and2b_1
XFILLER_217_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_231_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19311_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[7\] _06346_ _06310_
+ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__a31o_1
X_28509_ clknet_leaf_111_clk _02307_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_231_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16523_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[12\]\[23\]
+ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_231_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13735_ B_in\[42\] deser_B.word_buffer\[42\] net84 VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__mux2_1
X_29489_ clknet_leaf_280_clk _03287_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[461\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19242_ _06277_ _06278_ _06279_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__o21ba_1
XFILLER_220_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16454_ net67 _03816_ _03818_ systolic_inst.acc_wires\[12\]\[12\] net108 VGND VGND
+ VPWR VPWR _01182_ sky130_fd_sc_hd__a32o_1
XFILLER_231_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13666_ deser_B.word_buffer\[102\] deser_B.serial_word\[102\] net123 VGND VGND VPWR
+ VPWR _00503_ sky130_fd_sc_hd__mux2_1
XFILLER_189_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15405_ _12463_ _12466_ VGND VGND VPWR VPWR _12467_ sky130_fd_sc_hd__xnor2_1
X_19173_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[7\]
+ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__o21ai_2
X_16385_ _03756_ _03758_ _03751_ _03754_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a211o_1
X_13597_ deser_B.word_buffer\[33\] deser_B.serial_word\[33\] net124 VGND VGND VPWR
+ VPWR _00434_ sky130_fd_sc_hd__mux2_1
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18124_ _05311_ _05312_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__nor2_1
XFILLER_200_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15336_ _12420_ _12421_ VGND VGND VPWR VPWR _12422_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_229_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_229_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18055_ _05188_ _05244_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__or2_1
XFILLER_144_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15267_ net107 systolic_inst.acc_wires\[14\]\[17\] _11712_ _12363_ VGND VGND VPWR
+ VPWR _01059_ sky130_fd_sc_hd__a22o_1
XANTENNA_2 _10501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17006_ net69 _04311_ _04313_ systolic_inst.acc_wires\[11\]\[5\] net105 VGND VGND
+ VPWR VPWR _01239_ sky130_fd_sc_hd__a32o_1
XFILLER_160_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14218_ systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[4\]
+ systolic_inst.A_outs\[15\]\[5\] VGND VGND VPWR VPWR _11406_ sky130_fd_sc_hd__and4_1
XFILLER_67_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15198_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[14\]\[8\]
+ VGND VGND VPWR VPWR _12304_ sky130_fd_sc_hd__nor2_1
XFILLER_99_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14149_ systolic_inst.B_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[2\] _11339_ _11340_
+ VGND VGND VPWR VPWR _11341_ sky130_fd_sc_hd__and4_1
XFILLER_67_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18957_ _06054_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__inv_2
XFILLER_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17908_ _05071_ _05074_ _05101_ _05102_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__a211oi_2
XFILLER_239_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18888_ _05989_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_176_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17839_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.B_outs\[9\]\[1\] systolic_inst.A_outs\[9\]\[3\]
+ systolic_inst.A_outs\[9\]\[4\] VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__and4_1
XFILLER_227_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20850_ systolic_inst.A_outs\[4\]\[0\] systolic_inst.A_outs\[4\]\[1\] systolic_inst.B_outs\[4\]\[1\]
+ systolic_inst.B_outs\[4\]\[2\] VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__and4_1
XFILLER_82_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19509_ _06546_ _06547_ _06541_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__or3b_1
X_20781_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[24\]
+ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__nor2_1
XFILLER_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22520_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[2\]\[8\]
+ VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__xor2_1
XFILLER_168_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22451_ _09189_ _09188_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__and2b_1
XFILLER_206_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21402_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[22\]
+ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__nand2_1
X_22382_ _08984_ _09122_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__or2_1
X_25170_ net110 ser_C.shift_reg\[413\] VGND VGND VPWR VPWR _11055_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_152_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21333_ _08182_ _08185_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__and2_1
X_24121_ systolic_inst.A_shift\[30\]\[0\] A_in\[112\] net59 VGND VGND VPWR VPWR _10562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24052_ _10543_ systolic_inst.B_shift\[0\]\[5\] _11332_ VGND VGND VPWR VPWR _02055_
+ sky130_fd_sc_hd__mux2_1
XFILLER_117_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21264_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[4\]\[2\]
+ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__or2_1
XFILLER_150_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23003_ _09676_ _09677_ VGND VGND VPWR VPWR _09680_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_165_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20215_ _07176_ _07177_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__nand2_1
XFILLER_116_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28860_ clknet_leaf_335_clk _02658_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[408\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21195_ _08061_ _08062_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__xor2_1
XFILLER_81_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27811_ clknet_leaf_140_clk _01609_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_20146_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[20\]
+ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_161_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28791_ clknet_leaf_201_clk _02589_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_104_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27742_ clknet_leaf_209_clk _01540_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_20077_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[6\]\[10\]
+ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__or2_1
X_24954_ net111 ser_C.shift_reg\[305\] VGND VGND VPWR VPWR _10947_ sky130_fd_sc_hd__and2_1
XFILLER_131_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23905_ _10485_ systolic_inst.B_shift\[13\]\[4\] net72 VGND VGND VPWR VPWR _01966_
+ sky130_fd_sc_hd__mux2_1
XFILLER_213_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27673_ clknet_leaf_142_clk _01471_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_73_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24885_ C_out\[269\] net101 net75 ser_C.shift_reg\[269\] _10912_ VGND VGND VPWR VPWR
+ _02519_ sky130_fd_sc_hd__a221o_1
X_29412_ clknet_leaf_327_clk _03210_ net136 VGND VGND VPWR VPWR C_out\[384\] sky130_fd_sc_hd__dfrtp_1
X_26624_ clknet_leaf_23_B_in_serial_clk _00427_ net143 VGND VGND VPWR VPWR deser_B.word_buffer\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_23836_ systolic_inst.acc_wires\[0\]\[20\] systolic_inst.acc_wires\[0\]\[21\] systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _10431_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_105_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29343_ clknet_leaf_223_clk _03141_ net149 VGND VGND VPWR VPWR C_out\[315\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_159_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26555_ clknet_leaf_27_A_in_serial_clk _00358_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[85\]
+ sky130_fd_sc_hd__dfrtp_1
X_23767_ _11258_ systolic_inst.acc_wires\[0\]\[11\] net63 _10372_ VGND VGND VPWR VPWR
+ _01941_ sky130_fd_sc_hd__a22o_1
XFILLER_54_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20979_ systolic_inst.A_outs\[4\]\[0\] _07852_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__nor2_1
XFILLER_198_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25506_ systolic_inst.cycle_cnt\[25\] _11279_ _11231_ VGND VGND VPWR VPWR _11234_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_207_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13520_ deser_A.shift_reg\[84\] deser_A.shift_reg\[85\] net129 VGND VGND VPWR VPWR
+ _00357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22718_ systolic_inst.B_outs\[1\]\[2\] systolic_inst.A_outs\[1\]\[2\] VGND VGND VPWR
+ VPWR _09403_ sky130_fd_sc_hd__and2_1
X_29274_ clknet_leaf_189_clk _03072_ net146 VGND VGND VPWR VPWR C_out\[246\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26486_ clknet_leaf_8_A_in_serial_clk _00289_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23698_ _10313_ VGND VGND VPWR VPWR _10314_ sky130_fd_sc_hd__inv_2
XFILLER_158_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28225_ clknet_leaf_98_clk _02023_ VGND VGND VPWR VPWR systolic_inst.B_shift\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25437_ systolic_inst.cycle_cnt\[1\] systolic_inst.cycle_cnt\[0\] _11306_ systolic_inst.cycle_cnt\[2\]
+ VGND VGND VPWR VPWR _11188_ sky130_fd_sc_hd__a31o_1
X_13451_ deser_A.shift_reg\[15\] deser_A.shift_reg\[16\] deser_A.receiving VGND VGND
+ VPWR VPWR _00288_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22649_ systolic_inst.acc_wires\[2\]\[26\] systolic_inst.acc_wires\[2\]\[27\] systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__o21a_1
XFILLER_186_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28156_ clknet_leaf_107_clk _01954_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16170_ net115 _03552_ _03553_ _03554_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__a31o_1
XFILLER_210_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25368_ ser_C.parallel_data\[511\] net98 net78 ser_C.shift_reg\[511\] VGND VGND VPWR
+ VPWR _02761_ sky130_fd_sc_hd__a22o_1
X_13382_ A_in\[91\] deser_A.word_buffer\[91\] net92 VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__mux2_1
XFILLER_194_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27107_ clknet_leaf_2_B_in_serial_clk _00905_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15121_ _12235_ _12236_ VGND VGND VPWR VPWR _12237_ sky130_fd_sc_hd__or2_1
XFILLER_177_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24319_ systolic_inst.A_shift\[11\]\[7\] A_in\[47\] net59 VGND VGND VPWR VPWR _10633_
+ sky130_fd_sc_hd__mux2_1
X_28087_ clknet_leaf_118_clk _01885_ net152 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_181_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25299_ ser_C.parallel_data\[476\] net102 net74 ser_C.shift_reg\[476\] _11119_ VGND
+ VGND VPWR VPWR _02726_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_75_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27038_ clknet_leaf_14_B_in_serial_clk _00836_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_15052_ _12134_ _12138_ _12169_ VGND VGND VPWR VPWR _12171_ sky130_fd_sc_hd__o21ai_1
XFILLER_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14003_ deser_B.shift_reg\[37\] deser_B.shift_reg\[38\] deser_B.receiving VGND VGND
+ VPWR VPWR _00829_ sky130_fd_sc_hd__mux2_1
XFILLER_181_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19860_ systolic_inst.A_outs\[6\]\[6\] _06858_ _06857_ VGND VGND VPWR VPWR _06859_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_134_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18811_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[8\]\[2\]
+ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__or2_1
X_19791_ _06790_ _06791_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28989_ clknet_leaf_57_clk _02787_ VGND VGND VPWR VPWR systolic_inst.A_shift\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15954_ net67 _12972_ _12973_ systolic_inst.acc_wires\[13\]\[30\] net107 VGND VGND
+ VPWR VPWR _01136_ sky130_fd_sc_hd__a32o_1
X_18742_ _05864_ _05865_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__and2_1
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14905_ _11963_ _11999_ _11997_ VGND VGND VPWR VPWR _12027_ sky130_fd_sc_hd__a21o_1
X_18673_ net108 _05797_ _05798_ _05799_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__o31ai_1
XFILLER_76_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_196_clk clknet_5_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_196_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15885_ _12895_ _12900_ _12905_ _12909_ VGND VGND VPWR VPWR _12915_ sky130_fd_sc_hd__or4_1
XFILLER_7_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14836_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[5\] _11959_
+ _11960_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__a22o_1
XFILLER_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17624_ _04862_ _04863_ _04864_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a21o_1
XFILLER_97_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17555_ _04741_ _04784_ _04783_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__o21a_1
X_14767_ _11887_ _11894_ VGND VGND VPWR VPWR _11895_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_28_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16506_ _03837_ _03840_ _03862_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__o21a_1
X_13718_ B_in\[25\] deser_B.word_buffer\[25\] net85 VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__mux2_1
XFILLER_232_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17486_ _04601_ _04738_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__or2_1
XFILLER_32_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14698_ net105 systolic_inst.acc_wires\[15\]\[24\] net69 _11851_ VGND VGND VPWR VPWR
+ _01002_ sky130_fd_sc_hd__a22o_1
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19225_ _06286_ _06287_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__xnor2_1
X_16437_ _03796_ _03798_ _03794_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__a21o_1
XFILLER_20_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13649_ deser_B.word_buffer\[85\] deser_B.serial_word\[85\] net124 VGND VGND VPWR
+ VPWR _00486_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19156_ _06184_ _06220_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__and2_1
X_16368_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[12\]\[1\]
+ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nand2_1
XFILLER_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_895 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18107_ systolic_inst.B_outs\[9\]\[5\] systolic_inst.A_outs\[9\]\[7\] VGND VGND VPWR
+ VPWR _05296_ sky130_fd_sc_hd__nand2_1
X_15319_ _11712_ _12406_ _12407_ systolic_inst.acc_wires\[14\]\[25\] net107 VGND VGND
+ VPWR VPWR _01067_ sky130_fd_sc_hd__a32o_1
X_19087_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[3\] _06151_ _06152_
+ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_120_clk clknet_5_28__leaf_clk VGND VGND VPWR VPWR clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_195_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16299_ _03590_ _03649_ _03648_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18038_ systolic_inst.A_outs\[9\]\[4\] systolic_inst.B_outs\[9\]\[6\] _11263_ systolic_inst.A_outs\[9\]\[3\]
+ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_A_in_serial_clk clknet_2_1__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_26_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_158_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20000_ _06992_ _06993_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19989_ _06958_ _06960_ _06983_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21951_ _08731_ _08733_ _08735_ _08738_ VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__o31ai_2
XFILLER_41_1258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_187_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_187_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_132_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _07751_ _07777_ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__or2_1
X_24670_ net110 ser_C.shift_reg\[163\] VGND VGND VPWR VPWR _10805_ sky130_fd_sc_hd__and2_1
XFILLER_82_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_195_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21882_ _08680_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__inv_2
X_23621_ _10228_ _10240_ VGND VGND VPWR VPWR _10242_ sky130_fd_sc_hd__nand2_1
XFILLER_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20833_ systolic_inst.A_outs\[4\]\[6\] systolic_inst.A_shift\[8\]\[6\] net121 VGND
+ VGND VPWR VPWR _01656_ sky130_fd_sc_hd__mux2_1
X_26340_ clknet_leaf_24_clk _00147_ net135 VGND VGND VPWR VPWR A_in\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_165_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23552_ _10109_ _10111_ _10172_ _10174_ VGND VGND VPWR VPWR _10175_ sky130_fd_sc_hd__a211oi_1
XFILLER_74_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_194_Right_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20764_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[22\]
+ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_154_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22503_ _09231_ _09232_ _09233_ VGND VGND VPWR VPWR _09235_ sky130_fd_sc_hd__and3_1
XFILLER_196_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26271_ clknet_leaf_22_A_in_serial_clk _00079_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_195_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20695_ net109 systolic_inst.acc_wires\[5\]\[11\] net64 _07612_ VGND VGND VPWR VPWR
+ _01629_ sky130_fd_sc_hd__a22o_1
X_23483_ systolic_inst.A_outs\[0\]\[4\] systolic_inst.B_outs\[0\]\[5\] _10025_ VGND
+ VGND VPWR VPWR _10107_ sky130_fd_sc_hd__a21oi_1
XFILLER_126_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28010_ clknet_leaf_167_clk _01808_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25222_ net110 ser_C.shift_reg\[439\] VGND VGND VPWR VPWR _11081_ sky130_fd_sc_hd__and2_1
X_22434_ _09142_ _09145_ _09173_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_150_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25153_ C_out\[403\] net101 net73 ser_C.shift_reg\[403\] _11046_ VGND VGND VPWR VPWR
+ _02653_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_111_clk clknet_5_29__leaf_clk VGND VGND VPWR VPWR clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
X_22365_ _09069_ _09071_ _09106_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__a21o_1
XFILLER_164_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24104_ _10561_ systolic_inst.B_shift\[19\]\[7\] net72 VGND VGND VPWR VPWR _02089_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21316_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[4\]\[10\]
+ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__nand2_1
X_22296_ _09001_ _09003_ _09038_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__nand3_1
XFILLER_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25084_ net113 ser_C.shift_reg\[370\] VGND VGND VPWR VPWR _11012_ sky130_fd_sc_hd__and2_1
XFILLER_102_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24035_ systolic_inst.B_shift\[8\]\[5\] B_in\[37\] _00008_ VGND VGND VPWR VPWR _10535_
+ sky130_fd_sc_hd__mux2_1
X_21247_ _08111_ _08112_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__xnor2_1
X_28912_ clknet_leaf_280_clk _02710_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[460\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21178_ _08030_ _08046_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__xor2_1
X_28843_ clknet_leaf_333_clk _02641_ net131 VGND VGND VPWR VPWR ser_C.shift_reg\[391\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20129_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[17\]
+ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__xor2_2
X_28774_ clknet_leaf_251_clk _02572_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[322\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25986_ systolic_inst.acc_wires\[14\]\[14\] ser_C.parallel_data\[462\] net26 VGND
+ VGND VPWR VPWR _03288_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27725_ clknet_leaf_215_clk _01523_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24937_ C_out\[295\] net102 net76 ser_C.shift_reg\[295\] _10938_ VGND VGND VPWR VPWR
+ _02545_ sky130_fd_sc_hd__a221o_1
XFILLER_92_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_178_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_178_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_133_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15670_ _12723_ _12722_ VGND VGND VPWR VPWR _12724_ sky130_fd_sc_hd__nand2b_1
XFILLER_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27656_ clknet_leaf_302_clk _01454_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24868_ net110 ser_C.shift_reg\[262\] VGND VGND VPWR VPWR _10904_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_103_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26607_ clknet_leaf_15_B_in_serial_clk _00410_ net151 VGND VGND VPWR VPWR deser_B.word_buffer\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14621_ _11781_ _11783_ _11785_ systolic_inst.acc_wires\[15\]\[13\] net105 VGND VGND
+ VPWR VPWR _00991_ sky130_fd_sc_hd__a32o_1
X_23819_ _10412_ _10414_ _10411_ VGND VGND VPWR VPWR _10417_ sky130_fd_sc_hd__o21ai_1
XFILLER_57_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27587_ clknet_leaf_216_clk _01385_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ C_out\[226\] net99 net79 ser_C.shift_reg\[226\] _10869_ VGND VGND VPWR VPWR
+ _02476_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17340_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[7\] _04597_ net118
+ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__mux2_1
X_29326_ clknet_leaf_221_clk _03124_ net139 VGND VGND VPWR VPWR C_out\[298\] sky130_fd_sc_hd__dfrtp_1
XFILLER_198_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14552_ net69 _11724_ _11726_ systolic_inst.acc_wires\[15\]\[3\] net107 VGND VGND
+ VPWR VPWR _00981_ sky130_fd_sc_hd__a32o_1
X_26538_ clknet_leaf_21_A_in_serial_clk _00341_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13503_ deser_A.shift_reg\[67\] deser_A.shift_reg\[68\] net129 VGND VGND VPWR VPWR
+ _00340_ sky130_fd_sc_hd__mux2_1
X_29257_ clknet_leaf_196_clk _03055_ net146 VGND VGND VPWR VPWR C_out\[229\] sky130_fd_sc_hd__dfrtp_1
X_17271_ _04491_ _04510_ _04509_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__a21bo_1
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26469_ clknet_leaf_346_clk deser_A.serial_toggle net132 VGND VGND VPWR VPWR deser_A.serial_toggle_sync1
+ sky130_fd_sc_hd__dfrtp_2
X_14483_ _11661_ _11662_ VGND VGND VPWR VPWR _11664_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_12_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19010_ _06099_ _06098_ systolic_inst.acc_wires\[8\]\[31\] net108 VGND VGND VPWR
+ VPWR _01457_ sky130_fd_sc_hd__a2bb2o_1
X_28208_ clknet_leaf_98_clk _02006_ VGND VGND VPWR VPWR systolic_inst.B_shift\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16222_ _03596_ _03604_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__nand2_1
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13434_ deser_A.bit_idx\[5\] _11316_ _11310_ _11282_ VGND VGND VPWR VPWR _00272_
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29188_ clknet_leaf_40_clk _02986_ net141 VGND VGND VPWR VPWR C_out\[160\] sky130_fd_sc_hd__dfrtp_1
Xclkload208 clknet_leaf_39_clk VGND VGND VPWR VPWR clkload208/X sky130_fd_sc_hd__clkbuf_4
X_28139_ clknet_leaf_125_clk _01937_ net144 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload219 clknet_leaf_52_clk VGND VGND VPWR VPWR clkload219/Y sky130_fd_sc_hd__inv_6
X_16153_ _03536_ _03537_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_102_clk clknet_5_23__leaf_clk VGND VGND VPWR VPWR clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13365_ A_in\[74\] deser_A.word_buffer\[74\] net94 VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__mux2_1
XFILLER_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15104_ _12176_ _12190_ _12188_ VGND VGND VPWR VPWR _12221_ sky130_fd_sc_hd__o21a_1
XFILLER_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16084_ _13077_ _13078_ _13047_ _13050_ VGND VGND VPWR VPWR _13080_ sky130_fd_sc_hd__o211a_1
XFILLER_138_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13296_ A_in\[5\] deser_A.word_buffer\[5\] net94 VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__mux2_1
XFILLER_54_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19912_ _06856_ _06874_ _06873_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__o21a_1
X_15035_ _12151_ _12152_ VGND VGND VPWR VPWR _12154_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19843_ _06802_ _06803_ _06805_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__o21a_1
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19774_ _06736_ _06739_ _06775_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_53_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_166_Left_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16986_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[11\]\[3\]
+ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__nand2_1
XFILLER_110_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18725_ _05849_ _05848_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__and2b_1
XFILLER_95_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_169_clk clknet_5_30__leaf_clk VGND VGND VPWR VPWR clknet_leaf_169_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15937_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[28\]
+ VGND VGND VPWR VPWR _12959_ sky130_fd_sc_hd__or2_1
XFILLER_225_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15868_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[16\]
+ _12897_ VGND VGND VPWR VPWR _12901_ sky130_fd_sc_hd__a21oi_1
X_18656_ _05781_ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__nand2b_1
XFILLER_97_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14819_ systolic_inst.A_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[2\] systolic_inst.B_outs\[14\]\[3\]
+ systolic_inst.B_outs\[14\]\[4\] VGND VGND VPWR VPWR _11944_ sky130_fd_sc_hd__and4_1
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17607_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[10\]\[5\]
+ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__or2_1
XFILLER_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15799_ _12838_ _12839_ _12840_ VGND VGND VPWR VPWR _12842_ sky130_fd_sc_hd__nand3_1
X_18587_ _05713_ _05714_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__xor2_1
XFILLER_75_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17538_ _04740_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_190_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17469_ _04714_ _04722_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__nand2_1
XFILLER_177_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_341_clk clknet_5_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_341_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_225_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_175_Left_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19208_ _06235_ _06241_ _06240_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__a21o_1
X_20480_ _07396_ _07414_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__xor2_1
XFILLER_203_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19139_ _06204_ _06200_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__nand2b_1
XFILLER_192_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22150_ systolic_inst.A_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[2\] systolic_inst.B_outs\[2\]\[3\]
+ systolic_inst.B_outs\[2\]\[4\] VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__and4_1
XFILLER_106_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21101_ _07926_ _07934_ _07933_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__a21o_1
XFILLER_218_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22081_ systolic_inst.A_outs\[2\]\[3\] systolic_inst.A_outs\[1\]\[3\] net122 VGND
+ VGND VPWR VPWR _01781_ sky130_fd_sc_hd__mux2_1
XFILLER_236_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21032_ _07904_ _07872_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_5_28__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_5_28__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_236_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_184_Left_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25840_ systolic_inst.acc_wires\[9\]\[28\] C_out\[316\] net13 VGND VGND VPWR VPWR
+ _03142_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25771_ systolic_inst.acc_wires\[7\]\[23\] C_out\[247\] net44 VGND VGND VPWR VPWR
+ _03073_ sky130_fd_sc_hd__mux2_1
XFILLER_80_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22983_ systolic_inst.B_outs\[1\]\[5\] systolic_inst.A_outs\[1\]\[7\] VGND VGND VPWR
+ VPWR _09660_ sky130_fd_sc_hd__nand2_1
XFILLER_41_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27510_ clknet_leaf_231_clk _01308_ net140 VGND VGND VPWR VPWR systolic_inst.acc_wires\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24722_ net113 ser_C.shift_reg\[189\] VGND VGND VPWR VPWR _10831_ sky130_fd_sc_hd__and2_1
XFILLER_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28490_ clknet_leaf_116_clk _02288_ net152 VGND VGND VPWR VPWR ser_C.shift_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_21934_ net68 _08723_ _08724_ systolic_inst.acc_wires\[3\]\[10\] net106 VGND VGND
+ VPWR VPWR _01756_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_156_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27441_ clknet_leaf_249_clk _01239_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24653_ C_out\[153\] net104 _10643_ ser_C.shift_reg\[153\] _10796_ VGND VGND VPWR
+ VPWR _02403_ sky130_fd_sc_hd__a221o_1
XFILLER_231_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21865_ net122 _08656_ _08666_ VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__and3_1
XFILLER_242_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23604_ _10221_ _10223_ VGND VGND VPWR VPWR _10225_ sky130_fd_sc_hd__xnor2_1
X_20816_ _07705_ _07708_ _07711_ _07714_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__o31a_1
X_27372_ clknet_leaf_327_clk _01170_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24584_ net114 ser_C.shift_reg\[120\] VGND VGND VPWR VPWR _10762_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_193_Left_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21796_ _08553_ _08569_ _08567_ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__o21a_1
X_29111_ clknet_leaf_154_clk _02909_ net150 VGND VGND VPWR VPWR C_out\[83\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26323_ clknet_leaf_29_A_in_serial_clk _00131_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_23535_ _10156_ _10157_ VGND VGND VPWR VPWR _10158_ sky130_fd_sc_hd__or2_1
XFILLER_168_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20747_ _07652_ _07654_ _07651_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_332_clk clknet_5_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_332_clk
+ sky130_fd_sc_hd__clkbuf_8
X_29042_ clknet_leaf_99_clk _02840_ net152 VGND VGND VPWR VPWR C_out\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_196_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26254_ clknet_leaf_3_A_in_serial_clk _00062_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23466_ _10072_ _10089_ _10090_ VGND VGND VPWR VPWR _10091_ sky130_fd_sc_hd__and3_1
XFILLER_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20678_ _07593_ _07595_ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__nand2_1
X_25205_ C_out\[429\] net101 net73 ser_C.shift_reg\[429\] _11072_ VGND VGND VPWR VPWR
+ _02679_ sky130_fd_sc_hd__a221o_1
XFILLER_52_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22417_ _09130_ _09156_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__nand2b_1
X_26185_ ser_C.bit_idx\[5\] _11250_ VGND VGND VPWR VPWR _11252_ sky130_fd_sc_hd__and2_1
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23397_ _11258_ _10021_ _10022_ _10023_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__o31ai_1
X_13150_ net7 net10 VGND VGND VPWR VPWR _11302_ sky130_fd_sc_hd__and2b_4
XFILLER_124_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25136_ net110 ser_C.shift_reg\[396\] VGND VGND VPWR VPWR _11038_ sky130_fd_sc_hd__and2_1
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22348_ systolic_inst.A_outs\[2\]\[6\] _09060_ _09061_ _09025_ VGND VGND VPWR VPWR
+ _09090_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_192_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25067_ C_out\[360\] net97 net77 ser_C.shift_reg\[360\] _11003_ VGND VGND VPWR VPWR
+ _02610_ sky130_fd_sc_hd__a221o_1
X_22279_ _08985_ _09021_ VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__and2_1
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24018_ systolic_inst.B_shift\[6\]\[1\] _11332_ net83 systolic_inst.B_shift\[10\]\[1\]
+ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__a22o_1
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28826_ clknet_leaf_238_clk _02624_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[374\]
+ sky130_fd_sc_hd__dfrtp_1
X_16840_ _04086_ _04121_ _04122_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_6_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_230_Right_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16771_ net119 _04089_ _04090_ _04091_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__a31o_1
XFILLER_92_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13983_ deser_B.shift_reg\[17\] deser_B.shift_reg\[18\] net125 VGND VGND VPWR VPWR
+ _00809_ sky130_fd_sc_hd__mux2_1
X_28757_ clknet_leaf_223_clk _02555_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[305\]
+ sky130_fd_sc_hd__dfrtp_1
X_25969_ systolic_inst.acc_wires\[13\]\[29\] ser_C.parallel_data\[445\] net26 VGND
+ VGND VPWR VPWR _03271_ sky130_fd_sc_hd__mux2_1
XFILLER_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15722_ systolic_inst.B_outs\[13\]\[5\] systolic_inst.B_outs\[13\]\[6\] systolic_inst.A_outs\[13\]\[7\]
+ _12773_ VGND VGND VPWR VPWR _12774_ sky130_fd_sc_hd__a31o_1
X_18510_ _05635_ _05636_ _05640_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__nand3_2
X_27708_ clknet_leaf_192_clk _01506_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_185_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19490_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[7\]\[13\]
+ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__xor2_1
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28688_ clknet_leaf_192_clk _02486_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[236\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15653_ _12667_ _12669_ _12706_ VGND VGND VPWR VPWR _12708_ sky130_fd_sc_hd__a21o_1
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18441_ _05573_ _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__and2_1
XFILLER_59_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27639_ clknet_leaf_316_clk _01437_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14604_ _11769_ _11770_ VGND VGND VPWR VPWR _11771_ sky130_fd_sc_hd__xnor2_1
X_18372_ net105 systolic_inst.acc_wires\[9\]\[26\] net66 _05530_ VGND VGND VPWR VPWR
+ _01388_ sky130_fd_sc_hd__a22o_1
XFILLER_57_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _12605_ _12608_ _12640_ VGND VGND VPWR VPWR _12641_ sky130_fd_sc_hd__o21ai_1
XFILLER_226_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17323_ _04577_ _04580_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14535_ net106 systolic_inst.load_acc VGND VGND VPWR VPWR _11712_ sky130_fd_sc_hd__nor2_8
XFILLER_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29309_ clknet_leaf_313_clk _03107_ net141 VGND VGND VPWR VPWR C_out\[281\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_323_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_323_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_222_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17254_ systolic_inst.A_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[2\] systolic_inst.B_outs\[10\]\[3\]
+ systolic_inst.B_outs\[10\]\[4\] VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__nand4_1
X_14466_ _11645_ _11646_ VGND VGND VPWR VPWR _11648_ sky130_fd_sc_hd__nor2_1
XFILLER_175_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16205_ net115 _03586_ _03587_ _03588_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__a31o_1
XFILLER_179_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13417_ A_in\[126\] deser_A.word_buffer\[126\] net92 VGND VGND VPWR VPWR _00265_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17185_ systolic_inst.A_outs\[10\]\[7\] systolic_inst.A_outs\[9\]\[7\] net120 VGND
+ VGND VPWR VPWR _01273_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14397_ _11541_ _11544_ _11579_ VGND VGND VPWR VPWR _11581_ sky130_fd_sc_hd__and3_1
XFILLER_122_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16136_ _03514_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__xnor2_1
X_13348_ A_in\[57\] deser_A.word_buffer\[57\] net91 VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__mux2_1
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16067_ systolic_inst.B_outs\[12\]\[2\] systolic_inst.A_outs\[12\]\[4\] VGND VGND
+ VPWR VPWR _13063_ sky130_fd_sc_hd__nand2_1
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13279_ deser_A.word_buffer\[117\] deser_A.serial_word\[117\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15018_ _12062_ _12066_ _12100_ _12135_ _12098_ VGND VGND VPWR VPWR _12138_ sky130_fd_sc_hd__o311a_1
XFILLER_130_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19826_ systolic_inst.B_outs\[6\]\[4\] systolic_inst.A_outs\[6\]\[5\] systolic_inst.A_outs\[6\]\[6\]
+ systolic_inst.B_outs\[6\]\[3\] VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__a22oi_1
XFILLER_116_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_200_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19757_ systolic_inst.A_outs\[6\]\[1\] systolic_inst.B_outs\[6\]\[6\] _06758_ VGND
+ VGND VPWR VPWR _06759_ sky130_fd_sc_hd__and3_1
XFILLER_96_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16969_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[11\]\[0\]
+ systolic_inst.load_acc VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__a21o_1
XFILLER_37_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18708_ _05694_ _05832_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__or2_1
XFILLER_225_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19688_ _06670_ _06690_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_192_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18639_ _05764_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__or2_1
XFILLER_224_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21650_ _08458_ _08457_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__nand2b_1
XFILLER_40_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20601_ _07464_ _07507_ _07506_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__o21a_1
XFILLER_220_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21581_ _08360_ _08391_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_314_clk clknet_5_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_314_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_178_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23320_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.B_outs\[0\]\[2\] systolic_inst.A_outs\[0\]\[2\]
+ systolic_inst.A_outs\[0\]\[3\] VGND VGND VPWR VPWR _09949_ sky130_fd_sc_hd__nand4_2
X_20532_ _07464_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__inv_2
XFILLER_138_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23251_ net109 systolic_inst.acc_wires\[1\]\[27\] net65 _09896_ VGND VGND VPWR VPWR
+ _01901_ sky130_fd_sc_hd__a22o_1
X_20463_ systolic_inst.B_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[7\]
+ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__and3_1
XFILLER_203_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22202_ systolic_inst.B_outs\[2\]\[1\] systolic_inst.A_outs\[2\]\[6\] systolic_inst.A_outs\[2\]\[7\]
+ systolic_inst.B_outs\[2\]\[0\] VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__a22o_1
X_23182_ _11713_ _09838_ VGND VGND VPWR VPWR _09839_ sky130_fd_sc_hd__nor2_1
X_20394_ _07287_ _07330_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__xnor2_1
X_22133_ _08880_ _08881_ _08862_ VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__o21ai_1
X_27990_ clknet_leaf_121_clk _01788_ net152 VGND VGND VPWR VPWR systolic_inst.B_outs\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_160_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26941_ clknet_leaf_19_A_in_serial_clk _00739_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_22064_ _08834_ _08835_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__nor2_1
XFILLER_82_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21015_ systolic_inst.A_outs\[4\]\[2\] systolic_inst.B_outs\[4\]\[6\] VGND VGND VPWR
+ VPWR _07888_ sky130_fd_sc_hd__nand2_1
X_29660_ clknet_leaf_8_B_in_serial_clk _03455_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_26872_ clknet_leaf_15_A_in_serial_clk _00670_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28611_ clknet_leaf_137_clk _02409_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[159\]
+ sky130_fd_sc_hd__dfrtp_1
X_25823_ systolic_inst.acc_wires\[9\]\[11\] C_out\[299\] net15 VGND VGND VPWR VPWR
+ _03125_ sky130_fd_sc_hd__mux2_1
X_29591_ clknet_leaf_12_B_in_serial_clk _03386_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_229_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28542_ clknet_leaf_163_clk _02340_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_25754_ systolic_inst.acc_wires\[7\]\[6\] C_out\[230\] net40 VGND VGND VPWR VPWR
+ _03056_ sky130_fd_sc_hd__mux2_1
X_22966_ _09641_ _09642_ VGND VGND VPWR VPWR _09644_ sky130_fd_sc_hd__and2b_1
XFILLER_228_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24705_ C_out\[179\] net99 net79 ser_C.shift_reg\[179\] _10822_ VGND VGND VPWR VPWR
+ _02429_ sky130_fd_sc_hd__a221o_1
X_28473_ clknet_leaf_102_clk _02271_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_21917_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[3\]\[8\]
+ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_28_B_in_serial_clk clknet_2_0__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_28_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_25685_ systolic_inst.acc_wires\[5\]\[1\] C_out\[161\] net16 VGND VGND VPWR VPWR
+ _02987_ sky130_fd_sc_hd__mux2_1
XFILLER_82_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22897_ _09576_ _09575_ VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__nand2b_1
XFILLER_70_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27424_ clknet_leaf_248_clk _01222_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24636_ net7 ser_C.shift_reg\[146\] VGND VGND VPWR VPWR _10788_ sky130_fd_sc_hd__and2_1
X_21848_ _08650_ _08649_ VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_175_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27355_ clknet_leaf_231_clk _01153_ net140 VGND VGND VPWR VPWR systolic_inst.B_outs\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_24567_ C_out\[110\] net100 net80 ser_C.shift_reg\[110\] _10753_ VGND VGND VPWR VPWR
+ _02360_ sky130_fd_sc_hd__a221o_1
XFILLER_54_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_305_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_305_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21779_ _08442_ _08582_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__nand2_2
XFILLER_169_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14320_ _11474_ _11504_ VGND VGND VPWR VPWR _11506_ sky130_fd_sc_hd__xnor2_1
X_26306_ clknet_leaf_25_A_in_serial_clk _00114_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_23518_ _10140_ _10141_ VGND VGND VPWR VPWR _10142_ sky130_fd_sc_hd__and2_1
XFILLER_19_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27286_ clknet_leaf_320_clk _01084_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_24498_ net113 ser_C.shift_reg\[77\] VGND VGND VPWR VPWR _10719_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_134_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29025_ clknet_leaf_92_clk _02823_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_134_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14251_ systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[5\] systolic_inst.A_outs\[15\]\[6\]
+ systolic_inst.B_outs\[15\]\[1\] VGND VGND VPWR VPWR _11438_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26237_ clknet_leaf_16_A_in_serial_clk _00045_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_23449_ systolic_inst.B_outs\[0\]\[3\] systolic_inst.B_outs\[0\]\[4\] systolic_inst.A_outs\[0\]\[4\]
+ systolic_inst.A_outs\[0\]\[5\] VGND VGND VPWR VPWR _10074_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_59_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ deser_A.word_buffer\[40\] deser_A.serial_word\[40\] net127 VGND VGND VPWR
+ VPWR _00050_ sky130_fd_sc_hd__mux2_1
XFILLER_165_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26168_ deser_B.serial_word\[123\] deser_B.shift_reg\[123\] net56 VGND VGND VPWR
+ VPWR _03470_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14182_ _11340_ _11348_ _11349_ _11352_ VGND VGND VPWR VPWR _11372_ sky130_fd_sc_hd__o22ai_2
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13133_ systolic_inst.cycle_cnt\[23\] systolic_inst.cycle_cnt\[22\] systolic_inst.cycle_cnt\[21\]
+ systolic_inst.cycle_cnt\[20\] VGND VGND VPWR VPWR _11286_ sky130_fd_sc_hd__or4_1
X_25119_ C_out\[386\] net101 net73 ser_C.shift_reg\[386\] _11029_ VGND VGND VPWR VPWR
+ _02636_ sky130_fd_sc_hd__a221o_1
XFILLER_48_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26099_ deser_B.serial_word\[54\] deser_B.shift_reg\[54\] net56 VGND VGND VPWR VPWR
+ _03401_ sky130_fd_sc_hd__mux2_1
XFILLER_139_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18990_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[28\]
+ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__nand2_1
XFILLER_87_1088 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_240_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_240_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17941_ _05118_ _05134_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_11__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_11__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_17872_ _05067_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__inv_2
XFILLER_152_1356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19611_ _06636_ _06635_ systolic_inst.acc_wires\[7\]\[31\] net105 VGND VGND VPWR
+ VPWR _01521_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_128_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28809_ clknet_leaf_244_clk _02607_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[357\]
+ sky130_fd_sc_hd__dfrtp_1
X_16823_ _04139_ _04140_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19542_ _06576_ _06577_ _06574_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__o21ai_2
XFILLER_150_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13966_ deser_A.serial_word\[127\] deser_A.shift_reg\[127\] _00002_ VGND VGND VPWR
+ VPWR _00792_ sky130_fd_sc_hd__mux2_1
X_16754_ _04066_ _04074_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_238_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_238_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15705_ _12756_ _12757_ VGND VGND VPWR VPWR _12758_ sky130_fd_sc_hd__nand2b_1
XFILLER_228_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19473_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[7\]\[11\]
+ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__nor2_1
X_16685_ _04005_ _04006_ _03994_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__o21bai_1
XFILLER_111_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13897_ deser_A.serial_word\[58\] deser_A.shift_reg\[58\] _00002_ VGND VGND VPWR
+ VPWR _00723_ sky130_fd_sc_hd__mux2_1
XFILLER_235_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18424_ _05559_ _05557_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[1\]
+ net108 VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_234_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15636_ _12689_ _12690_ VGND VGND VPWR VPWR _12691_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_234_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18355_ _05495_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__nor2_1
X_15567_ _12622_ _12623_ VGND VGND VPWR VPWR _12624_ sky130_fd_sc_hd__nor2_1
XFILLER_226_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _11695_ _11697_ VGND VGND VPWR VPWR _11698_ sky130_fd_sc_hd__xnor2_1
X_17306_ systolic_inst.B_outs\[10\]\[1\] systolic_inst.A_outs\[10\]\[6\] systolic_inst.A_outs\[10\]\[7\]
+ systolic_inst.B_outs\[10\]\[0\] VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__a22o_1
XFILLER_222_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15498_ _12521_ _12556_ VGND VGND VPWR VPWR _12557_ sky130_fd_sc_hd__xnor2_1
X_18286_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[9\]\[14\]
+ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__nand2_1
XFILLER_175_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14449_ _11593_ _11630_ VGND VGND VPWR VPWR _11631_ sky130_fd_sc_hd__xnor2_1
X_17237_ _04479_ _04481_ _04497_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_185_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_185_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17168_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[11\]\[30\]
+ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__nand2_1
XFILLER_196_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_185_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16119_ _03502_ _03503_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_181_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17099_ _04391_ _04392_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_181_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19809_ _06809_ _06779_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__nand2b_1
XFILLER_131_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22820_ _09466_ _09468_ VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_179_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22751_ _09428_ _09433_ _09434_ VGND VGND VPWR VPWR _09435_ sky130_fd_sc_hd__and3_1
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_91_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
X_21702_ _08507_ _08508_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25470_ systolic_inst.cycle_cnt\[13\] systolic_inst.cycle_cnt\[12\] _11206_ VGND
+ VGND VPWR VPWR _11210_ sky130_fd_sc_hd__and3_1
XFILLER_240_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22682_ systolic_inst.B_outs\[0\]\[1\] systolic_inst.B_shift\[0\]\[1\] net121 VGND
+ VGND VPWR VPWR _01851_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24421_ C_out\[37\] _11302_ net81 ser_C.shift_reg\[37\] _10680_ VGND VGND VPWR VPWR
+ _02287_ sky130_fd_sc_hd__a221o_1
XFILLER_80_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21633_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[7\]
+ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__o21a_1
XFILLER_240_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27140_ clknet_leaf_6_clk _00938_ VGND VGND VPWR VPWR systolic_inst.A_shift\[21\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24352_ net7 ser_C.shift_reg\[4\] VGND VGND VPWR VPWR _10646_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_170_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21564_ systolic_inst.B_outs\[3\]\[0\] systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[5\]
+ systolic_inst.A_outs\[3\]\[6\] VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_170_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23303_ _09930_ _09931_ _09923_ VGND VGND VPWR VPWR _09933_ sky130_fd_sc_hd__a21bo_1
X_27071_ clknet_leaf_10_B_in_serial_clk _00869_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_193_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20515_ _07432_ _07448_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__xor2_1
XFILLER_176_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24283_ systolic_inst.B_shift\[27\]\[5\] B_in\[93\] _00008_ VGND VGND VPWR VPWR _10615_
+ sky130_fd_sc_hd__mux2_1
X_21495_ net106 systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[2\] _08308_
+ _08309_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__a22o_1
XFILLER_166_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26022_ systolic_inst.acc_wires\[15\]\[18\] ser_C.parallel_data\[498\] net23 VGND
+ VGND VPWR VPWR _03324_ sky130_fd_sc_hd__mux2_1
X_23234_ _09877_ _09879_ _09882_ VGND VGND VPWR VPWR _09883_ sky130_fd_sc_hd__a21oi_2
XFILLER_140_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20446_ _07380_ _07381_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__and2_1
XFILLER_181_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23165_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[1\]\[13\]
+ _09818_ VGND VGND VPWR VPWR _09824_ sky130_fd_sc_hd__a21oi_1
Xclkload380 clknet_leaf_21_B_in_serial_clk VGND VGND VPWR VPWR clkload380/Y sky130_fd_sc_hd__clkinv_2
XFILLER_162_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20377_ _07312_ _07313_ _07277_ _07279_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__o211ai_1
Xclkload391 clknet_leaf_12_B_in_serial_clk VGND VGND VPWR VPWR clkload391/Y sky130_fd_sc_hd__bufinv_16
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22116_ _08864_ _08865_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__and2_1
XFILLER_136_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27973_ clknet_leaf_174_clk _01771_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_23096_ _09761_ _09762_ _09763_ VGND VGND VPWR VPWR _09765_ sky130_fd_sc_hd__and3_1
XFILLER_161_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22047_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[27\]
+ VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__xnor2_1
X_26924_ clknet_leaf_6_A_in_serial_clk _00722_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_212_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29643_ clknet_leaf_31_B_in_serial_clk _03438_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26855_ clknet_leaf_70_clk _00657_ net135 VGND VGND VPWR VPWR B_in\[127\] sky130_fd_sc_hd__dfrtp_1
XFILLER_76_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13820_ B_in\[127\] deser_B.word_buffer\[127\] net89 VGND VGND VPWR VPWR _00657_
+ sky130_fd_sc_hd__mux2_1
X_25806_ systolic_inst.acc_wires\[8\]\[26\] C_out\[282\] net28 VGND VGND VPWR VPWR
+ _03108_ sky130_fd_sc_hd__mux2_1
X_29574_ clknet_leaf_22_B_in_serial_clk _03369_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_26786_ clknet_leaf_63_clk _00588_ net144 VGND VGND VPWR VPWR B_in\[58\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23998_ _10524_ systolic_inst.B_shift\[5\]\[2\] _11332_ VGND VGND VPWR VPWR _02020_
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28525_ clknet_leaf_161_clk _02323_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_25737_ systolic_inst.acc_wires\[6\]\[21\] C_out\[213\] net46 VGND VGND VPWR VPWR
+ _03039_ sky130_fd_sc_hd__mux2_1
X_13751_ B_in\[58\] deser_B.word_buffer\[58\] net89 VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__mux2_1
XFILLER_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22949_ _09557_ _09626_ VGND VGND VPWR VPWR _09627_ sky130_fd_sc_hd__xnor2_4
XFILLER_21_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_82_clk clknet_5_21__leaf_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_84_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16470_ _03825_ _03828_ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__a21oi_1
X_28456_ clknet_leaf_126_clk _02254_ net144 VGND VGND VPWR VPWR ser_C.shift_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13682_ deser_B.word_buffer\[118\] deser_B.serial_word\[118\] net124 VGND VGND VPWR
+ VPWR _00519_ sky130_fd_sc_hd__mux2_1
X_25668_ systolic_inst.acc_wires\[4\]\[16\] C_out\[144\] net30 VGND VGND VPWR VPWR
+ _02970_ sky130_fd_sc_hd__mux2_1
X_15421_ _12471_ _12474_ VGND VGND VPWR VPWR _12482_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_80_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27407_ clknet_leaf_227_clk _01205_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_24619_ C_out\[136\] net103 net75 ser_C.shift_reg\[136\] _10779_ VGND VGND VPWR VPWR
+ _02386_ sky130_fd_sc_hd__a221o_1
X_28387_ clknet_leaf_31_clk _02185_ VGND VGND VPWR VPWR systolic_inst.A_shift\[18\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25599_ systolic_inst.acc_wires\[2\]\[11\] C_out\[75\] net51 VGND VGND VPWR VPWR
+ _02901_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27338_ clknet_leaf_285_clk _01136_ net136 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_15352_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[31\]
+ VGND VGND VPWR VPWR _12435_ sky130_fd_sc_hd__xnor2_1
X_18140_ _05325_ _05326_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__xnor2_1
XFILLER_223_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14303_ systolic_inst.A_outs\[15\]\[2\] systolic_inst.B_outs\[15\]\[6\] VGND VGND
+ VPWR VPWR _11489_ sky130_fd_sc_hd__nand2_1
XFILLER_200_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18071_ _05224_ _05260_ systolic_inst.A_outs\[9\]\[7\] VGND VGND VPWR VPWR _05261_
+ sky130_fd_sc_hd__and3b_1
XFILLER_157_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15283_ _12355_ _12376_ VGND VGND VPWR VPWR _12377_ sky130_fd_sc_hd__nor2_1
X_27269_ clknet_leaf_268_clk _01067_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17022_ _04325_ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__and2_1
X_29008_ clknet_leaf_104_clk _02806_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14234_ _11419_ _11420_ _11392_ VGND VGND VPWR VPWR _11422_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_242_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_242_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14165_ _11345_ _11355_ VGND VGND VPWR VPWR _11356_ sky130_fd_sc_hd__or2_1
XFILLER_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13116_ systolic_inst.B_outs\[13\]\[7\] VGND VGND VPWR VPWR _11272_ sky130_fd_sc_hd__inv_2
XFILLER_154_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14096_ net126 net4 net3 VGND VGND VPWR VPWR _11331_ sky130_fd_sc_hd__and3b_1
XFILLER_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18973_ _06063_ _06065_ _06067_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew136 net137 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_16
X_17924_ _05081_ _05117_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__xnor2_1
XFILLER_230_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17855_ _05029_ _05031_ _05030_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a21bo_1
X_16806_ _04086_ _04089_ _04124_ net105 VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__a31oi_1
XFILLER_94_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_236_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17786_ systolic_inst.A_outs\[9\]\[1\] systolic_inst.A_outs\[8\]\[1\] net117 VGND
+ VGND VPWR VPWR _01331_ sky130_fd_sc_hd__mux2_1
XFILLER_208_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14998_ _12117_ _12116_ VGND VGND VPWR VPWR _12118_ sky130_fd_sc_hd__nand2b_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19525_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[18\]
+ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__nand2_1
X_16737_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] _04057_ VGND
+ VGND VPWR VPWR _04058_ sky130_fd_sc_hd__a21o_1
X_13949_ deser_A.serial_word\[110\] deser_A.shift_reg\[110\] net57 VGND VGND VPWR
+ VPWR _00775_ sky130_fd_sc_hd__mux2_1
XFILLER_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_clk clknet_5_20__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19456_ _06503_ _06504_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__nor2_1
X_16668_ _03989_ _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__or2_1
XFILLER_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18407_ systolic_inst.A_outs\[8\]\[4\] systolic_inst.A_shift\[16\]\[4\] net115 VGND
+ VGND VPWR VPWR _01398_ sky130_fd_sc_hd__mux2_1
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15619_ _12605_ _12638_ _12639_ VGND VGND VPWR VPWR _12675_ sky130_fd_sc_hd__a21o_1
XFILLER_241_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19387_ _06374_ _06422_ _06421_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16599_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[1\]
+ systolic_inst.A_outs\[11\]\[2\] VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__and4_1
XFILLER_163_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18338_ _05501_ _05500_ systolic_inst.acc_wires\[9\]\[21\] net106 VGND VGND VPWR
+ VPWR _01383_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_187_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18269_ _05419_ _05423_ _05424_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__o21ai_1
X_20300_ _07237_ _07238_ _07236_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__o21ai_1
XFILLER_135_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21280_ _08131_ _08135_ _08138_ _08139_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__o211a_1
X_20231_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.B_outs\[0\]\[0\] net117 VGND
+ VGND VPWR VPWR _01594_ sky130_fd_sc_hd__mux2_1
XFILLER_116_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20162_ systolic_inst.acc_wires\[6\]\[20\] systolic_inst.acc_wires\[6\]\[21\] systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__o21a_1
XFILLER_171_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20093_ _07059_ _07065_ _07067_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__o21a_1
X_24970_ net111 ser_C.shift_reg\[313\] VGND VGND VPWR VPWR _10955_ sky130_fd_sc_hd__and2_1
XFILLER_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_163_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23921_ _10493_ systolic_inst.B_shift\[18\]\[4\] net71 VGND VGND VPWR VPWR _01974_
+ sky130_fd_sc_hd__mux2_1
XFILLER_218_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26640_ clknet_leaf_13_B_in_serial_clk _00443_ net5 VGND VGND VPWR VPWR deser_B.word_buffer\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23852_ _10443_ _10444_ VGND VGND VPWR VPWR _10445_ sky130_fd_sc_hd__or2_1
XFILLER_217_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22803_ _09478_ _09484_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__and2_1
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26571_ clknet_leaf_24_A_in_serial_clk _00374_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_23783_ _10382_ _10384_ _10386_ systolic_inst.acc_wires\[0\]\[13\] _11258_ VGND VGND
+ VPWR VPWR _01943_ sky130_fd_sc_hd__a32o_1
XFILLER_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20995_ _07834_ _07867_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_64_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
X_25522_ systolic_inst.cycle_cnt\[31\] _11243_ _11241_ VGND VGND VPWR VPWR _11244_
+ sky130_fd_sc_hd__mux2_1
XFILLER_213_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28310_ clknet_leaf_347_clk _02108_ VGND VGND VPWR VPWR systolic_inst.A_shift\[29\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_22734_ _09416_ _09417_ _09395_ _09398_ VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__o211ai_2
XFILLER_164_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29290_ clknet_leaf_315_clk _03088_ net142 VGND VGND VPWR VPWR C_out\[262\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28241_ clknet_leaf_134_clk _02039_ VGND VGND VPWR VPWR systolic_inst.B_shift\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25453_ systolic_inst.cycle_cnt\[7\] systolic_inst.cycle_cnt\[6\] _11195_ VGND VGND
+ VPWR VPWR _11199_ sky130_fd_sc_hd__and3_1
XFILLER_201_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22665_ _09370_ _09371_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__nand2_1
XFILLER_52_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24404_ net114 ser_C.shift_reg\[30\] VGND VGND VPWR VPWR _10672_ sky130_fd_sc_hd__and2_1
XFILLER_142_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28172_ clknet_leaf_79_clk _01970_ VGND VGND VPWR VPWR systolic_inst.B_shift\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_21616_ _08390_ _08425_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__or2_1
XFILLER_90_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25384_ _11161_ systolic_inst.B_shift\[14\]\[7\] net71 VGND VGND VPWR VPWR _02769_
+ sky130_fd_sc_hd__mux2_1
X_22596_ _09309_ _09311_ _09308_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27123_ clknet_leaf_3_B_in_serial_clk _00921_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24335_ systolic_inst.A_shift\[10\]\[7\] A_in\[39\] net59 VGND VGND VPWR VPWR _10641_
+ sky130_fd_sc_hd__mux2_1
X_21547_ _08355_ _08358_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27054_ clknet_leaf_27_B_in_serial_clk _00852_ net135 VGND VGND VPWR VPWR deser_B.shift_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_24266_ systolic_inst.B_shift\[17\]\[1\] net72 _11333_ B_in\[105\] VGND VGND VPWR
+ VPWR _02203_ sky130_fd_sc_hd__a22o_1
XFILLER_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21478_ systolic_inst.B_outs\[2\]\[6\] systolic_inst.B_shift\[2\]\[6\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__mux2_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26005_ systolic_inst.acc_wires\[15\]\[1\] ser_C.parallel_data\[481\] net23 VGND
+ VGND VPWR VPWR _03307_ sky130_fd_sc_hd__mux2_1
X_23217_ systolic_inst.acc_wires\[1\]\[20\] systolic_inst.acc_wires\[1\]\[21\] systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _09868_ sky130_fd_sc_hd__o21a_1
X_20429_ systolic_inst.B_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[5\] systolic_inst.A_outs\[5\]\[6\]
+ systolic_inst.B_outs\[5\]\[3\] VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__a22oi_1
XFILLER_134_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24197_ systolic_inst.B_shift\[22\]\[4\] net71 _11333_ B_in\[116\] VGND VGND VPWR
+ VPWR _02158_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_112_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23148_ _09794_ _09800_ _09802_ VGND VGND VPWR VPWR _09809_ sky130_fd_sc_hd__o21a_1
XFILLER_161_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23079_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[1\]\[2\]
+ VGND VGND VPWR VPWR _09750_ sky130_fd_sc_hd__or2_1
X_27956_ clknet_leaf_170_clk _01754_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15970_ systolic_inst.B_outs\[11\]\[3\] systolic_inst.B_outs\[7\]\[3\] net119 VGND
+ VGND VPWR VPWR _01149_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14921_ systolic_inst.A_outs\[14\]\[2\] systolic_inst.B_outs\[14\]\[6\] _11264_ systolic_inst.A_outs\[14\]\[1\]
+ VGND VGND VPWR VPWR _12043_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26907_ clknet_leaf_11_A_in_serial_clk _00705_ net135 VGND VGND VPWR VPWR deser_A.serial_word\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27887_ clknet_leaf_309_clk _01685_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29626_ clknet_leaf_9_B_in_serial_clk _03421_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_17640_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[9\] systolic_inst.acc_wires\[10\]\[9\]
+ _04874_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__a21oi_1
X_26838_ clknet_leaf_83_clk _00640_ net144 VGND VGND VPWR VPWR B_in\[110\] sky130_fd_sc_hd__dfrtp_1
X_14852_ _11942_ _11975_ VGND VGND VPWR VPWR _11976_ sky130_fd_sc_hd__nor2_1
XFILLER_29_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13803_ B_in\[110\] deser_B.word_buffer\[110\] net88 VGND VGND VPWR VPWR _00640_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29557_ clknet_leaf_16_B_in_serial_clk _03352_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14783_ _11888_ _11894_ _11897_ VGND VGND VPWR VPWR _11910_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_82_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17571_ _04819_ _04820_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__xnor2_1
X_26769_ clknet_leaf_95_clk _00571_ net5 VGND VGND VPWR VPWR B_in\[41\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_clk clknet_5_17__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_17_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_231_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19310_ net105 _06370_ _06371_ _06341_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__o31a_1
X_28508_ clknet_leaf_111_clk _02306_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_13734_ B_in\[41\] deser_B.word_buffer\[41\] net84 VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__mux2_1
X_16522_ net67 _03875_ _03876_ systolic_inst.acc_wires\[12\]\[22\] net108 VGND VGND
+ VPWR VPWR _01192_ sky130_fd_sc_hd__a32o_1
XFILLER_1_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_231_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_231_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29488_ clknet_leaf_279_clk _03286_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[460\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19241_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[9\] _06304_ net119
+ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13665_ deser_B.word_buffer\[101\] deser_B.serial_word\[101\] net123 VGND VGND VPWR
+ VPWR _00502_ sky130_fd_sc_hd__mux2_1
XFILLER_189_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16453_ _03817_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__inv_2
X_28439_ clknet_leaf_35_clk _02237_ VGND VGND VPWR VPWR systolic_inst.A_shift\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15404_ _12464_ _12465_ VGND VGND VPWR VPWR _12466_ sky130_fd_sc_hd__nand2_1
X_19172_ systolic_inst.B_outs\[7\]\[0\] systolic_inst.B_outs\[7\]\[1\] systolic_inst.A_outs\[7\]\[7\]
+ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__o21a_1
X_16384_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[3\] systolic_inst.acc_wires\[12\]\[3\]
+ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__or2_1
X_13596_ deser_B.word_buffer\[32\] deser_B.serial_word\[32\] net124 VGND VGND VPWR
+ VPWR _00433_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15335_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[28\]
+ VGND VGND VPWR VPWR _12421_ sky130_fd_sc_hd__nand2_1
X_18123_ _05220_ _05280_ _05278_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_229_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_229_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15266_ _12360_ _12362_ VGND VGND VPWR VPWR _12363_ sky130_fd_sc_hd__xnor2_1
X_18054_ _05188_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__nand2_1
XANTENNA_3 _10506_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14217_ systolic_inst.B_outs\[15\]\[2\] systolic_inst.A_outs\[15\]\[4\] systolic_inst.A_outs\[15\]\[5\]
+ systolic_inst.B_outs\[15\]\[1\] VGND VGND VPWR VPWR _11405_ sky130_fd_sc_hd__a22oi_1
X_17005_ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__inv_2
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15197_ _12298_ _12301_ VGND VGND VPWR VPWR _12303_ sky130_fd_sc_hd__nand2_1
XFILLER_153_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_9__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_5_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_14148_ systolic_inst.A_outs\[15\]\[0\] systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[1\]
+ systolic_inst.B_outs\[15\]\[2\] VGND VGND VPWR VPWR _11340_ sky130_fd_sc_hd__nand4_2
XFILLER_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14079_ deser_B.shift_reg\[113\] deser_B.shift_reg\[114\] deser_B.receiving VGND
+ VGND VPWR VPWR _00905_ sky130_fd_sc_hd__mux2_1
X_18956_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[8\]\[23\]
+ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__xor2_1
XFILLER_234_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17907_ _05055_ _05057_ _05100_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__and3_1
XFILLER_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18887_ _05993_ _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__nand2_1
XFILLER_230_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_175_Right_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17838_ systolic_inst.B_outs\[9\]\[0\] systolic_inst.A_outs\[9\]\[4\] VGND VGND VPWR
+ VPWR _05035_ sky130_fd_sc_hd__nand2_1
XFILLER_242_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17769_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_46_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19508_ net62 _06548_ _06549_ systolic_inst.acc_wires\[7\]\[15\] net105 VGND VGND
+ VPWR VPWR _01505_ sky130_fd_sc_hd__a32o_1
XFILLER_35_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20780_ _07664_ _07684_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__nor2_1
XFILLER_50_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19439_ net62 _06488_ _06490_ systolic_inst.acc_wires\[7\]\[5\] net105 VGND VGND
+ VPWR VPWR _01495_ sky130_fd_sc_hd__a32o_1
XFILLER_168_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_214_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22450_ _09125_ _09167_ _09166_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__o21a_1
XFILLER_50_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21401_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[4\]\[22\]
+ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__or2_1
XFILLER_202_1227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22381_ systolic_inst.B_outs\[2\]\[2\] systolic_inst.A_outs\[2\]\[7\] _09094_ _09060_
+ VGND VGND VPWR VPWR _09122_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_152_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24120_ systolic_inst.B_shift\[27\]\[7\] net72 _11333_ B_in\[127\] VGND VGND VPWR
+ VPWR _02105_ sky130_fd_sc_hd__a22o_1
X_21332_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[4\]\[11\]
+ _08180_ _08183_ _08184_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__a221oi_1
XFILLER_11_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24051_ systolic_inst.B_shift\[4\]\[5\] B_in\[5\] _00008_ VGND VGND VPWR VPWR _10543_
+ sky130_fd_sc_hd__mux2_1
X_21263_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[4\]\[2\]
+ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__nand2_1
XFILLER_11_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23002_ _09678_ VGND VGND VPWR VPWR _09679_ sky130_fd_sc_hd__inv_2
XFILLER_85_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20214_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[30\]
+ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__or2_1
XFILLER_85_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21194_ systolic_inst.B_outs\[4\]\[6\] systolic_inst.A_outs\[4\]\[7\] VGND VGND VPWR
+ VPWR _08062_ sky130_fd_sc_hd__nand2_1
XFILLER_116_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27810_ clknet_leaf_140_clk _01608_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_20145_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[20\]
+ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__or2_1
XFILLER_213_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28790_ clknet_leaf_201_clk _02588_ net147 VGND VGND VPWR VPWR ser_C.shift_reg\[338\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27741_ clknet_leaf_209_clk _01539_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24953_ C_out\[303\] net103 net76 ser_C.shift_reg\[303\] _10946_ VGND VGND VPWR VPWR
+ _02553_ sky130_fd_sc_hd__a221o_1
XFILLER_213_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20076_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[6\]\[10\]
+ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__nand2_1
XFILLER_100_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23904_ systolic_inst.B_shift\[17\]\[4\] B_in\[76\] _00008_ VGND VGND VPWR VPWR _10485_
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27672_ clknet_leaf_147_clk _01470_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24884_ net110 ser_C.shift_reg\[270\] VGND VGND VPWR VPWR _10912_ sky130_fd_sc_hd__and2_1
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29411_ clknet_leaf_234_clk _03209_ net147 VGND VGND VPWR VPWR C_out\[383\] sky130_fd_sc_hd__dfrtp_1
X_23835_ _10428_ _10429_ VGND VGND VPWR VPWR _10430_ sky130_fd_sc_hd__and2_1
X_26623_ clknet_leaf_22_B_in_serial_clk _00426_ net137 VGND VGND VPWR VPWR deser_B.word_buffer\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk clknet_5_18__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29342_ clknet_leaf_223_clk _03140_ net149 VGND VGND VPWR VPWR C_out\[314\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26554_ clknet_leaf_27_A_in_serial_clk _00357_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_23766_ _10370_ _10371_ VGND VGND VPWR VPWR _10372_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20978_ systolic_inst.B_outs\[4\]\[0\] systolic_inst.B_outs\[4\]\[7\] systolic_inst.A_outs\[4\]\[7\]
+ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__nand3_4
XFILLER_92_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25505_ systolic_inst.cycle_cnt\[25\] _11231_ VGND VGND VPWR VPWR _11233_ sky130_fd_sc_hd__and2_1
X_22717_ _11258_ _09400_ _09401_ _09402_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__o31ai_1
X_29273_ clknet_leaf_189_clk _03071_ net146 VGND VGND VPWR VPWR C_out\[245\] sky130_fd_sc_hd__dfrtp_1
X_26485_ clknet_leaf_9_A_in_serial_clk _00288_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23697_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[0\]\[0\]
+ _10311_ _10312_ VGND VGND VPWR VPWR _10313_ sky130_fd_sc_hd__and4_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25436_ systolic_inst.ce_local _11186_ _11187_ _11307_ systolic_inst.cycle_cnt\[1\]
+ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__a32o_1
X_28224_ clknet_leaf_98_clk _02022_ VGND VGND VPWR VPWR systolic_inst.B_shift\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13450_ deser_A.shift_reg\[14\] deser_A.shift_reg\[15\] deser_A.receiving VGND VGND
+ VPWR VPWR _00287_ sky130_fd_sc_hd__mux2_1
X_22648_ _09350_ _09354_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__nor2_1
XFILLER_139_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28155_ clknet_leaf_104_clk _01953_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25367_ ser_C.parallel_data\[510\] net98 net78 ser_C.shift_reg\[510\] _11153_ VGND
+ VGND VPWR VPWR _02760_ sky130_fd_sc_hd__a221o_1
X_13381_ A_in\[90\] deser_A.word_buffer\[90\] net92 VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__mux2_1
X_22579_ _09298_ _09299_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__nand2_1
XFILLER_210_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15120_ _12146_ _12234_ VGND VGND VPWR VPWR _12236_ sky130_fd_sc_hd__and2_1
X_27106_ clknet_leaf_4_B_in_serial_clk _00904_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_24318_ _10632_ systolic_inst.A_shift\[10\]\[6\] net71 VGND VGND VPWR VPWR _02232_
+ sky130_fd_sc_hd__mux2_1
X_28086_ clknet_leaf_118_clk _01884_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25298_ net111 ser_C.shift_reg\[477\] VGND VGND VPWR VPWR _11119_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27037_ clknet_leaf_14_B_in_serial_clk _00835_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_15051_ _12134_ _12138_ _12169_ VGND VGND VPWR VPWR _12170_ sky130_fd_sc_hd__or3_1
X_24249_ systolic_inst.A_shift\[17\]\[0\] net70 net83 systolic_inst.A_shift\[18\]\[0\]
+ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__a22o_1
XFILLER_107_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_224_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14002_ deser_B.shift_reg\[36\] deser_B.shift_reg\[37\] deser_B.receiving VGND VGND
+ VPWR VPWR _00828_ sky130_fd_sc_hd__mux2_1
XFILLER_107_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_79_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18810_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[8\]\[2\]
+ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_220_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19790_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[6\] VGND VGND VPWR
+ VPWR _06791_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28988_ clknet_leaf_56_clk _02786_ VGND VGND VPWR VPWR systolic_inst.A_shift\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18741_ systolic_inst.A_outs\[8\]\[6\] _11259_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__or2_1
X_27939_ clknet_leaf_170_clk _01737_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15953_ _12968_ _12971_ VGND VGND VPWR VPWR _12973_ sky130_fd_sc_hd__or2_1
XFILLER_7_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_A_in_serial_clk clknet_2_3__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_13_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_3_1209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14904_ net107 systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[7\] _12025_
+ _12026_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__a22o_1
XFILLER_236_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18672_ net108 systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[10\] VGND
+ VGND VPWR VPWR _05799_ sky130_fd_sc_hd__nand2_1
X_15884_ _12912_ _12913_ VGND VGND VPWR VPWR _12914_ sky130_fd_sc_hd__and2_1
XFILLER_149_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29609_ clknet_leaf_24_B_in_serial_clk _03404_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_17623_ _04862_ _04863_ _04864_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__nand3_1
XFILLER_188_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14835_ _11928_ _11931_ _11957_ net118 VGND VGND VPWR VPWR _11960_ sky130_fd_sc_hd__o31a_1
XFILLER_17_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_clk clknet_5_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_218_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_218_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17554_ _04741_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__xnor2_1
X_14766_ _11891_ _11892_ _11893_ VGND VGND VPWR VPWR _11894_ sky130_fd_sc_hd__a21o_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16505_ _03844_ _03847_ _03861_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__and3_1
X_13717_ B_in\[24\] deser_B.word_buffer\[24\] net85 VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14697_ _11849_ _11850_ VGND VGND VPWR VPWR _11851_ sky130_fd_sc_hd__nor2_1
X_17485_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[7\] _04712_ _04676_
+ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__a31o_1
X_19224_ _06287_ _06286_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__nand2b_1
XFILLER_34_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16436_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[12\]\[11\]
+ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__nand2_1
X_13648_ deser_B.word_buffer\[84\] deser_B.serial_word\[84\] net124 VGND VGND VPWR
+ VPWR _00485_ sky130_fd_sc_hd__mux2_1
XFILLER_72_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19155_ _06184_ _06220_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__or2_1
X_13579_ deser_B.word_buffer\[15\] deser_B.serial_word\[15\] net124 VGND VGND VPWR
+ VPWR _00416_ sky130_fd_sc_hd__mux2_1
X_16367_ net115 _03742_ _03743_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18106_ _05293_ _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__nor2_1
X_15318_ _12401_ _12403_ _12405_ VGND VGND VPWR VPWR _12407_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19086_ _06151_ _06153_ systolic_inst.B_outs\[7\]\[2\] systolic_inst.A_outs\[7\]\[3\]
+ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__and4b_1
X_16298_ _03627_ _03677_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__xor2_1
XFILLER_195_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18037_ systolic_inst.A_outs\[9\]\[3\] systolic_inst.A_outs\[9\]\[4\] systolic_inst.B_outs\[9\]\[6\]
+ systolic_inst.B_outs\[9\]\[7\] VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__and4b_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15249_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[15\]
+ VGND VGND VPWR VPWR _12348_ sky130_fd_sc_hd__and2_1
XFILLER_114_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19988_ _06981_ _06982_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__nand2_1
XFILLER_140_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18939_ systolic_inst.acc_wires\[8\]\[16\] systolic_inst.acc_wires\[8\]\[17\] systolic_inst.acc_wires\[8\]\[18\]
+ systolic_inst.acc_wires\[8\]\[19\] systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__o41a_1
XFILLER_234_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_203_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21950_ _08731_ _08733_ _08735_ _08738_ VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__or4_1
XFILLER_239_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_228_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20901_ _07759_ _07776_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21881_ _08670_ _08673_ _08677_ _08678_ VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__o211a_1
XFILLER_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_clk clknet_5_16__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_43_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23620_ _10228_ _10240_ VGND VGND VPWR VPWR _10241_ sky130_fd_sc_hd__or2_1
XFILLER_54_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20832_ systolic_inst.A_outs\[4\]\[5\] systolic_inst.A_shift\[8\]\[5\] net121 VGND
+ VGND VPWR VPWR _01655_ sky130_fd_sc_hd__mux2_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23551_ _10130_ _10132_ _10171_ VGND VGND VPWR VPWR _10174_ sky130_fd_sc_hd__nor3_1
X_20763_ _07670_ _07669_ systolic_inst.acc_wires\[5\]\[21\] net106 VGND VGND VPWR
+ VPWR _01639_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22502_ _09231_ _09232_ _09233_ VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_154_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26270_ clknet_leaf_21_A_in_serial_clk _00078_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[68\]
+ sky130_fd_sc_hd__dfrtp_1
X_23482_ systolic_inst.A_outs\[0\]\[4\] systolic_inst.B_outs\[0\]\[5\] _10025_ VGND
+ VGND VPWR VPWR _10106_ sky130_fd_sc_hd__and3_1
XFILLER_52_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20694_ _07610_ _07611_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25221_ C_out\[437\] net101 net73 ser_C.shift_reg\[437\] _11080_ VGND VGND VPWR VPWR
+ _02687_ sky130_fd_sc_hd__a221o_1
XFILLER_104_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22433_ _09124_ _09172_ VGND VGND VPWR VPWR _09173_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25152_ net110 ser_C.shift_reg\[404\] VGND VGND VPWR VPWR _11046_ sky130_fd_sc_hd__and2_1
X_22364_ _09096_ _09104_ VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__xnor2_1
XFILLER_191_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24103_ systolic_inst.B_shift\[23\]\[7\] B_in\[63\] _00008_ VGND VGND VPWR VPWR _10561_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21315_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[4\]\[10\]
+ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__or2_1
X_25083_ C_out\[368\] net97 net77 ser_C.shift_reg\[368\] _11011_ VGND VGND VPWR VPWR
+ _02618_ sky130_fd_sc_hd__a221o_1
X_22295_ _09001_ _09003_ _09038_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__a21o_1
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_211_Right_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24034_ _10534_ systolic_inst.B_shift\[4\]\[4\] net72 VGND VGND VPWR VPWR _02046_
+ sky130_fd_sc_hd__mux2_1
X_28911_ clknet_leaf_280_clk _02709_ net139 VGND VGND VPWR VPWR ser_C.shift_reg\[459\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_151_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21246_ _08094_ _08095_ _08097_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__o21a_1
XFILLER_117_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28842_ clknet_leaf_333_clk _02640_ net136 VGND VGND VPWR VPWR ser_C.shift_reg\[390\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21177_ _08044_ _08045_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20128_ net106 systolic_inst.acc_wires\[6\]\[16\] _07102_ _07104_ VGND VGND VPWR
+ VPWR _01570_ sky130_fd_sc_hd__a22o_1
X_28773_ clknet_leaf_295_clk _02571_ net138 VGND VGND VPWR VPWR ser_C.shift_reg\[321\]
+ sky130_fd_sc_hd__dfrtp_1
X_25985_ systolic_inst.acc_wires\[14\]\[13\] ser_C.parallel_data\[461\] net26 VGND
+ VGND VPWR VPWR _03287_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27724_ clknet_leaf_215_clk _01522_ net149 VGND VGND VPWR VPWR systolic_inst.A_outs\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_20059_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[7\] systolic_inst.acc_wires\[6\]\[7\]
+ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__or2_1
X_24936_ net111 ser_C.shift_reg\[296\] VGND VGND VPWR VPWR _10938_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_107_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27655_ clknet_leaf_303_clk _01453_ net141 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24867_ C_out\[260\] net101 net73 ser_C.shift_reg\[260\] _10903_ VGND VGND VPWR VPWR
+ _02510_ sky130_fd_sc_hd__a221o_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26606_ clknet_leaf_15_B_in_serial_clk _00409_ net152 VGND VGND VPWR VPWR deser_B.word_buffer\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14620_ net61 _11784_ VGND VGND VPWR VPWR _11785_ sky130_fd_sc_hd__nor2_1
X_23818_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[19\]
+ VGND VGND VPWR VPWR _10416_ sky130_fd_sc_hd__xnor2_1
X_27586_ clknet_leaf_215_clk _01384_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_24798_ net112 ser_C.shift_reg\[227\] VGND VGND VPWR VPWR _10869_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_64_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14551_ _11725_ VGND VGND VPWR VPWR _11726_ sky130_fd_sc_hd__inv_2
X_29325_ clknet_leaf_304_clk _03123_ net139 VGND VGND VPWR VPWR C_out\[297\] sky130_fd_sc_hd__dfrtp_1
XFILLER_242_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23749_ _10352_ _10355_ VGND VGND VPWR VPWR _10357_ sky130_fd_sc_hd__nand2_1
XFILLER_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26537_ clknet_leaf_21_A_in_serial_clk _00340_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_199_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13502_ deser_A.shift_reg\[66\] deser_A.shift_reg\[67\] net129 VGND VGND VPWR VPWR
+ _00339_ sky130_fd_sc_hd__mux2_1
X_29256_ clknet_leaf_196_clk _03054_ net146 VGND VGND VPWR VPWR C_out\[228\] sky130_fd_sc_hd__dfrtp_1
X_14482_ _11661_ _11662_ VGND VGND VPWR VPWR _11663_ sky130_fd_sc_hd__and2b_1
X_17270_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[5\] _04529_ net118
+ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__mux2_1
X_26468_ clknet_leaf_1_A_in_serial_clk _00002_ net132 VGND VGND VPWR VPWR deser_A.serial_word_ready
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_105_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28207_ clknet_leaf_103_clk _02005_ VGND VGND VPWR VPWR systolic_inst.B_shift\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16221_ _03601_ _03602_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__xnor2_1
X_13433_ _11310_ _11315_ _11317_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__and3_1
X_25419_ systolic_inst.A_shift\[1\]\[1\] A_in\[1\] net59 VGND VGND VPWR VPWR _11179_
+ sky130_fd_sc_hd__mux2_1
X_29187_ clknet_leaf_136_clk _02985_ net142 VGND VGND VPWR VPWR C_out\[159\] sky130_fd_sc_hd__dfrtp_1
X_26399_ clknet_leaf_31_clk _00206_ net137 VGND VGND VPWR VPWR A_in\[67\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload209 clknet_leaf_42_clk VGND VGND VPWR VPWR clkload209/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16152_ _13070_ _03495_ _03497_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__a21oi_1
X_28138_ clknet_leaf_125_clk _01936_ net144 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13364_ A_in\[73\] deser_A.word_buffer\[73\] net94 VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__mux2_1
X_15103_ _12177_ _12219_ VGND VGND VPWR VPWR _12220_ sky130_fd_sc_hd__xnor2_1
X_16083_ _13047_ _13050_ _13077_ _13078_ VGND VGND VPWR VPWR _13079_ sky130_fd_sc_hd__a211oi_2
X_28069_ clknet_leaf_119_clk _01867_ net149 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13295_ A_in\[4\] deser_A.word_buffer\[4\] net94 VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__mux2_1
X_19911_ _06892_ _06908_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__xor2_1
X_15034_ _12152_ _12151_ VGND VGND VPWR VPWR _12153_ sky130_fd_sc_hd__nand2b_1
XFILLER_218_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19842_ _06824_ _06841_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__xor2_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19773_ _06741_ _06773_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__xnor2_1
XFILLER_231_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16985_ net69 _04293_ _04295_ systolic_inst.acc_wires\[11\]\[2\] net105 VGND VGND
+ VPWR VPWR _01236_ sky130_fd_sc_hd__a32o_1
XFILLER_84_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18724_ _05803_ _05819_ _05817_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__o21a_1
X_15936_ _12942_ _12944_ _12956_ _12957_ _12950_ VGND VGND VPWR VPWR _12958_ sky130_fd_sc_hd__a311oi_4
XFILLER_37_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18655_ _05739_ _05747_ _05746_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__a21bo_1
XFILLER_188_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15867_ _12899_ VGND VGND VPWR VPWR _12900_ sky130_fd_sc_hd__inv_2
XFILLER_64_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17606_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[10\]\[5\]
+ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__nand2_1
X_14818_ systolic_inst.B_outs\[14\]\[2\] systolic_inst.A_outs\[14\]\[3\] VGND VGND
+ VPWR VPWR _11943_ sky130_fd_sc_hd__nand2_1
X_18586_ _05714_ _05713_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__and2b_1
X_15798_ _12838_ _12839_ _12840_ VGND VGND VPWR VPWR _12841_ sky130_fd_sc_hd__a21o_1
XFILLER_225_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17537_ _04787_ _04788_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_190_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14749_ systolic_inst.B_outs\[13\]\[1\] systolic_inst.B_outs\[9\]\[1\] net115 VGND
+ VGND VPWR VPWR _01019_ sky130_fd_sc_hd__mux2_1
XFILLER_178_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17468_ _04719_ _04720_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_220_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19207_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[8\] _06271_ net119
+ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__mux2_1
XFILLER_32_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16419_ _03787_ _03786_ systolic_inst.acc_wires\[12\]\[8\] net108 VGND VGND VPWR
+ VPWR _01178_ sky130_fd_sc_hd__a2bb2o_1
X_17399_ _04652_ _04653_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19138_ _11261_ _06203_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19069_ _06135_ _06136_ _06129_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_8_clk clknet_5_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_209_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21100_ _07962_ _07970_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_8_A_in_serial_clk clknet_2_2__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_8_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_209_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22080_ systolic_inst.A_outs\[2\]\[2\] systolic_inst.A_outs\[1\]\[2\] net122 VGND
+ VGND VPWR VPWR _01780_ sky130_fd_sc_hd__mux2_1
XFILLER_218_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21031_ _07901_ _07902_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__xor2_1
XFILLER_101_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22982_ _09657_ _09658_ VGND VGND VPWR VPWR _09659_ sky130_fd_sc_hd__nor2_1
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25770_ systolic_inst.acc_wires\[7\]\[22\] C_out\[246\] net44 VGND VGND VPWR VPWR
+ _03072_ sky130_fd_sc_hd__mux2_1
X_21933_ _08720_ _08722_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__nand2_1
X_24721_ C_out\[187\] net99 net79 ser_C.shift_reg\[187\] _10830_ VGND VGND VPWR VPWR
+ _02437_ sky130_fd_sc_hd__a221o_1
XFILLER_28_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24652_ net7 ser_C.shift_reg\[154\] VGND VGND VPWR VPWR _10796_ sky130_fd_sc_hd__and2_1
X_27440_ clknet_leaf_245_clk _01238_ net145 VGND VGND VPWR VPWR systolic_inst.acc_wires\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_21864_ _08662_ _08665_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23603_ _10223_ _10221_ VGND VGND VPWR VPWR _10224_ sky130_fd_sc_hd__nand2b_1
XFILLER_82_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20815_ systolic_inst.acc_wires\[5\]\[28\] systolic_inst.acc_wires\[5\]\[29\] systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__o21ai_1
X_24583_ C_out\[118\] net100 net82 ser_C.shift_reg\[118\] _10761_ VGND VGND VPWR VPWR
+ _02368_ sky130_fd_sc_hd__a221o_1
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27371_ clknet_leaf_344_clk _01169_ net131 VGND VGND VPWR VPWR systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_21795_ _08586_ _08599_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29110_ clknet_leaf_160_clk _02908_ net150 VGND VGND VPWR VPWR C_out\[82\] sky130_fd_sc_hd__dfrtp_1
XFILLER_169_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23534_ systolic_inst.A_outs\[0\]\[4\] systolic_inst.B_outs\[0\]\[6\] _10155_ VGND
+ VGND VPWR VPWR _10157_ sky130_fd_sc_hd__a21oi_1
X_26322_ clknet_leaf_0_A_in_serial_clk _00130_ net132 VGND VGND VPWR VPWR deser_A.word_buffer\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_20746_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[19\]
+ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29041_ clknet_leaf_100_clk _02839_ net152 VGND VGND VPWR VPWR C_out\[13\] sky130_fd_sc_hd__dfrtp_1
X_26253_ clknet_leaf_3_A_in_serial_clk _00061_ net133 VGND VGND VPWR VPWR deser_A.word_buffer\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_23465_ _10044_ _10047_ _10088_ VGND VGND VPWR VPWR _10090_ sky130_fd_sc_hd__nand3_1
XFILLER_221_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20677_ _07592_ _07595_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__nand2_1
X_25204_ net110 ser_C.shift_reg\[430\] VGND VGND VPWR VPWR _11072_ sky130_fd_sc_hd__and2_1
XFILLER_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22416_ _09154_ _09155_ VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26184_ _11250_ _11251_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__nor2_1
X_23396_ _11258_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[6\] VGND
+ VGND VPWR VPWR _10023_ sky130_fd_sc_hd__nand2_1
XFILLER_52_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25135_ C_out\[394\] net101 net73 ser_C.shift_reg\[394\] _11037_ VGND VGND VPWR VPWR
+ _02644_ sky130_fd_sc_hd__a221o_1
X_22347_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[10\] _09089_ net122
+ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__mux2_1
XFILLER_192_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25066_ net112 ser_C.shift_reg\[361\] VGND VGND VPWR VPWR _11003_ sky130_fd_sc_hd__and2_1
X_22278_ _08985_ _09021_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__nor2_1
XFILLER_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24017_ systolic_inst.B_shift\[6\]\[0\] _11332_ net83 systolic_inst.B_shift\[10\]\[0\]
+ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__a22o_1
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21229_ _08094_ _08095_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28825_ clknet_leaf_238_clk _02623_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[373\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16770_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[8\] VGND
+ VGND VPWR VPWR _04091_ sky130_fd_sc_hd__and2_1
X_28756_ clknet_leaf_223_clk _02554_ net140 VGND VGND VPWR VPWR ser_C.shift_reg\[304\]
+ sky130_fd_sc_hd__dfrtp_1
X_13982_ deser_B.shift_reg\[16\] deser_B.shift_reg\[17\] net125 VGND VGND VPWR VPWR
+ _00808_ sky130_fd_sc_hd__mux2_1
X_25968_ systolic_inst.acc_wires\[13\]\[28\] ser_C.parallel_data\[444\] net26 VGND
+ VGND VPWR VPWR _03270_ sky130_fd_sc_hd__mux2_1
XFILLER_59_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27707_ clknet_leaf_190_clk _01505_ net146 VGND VGND VPWR VPWR systolic_inst.acc_wires\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15721_ systolic_inst.A_outs\[13\]\[6\] _11272_ _12746_ _12749_ _12772_ VGND VGND
+ VPWR VPWR _12773_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_66_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24919_ C_out\[286\] net103 net75 ser_C.shift_reg\[286\] _10929_ VGND VGND VPWR VPWR
+ _02536_ sky130_fd_sc_hd__a221o_1
X_28687_ clknet_leaf_192_clk _02485_ net146 VGND VGND VPWR VPWR ser_C.shift_reg\[235\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_215_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25899_ systolic_inst.acc_wires\[11\]\[23\] C_out\[375\] net41 VGND VGND VPWR VPWR
+ _03201_ sky130_fd_sc_hd__mux2_1
XFILLER_233_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _05571_ _05572_ _05562_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__a21o_1
XFILLER_74_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15652_ _12667_ _12669_ _12706_ VGND VGND VPWR VPWR _12707_ sky130_fd_sc_hd__and3_1
X_27638_ clknet_leaf_315_clk _01436_ net137 VGND VGND VPWR VPWR systolic_inst.acc_wires\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _11762_ _11764_ _11760_ VGND VGND VPWR VPWR _11770_ sky130_fd_sc_hd__a21bo_1
X_18371_ _05527_ _05529_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_17_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15583_ _12610_ _12637_ VGND VGND VPWR VPWR _12640_ sky130_fd_sc_hd__xnor2_1
X_27569_ clknet_leaf_298_clk _01367_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29308_ clknet_leaf_313_clk _03106_ net141 VGND VGND VPWR VPWR C_out\[280\] sky130_fd_sc_hd__dfrtp_1
X_17322_ _04543_ _04578_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14534_ _11710_ VGND VGND VPWR VPWR _11711_ sky130_fd_sc_hd__inv_2
XFILLER_183_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29239_ clknet_leaf_177_clk _03037_ net148 VGND VGND VPWR VPWR C_out\[211\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17253_ systolic_inst.B_outs\[10\]\[2\] systolic_inst.A_outs\[10\]\[3\] VGND VGND
+ VPWR VPWR _04513_ sky130_fd_sc_hd__and2_1
XFILLER_202_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14465_ _11645_ _11646_ VGND VGND VPWR VPWR _11647_ sky130_fd_sc_hd__and2_1
XFILLER_35_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16204_ net108 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[9\] VGND
+ VGND VPWR VPWR _03588_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13416_ A_in\[125\] deser_A.word_buffer\[125\] net92 VGND VGND VPWR VPWR _00264_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14396_ _11541_ _11544_ _11579_ VGND VGND VPWR VPWR _11580_ sky130_fd_sc_hd__a21oi_1
X_17184_ systolic_inst.A_outs\[10\]\[6\] systolic_inst.A_outs\[9\]\[6\] net120 VGND
+ VGND VPWR VPWR _01272_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16135_ _03515_ _03518_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__xnor2_1
X_13347_ A_in\[56\] deser_A.word_buffer\[56\] net91 VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__mux2_1
XFILLER_128_888 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16066_ _13060_ _13061_ VGND VGND VPWR VPWR _13062_ sky130_fd_sc_hd__or2_1
X_13278_ deser_A.word_buffer\[116\] deser_A.serial_word\[116\] deser_A.serial_word_ready
+ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__mux2_1
XFILLER_142_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_183_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15017_ _12135_ _12136_ VGND VGND VPWR VPWR _12137_ sky130_fd_sc_hd__and2b_1
XFILLER_111_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19825_ systolic_inst.B_outs\[6\]\[2\] systolic_inst.A_outs\[6\]\[7\] VGND VGND VPWR
+ VPWR _06825_ sky130_fd_sc_hd__nand2_4
XFILLER_155_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_229_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19756_ systolic_inst.A_outs\[6\]\[0\] systolic_inst.B_outs\[6\]\[7\] VGND VGND VPWR
+ VPWR _06758_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_196_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16968_ net105 systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[15\] _04274_
+ _04281_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__a22o_1
XFILLER_204_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18707_ systolic_inst.B_outs\[8\]\[2\] systolic_inst.A_outs\[8\]\[7\] _05804_ _05768_
+ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__a31o_1
X_15919_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[25\]
+ VGND VGND VPWR VPWR _12944_ sky130_fd_sc_hd__xor2_2
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19687_ _06670_ _06690_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_192_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16899_ _04213_ _04214_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_192_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18638_ _05695_ _05763_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__and2_1
XFILLER_224_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_227_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18569_ _05693_ _05696_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20600_ _07464_ _07530_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21580_ _08385_ _08389_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_15_B_in_serial_clk clknet_2_3__leaf_B_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_15_B_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_20531_ _07462_ _07463_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__nand2_1
XFILLER_221_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23250_ _09894_ _09895_ VGND VGND VPWR VPWR _09896_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20462_ systolic_inst.B_outs\[5\]\[4\] systolic_inst.A_outs\[5\]\[6\] systolic_inst.A_outs\[5\]\[7\]
+ systolic_inst.B_outs\[5\]\[3\] VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__a22o_1
XFILLER_192_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22201_ _08923_ _08925_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__nand2_1
XFILLER_10_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23181_ _09835_ _09836_ VGND VGND VPWR VPWR _09838_ sky130_fd_sc_hd__nor2_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20393_ _07328_ _07329_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_149_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22132_ _08877_ _08879_ _08860_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_238_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22063_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[29\]
+ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__and2_1
XFILLER_161_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26940_ clknet_leaf_20_A_in_serial_clk _00738_ net133 VGND VGND VPWR VPWR deser_A.serial_word\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21014_ _07883_ _07886_ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__xor2_1
XFILLER_134_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26871_ clknet_leaf_15_A_in_serial_clk _00669_ net137 VGND VGND VPWR VPWR deser_A.serial_word\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_34_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28610_ clknet_leaf_133_clk _02408_ net142 VGND VGND VPWR VPWR ser_C.shift_reg\[158\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_250_clk clknet_5_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_250_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_3_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25822_ systolic_inst.acc_wires\[9\]\[10\] C_out\[298\] net15 VGND VGND VPWR VPWR
+ _03124_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29590_ clknet_leaf_12_B_in_serial_clk _03385_ net153 VGND VGND VPWR VPWR deser_B.serial_word\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28541_ clknet_leaf_163_clk _02339_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22965_ _09642_ _09641_ VGND VGND VPWR VPWR _09643_ sky130_fd_sc_hd__and2b_1
X_25753_ systolic_inst.acc_wires\[7\]\[5\] C_out\[229\] net40 VGND VGND VPWR VPWR
+ _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_28_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24704_ net113 ser_C.shift_reg\[180\] VGND VGND VPWR VPWR _10822_ sky130_fd_sc_hd__and2_1
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28472_ clknet_leaf_102_clk _02270_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_215_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21916_ net68 _08708_ _08709_ systolic_inst.acc_wires\[3\]\[7\] net106 VGND VGND
+ VPWR VPWR _01753_ sky130_fd_sc_hd__a32o_1
XFILLER_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22896_ _09520_ _09538_ _09537_ VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__o21a_1
X_25684_ systolic_inst.acc_wires\[5\]\[0\] C_out\[160\] net16 VGND VGND VPWR VPWR
+ _02986_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27423_ clknet_leaf_248_clk _01221_ net145 VGND VGND VPWR VPWR systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21847_ _08585_ _08628_ _08627_ VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__o21a_1
X_24635_ C_out\[144\] net103 net76 ser_C.shift_reg\[144\] _10787_ VGND VGND VPWR VPWR
+ _02394_ sky130_fd_sc_hd__a221o_1
XFILLER_19_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24566_ net113 ser_C.shift_reg\[111\] VGND VGND VPWR VPWR _10753_ sky130_fd_sc_hd__and2_1
X_27354_ clknet_leaf_201_clk _01152_ net147 VGND VGND VPWR VPWR systolic_inst.B_outs\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21778_ _08442_ _08582_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__or2_1
XFILLER_208_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26305_ clknet_leaf_23_A_in_serial_clk _00113_ net131 VGND VGND VPWR VPWR deser_A.word_buffer\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_184_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20729_ systolic_inst.row_loop\[1\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[5\]\[16\]
+ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__xnor2_1
X_23517_ _10099_ _10102_ VGND VGND VPWR VPWR _10141_ sky130_fd_sc_hd__nor2_1
XFILLER_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24497_ C_out\[75\] net100 net80 ser_C.shift_reg\[75\] _10718_ VGND VGND VPWR VPWR
+ _02325_ sky130_fd_sc_hd__a221o_1
XFILLER_145_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27285_ clknet_leaf_320_clk _01083_ net136 VGND VGND VPWR VPWR systolic_inst.B_outs\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_141_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29024_ clknet_leaf_92_clk _02822_ net152 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14250_ _11411_ _11413_ VGND VGND VPWR VPWR _11437_ sky130_fd_sc_hd__nand2_1
X_23448_ systolic_inst.A_outs\[0\]\[2\] systolic_inst.B_outs\[0\]\[6\] VGND VGND VPWR
+ VPWR _10073_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_134_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26236_ clknet_leaf_15_A_in_serial_clk _00044_ net137 VGND VGND VPWR VPWR deser_A.word_buffer\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ deser_A.word_buffer\[39\] deser_A.serial_word\[39\] net127 VGND VGND VPWR
+ VPWR _00049_ sky130_fd_sc_hd__mux2_1
XFILLER_137_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14181_ _11364_ _11369_ VGND VGND VPWR VPWR _11371_ sky130_fd_sc_hd__xnor2_1
X_23379_ _10003_ _10004_ _09975_ VGND VGND VPWR VPWR _10006_ sky130_fd_sc_hd__o21bai_1
X_26167_ deser_B.serial_word\[122\] deser_B.shift_reg\[122\] net56 VGND VGND VPWR
+ VPWR _03469_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13132_ deser_B.bit_idx\[6\] _11284_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__and2_4
X_25118_ net110 ser_C.shift_reg\[387\] VGND VGND VPWR VPWR _11029_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_91_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26098_ deser_B.serial_word\[53\] deser_B.shift_reg\[53\] net56 VGND VGND VPWR VPWR
+ _03400_ sky130_fd_sc_hd__mux2_1
XFILLER_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17940_ _05096_ _05131_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__xor2_1
X_25049_ C_out\[351\] net98 net78 ser_C.shift_reg\[351\] _10994_ VGND VGND VPWR VPWR
+ _02601_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_240_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_240_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17871_ _05058_ _05066_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__nor2_1
XFILLER_61_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19610_ _06629_ _06633_ _06634_ net60 VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_128_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_241_clk clknet_5_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_241_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_152_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28808_ clknet_leaf_244_clk _02606_ net145 VGND VGND VPWR VPWR ser_C.shift_reg\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16822_ _04140_ _04139_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__nand2b_1
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19541_ _06574_ _06576_ _06577_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__or3_1
XFILLER_219_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28739_ clknet_leaf_291_clk _02537_ net141 VGND VGND VPWR VPWR ser_C.shift_reg\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16753_ _04071_ _04072_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__xor2_1
XFILLER_98_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13965_ deser_A.serial_word\[126\] deser_A.shift_reg\[126\] _00002_ VGND VGND VPWR
+ VPWR _00791_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_238_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_238_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15704_ _12687_ _12725_ _12724_ VGND VGND VPWR VPWR _12757_ sky130_fd_sc_hd__a21bo_1
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19472_ net105 systolic_inst.acc_wires\[7\]\[10\] net62 _06518_ VGND VGND VPWR VPWR
+ _01500_ sky130_fd_sc_hd__a22o_1
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16684_ _04005_ _04006_ _03994_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__or3b_1
XFILLER_98_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13896_ deser_A.serial_word\[57\] deser_A.shift_reg\[57\] net58 VGND VGND VPWR VPWR
+ _00722_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18423_ net115 _05558_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__nand2_1
XFILLER_94_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_234_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15635_ systolic_inst.A_outs\[13\]\[5\] systolic_inst.B_outs\[13\]\[6\] _11272_ systolic_inst.A_outs\[13\]\[4\]
+ VGND VGND VPWR VPWR _12690_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_234_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_226_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18354_ systolic_inst.acc_wires\[9\]\[20\] systolic_inst.acc_wires\[9\]\[21\] systolic_inst.acc_wires\[9\]\[22\]
+ systolic_inst.acc_wires\[9\]\[23\] systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[15\]
+ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_44_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ systolic_inst.A_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[6\] _11272_ systolic_inst.A_outs\[13\]\[2\]
+ VGND VGND VPWR VPWR _12623_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_221_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17305_ _04507_ _04536_ _04535_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14517_ _11647_ _11673_ _11696_ VGND VGND VPWR VPWR _11697_ sky130_fd_sc_hd__a21oi_1
X_18285_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[14\] systolic_inst.acc_wires\[9\]\[14\]
+ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__or2_1
XFILLER_187_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15497_ _12552_ _12555_ VGND VGND VPWR VPWR _12556_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17236_ _04489_ _04495_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__xnor2_1
X_14448_ _11627_ _11628_ VGND VGND VPWR VPWR _11630_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_185_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17167_ _04440_ _04443_ _04446_ _04449_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_185_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14379_ systolic_inst.A_outs\[15\]\[4\] systolic_inst.B_outs\[15\]\[6\] _11273_ systolic_inst.A_outs\[15\]\[3\]
+ VGND VGND VPWR VPWR _11563_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_183_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16118_ _03503_ _03502_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__nand2b_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17098_ _04387_ _04389_ _04386_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_181_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16049_ _13043_ _13045_ VGND VGND VPWR VPWR _13046_ sky130_fd_sc_hd__nor2_1
XFILLER_233_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_237_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_233_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_232_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_232_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19808_ _06806_ _06807_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__xor2_1
XFILLER_69_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19739_ _06702_ _06732_ _06734_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__o21ba_1
XFILLER_238_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22750_ _09431_ _09432_ _09430_ VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__o21ai_1
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21701_ _08508_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__inv_2
XFILLER_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_213_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22681_ systolic_inst.B_outs\[0\]\[0\] systolic_inst.B_shift\[0\]\[0\] net121 VGND
+ VGND VPWR VPWR _01850_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24420_ net114 ser_C.shift_reg\[38\] VGND VGND VPWR VPWR _10680_ sky130_fd_sc_hd__and2_1
X_21632_ _08413_ _08415_ _08414_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__o21bai_1
XFILLER_40_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24351_ C_out\[2\] net104 _10643_ ser_C.shift_reg\[2\] _10645_ VGND VGND VPWR VPWR
+ _02252_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_299_clk clknet_5_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_299_clk
+ sky130_fd_sc_hd__clkbuf_8
X_21563_ systolic_inst.B_outs\[3\]\[1\] systolic_inst.A_outs\[3\]\[5\] systolic_inst.A_outs\[3\]\[6\]
+ systolic_inst.B_outs\[3\]\[0\] VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_170_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23302_ _09923_ _09930_ _09931_ VGND VGND VPWR VPWR _09932_ sky130_fd_sc_hd__and3b_1
XFILLER_21_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27070_ clknet_leaf_9_B_in_serial_clk _00868_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_20514_ _07446_ _07447_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__nand2_1
X_24282_ _10614_ systolic_inst.B_shift\[23\]\[4\] net72 VGND VGND VPWR VPWR _02214_
+ sky130_fd_sc_hd__mux2_1
X_21494_ _08306_ _08307_ net122 VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__o21a_1
XFILLER_88_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23233_ _09880_ _09881_ VGND VGND VPWR VPWR _09882_ sky130_fd_sc_hd__or2_1
XFILLER_153_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26021_ systolic_inst.acc_wires\[15\]\[17\] ser_C.parallel_data\[497\] net23 VGND
+ VGND VPWR VPWR _03323_ sky130_fd_sc_hd__mux2_1
X_20445_ _07363_ _07379_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__nand2_1
XFILLER_147_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23164_ _09820_ _09821_ VGND VGND VPWR VPWR _09823_ sky130_fd_sc_hd__nand2_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload370 clknet_leaf_1_B_in_serial_clk VGND VGND VPWR VPWR clkload370/X sky130_fd_sc_hd__clkbuf_8
X_20376_ _07277_ _07279_ _07312_ _07313_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__a211oi_1
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload381 clknet_leaf_23_B_in_serial_clk VGND VGND VPWR VPWR clkload381/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload392 clknet_leaf_13_B_in_serial_clk VGND VGND VPWR VPWR clkload392/Y sky130_fd_sc_hd__clkinv_4
XFILLER_162_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22115_ _08862_ _08863_ _08853_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_189_Right_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27972_ clknet_leaf_175_clk _01770_ net150 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_23095_ _09761_ _09762_ _09763_ VGND VGND VPWR VPWR _09764_ sky130_fd_sc_hd__a21o_1
XFILLER_192_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22046_ net65 _08819_ _08820_ systolic_inst.acc_wires\[3\]\[26\] net106 VGND VGND
+ VPWR VPWR _01772_ sky130_fd_sc_hd__a32o_1
X_26923_ clknet_leaf_6_A_in_serial_clk _00721_ net134 VGND VGND VPWR VPWR deser_A.serial_word\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_216_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_223_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_223_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_102_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_212_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29642_ clknet_leaf_31_B_in_serial_clk _03437_ net135 VGND VGND VPWR VPWR deser_B.serial_word\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_26854_ clknet_leaf_70_clk _00656_ net135 VGND VGND VPWR VPWR B_in\[126\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25805_ systolic_inst.acc_wires\[8\]\[25\] C_out\[281\] net27 VGND VGND VPWR VPWR
+ _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29573_ clknet_leaf_22_B_in_serial_clk _03368_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26785_ clknet_leaf_60_clk _00587_ net144 VGND VGND VPWR VPWR B_in\[57\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23997_ systolic_inst.B_shift\[9\]\[2\] B_in\[10\] _00008_ VGND VGND VPWR VPWR _10524_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28524_ clknet_leaf_154_clk _02322_ net150 VGND VGND VPWR VPWR ser_C.shift_reg\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25736_ systolic_inst.acc_wires\[6\]\[20\] C_out\[212\] net46 VGND VGND VPWR VPWR
+ _03038_ sky130_fd_sc_hd__mux2_1
X_13750_ B_in\[57\] deser_B.word_buffer\[57\] net89 VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__mux2_1
XFILLER_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_217_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22948_ _09590_ _09625_ systolic_inst.A_outs\[1\]\[7\] VGND VGND VPWR VPWR _09626_
+ sky130_fd_sc_hd__and3b_1
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28455_ clknet_leaf_127_clk _02253_ net144 VGND VGND VPWR VPWR ser_C.shift_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13681_ deser_B.word_buffer\[117\] deser_B.serial_word\[117\] net124 VGND VGND VPWR
+ VPWR _00518_ sky130_fd_sc_hd__mux2_1
X_25667_ systolic_inst.acc_wires\[4\]\[15\] C_out\[143\] net30 VGND VGND VPWR VPWR
+ _02969_ sky130_fd_sc_hd__mux2_1
XFILLER_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22879_ systolic_inst.B_outs\[1\]\[3\] systolic_inst.B_outs\[1\]\[4\] systolic_inst.A_outs\[1\]\[5\]
+ systolic_inst.A_outs\[1\]\[6\] VGND VGND VPWR VPWR _09559_ sky130_fd_sc_hd__and4_1
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15420_ net107 systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[4\] _12481_
+ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__a21bo_1
X_27406_ clknet_leaf_228_clk _01204_ net140 VGND VGND VPWR VPWR systolic_inst.A_outs\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_80_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24618_ net110 ser_C.shift_reg\[137\] VGND VGND VPWR VPWR _10779_ sky130_fd_sc_hd__and2_1
XFILLER_169_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28386_ clknet_leaf_32_clk _02184_ VGND VGND VPWR VPWR systolic_inst.A_shift\[18\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25598_ systolic_inst.acc_wires\[2\]\[10\] C_out\[74\] net34 VGND VGND VPWR VPWR
+ _02900_ sky130_fd_sc_hd__mux2_1
XFILLER_197_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27337_ clknet_leaf_285_clk _01135_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_15351_ _11712_ _12433_ _12434_ systolic_inst.acc_wires\[14\]\[30\] net107 VGND VGND
+ VPWR VPWR _01072_ sky130_fd_sc_hd__a32o_1
X_24549_ C_out\[101\] net99 net79 ser_C.shift_reg\[101\] _10744_ VGND VGND VPWR VPWR
+ _02351_ sky130_fd_sc_hd__a221o_1
XFILLER_200_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14302_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[7\] VGND VGND
+ VPWR VPWR _11488_ sky130_fd_sc_hd__and2b_1
XFILLER_129_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18070_ systolic_inst.B_outs\[9\]\[3\] systolic_inst.B_outs\[9\]\[4\] VGND VGND VPWR
+ VPWR _05260_ sky130_fd_sc_hd__or2_1
X_15282_ _12356_ _12361_ _12366_ _12370_ VGND VGND VPWR VPWR _12376_ sky130_fd_sc_hd__or4_1
X_27268_ clknet_leaf_268_clk _01066_ net139 VGND VGND VPWR VPWR systolic_inst.acc_wires\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29007_ clknet_leaf_104_clk _02805_ net151 VGND VGND VPWR VPWR systolic_inst.cycle_cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_17021_ systolic_inst.row_loop\[2\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[11\]\[8\]
+ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__xor2_1
X_26219_ clknet_leaf_9_A_in_serial_clk _00027_ net135 VGND VGND VPWR VPWR deser_A.word_buffer\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14233_ _11392_ _11419_ _11420_ VGND VGND VPWR VPWR _11421_ sky130_fd_sc_hd__and3_1
XFILLER_172_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27199_ clknet_leaf_262_clk _00997_ net138 VGND VGND VPWR VPWR systolic_inst.acc_wires\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_242_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_242_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14164_ _11341_ _11353_ VGND VGND VPWR VPWR _11355_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13115_ systolic_inst.B_outs\[4\]\[7\] VGND VGND VPWR VPWR _11271_ sky130_fd_sc_hd__inv_2
XFILLER_98_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14095_ deser_A.receiving deser_A.shift_reg\[1\] deser_A.shift_reg\[0\] _11304_ _11330_
+ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__a221o_1
X_18972_ _06063_ _06065_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__or3_1
XFILLER_234_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _05115_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__nor2_1
Xload_slew137 net143 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_37_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew148 net152 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_16
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_214_clk clknet_5_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_214_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17854_ _05016_ _05037_ _05039_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16805_ _04086_ _04089_ _04124_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_236_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17785_ systolic_inst.A_outs\[9\]\[0\] systolic_inst.A_outs\[8\]\[0\] net117 VGND
+ VGND VPWR VPWR _01330_ sky130_fd_sc_hd__mux2_1
XFILLER_82_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14997_ _12080_ _12082_ _12081_ VGND VGND VPWR VPWR _12117_ sky130_fd_sc_hd__o21ba_1
XFILLER_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19524_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[7\]\[18\]
+ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__or2_1
X_16736_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[7\]
+ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__o21ai_2
XFILLER_228_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13948_ deser_A.serial_word\[109\] deser_A.shift_reg\[109\] net57 VGND VGND VPWR
+ VPWR _00774_ sky130_fd_sc_hd__mux2_1
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19455_ systolic_inst.row_loop\[1\].col_loop\[3\].pe_i.prod_reg\[8\] systolic_inst.acc_wires\[7\]\[8\]
+ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__and2_1
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16667_ systolic_inst.B_outs\[11\]\[0\] systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[5\]
+ systolic_inst.A_outs\[11\]\[6\] VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__and4_1
X_13879_ deser_A.serial_word\[40\] deser_A.shift_reg\[40\] net58 VGND VGND VPWR VPWR
+ _00705_ sky130_fd_sc_hd__mux2_1
X_18406_ systolic_inst.A_outs\[8\]\[3\] systolic_inst.A_shift\[16\]\[3\] net115 VGND
+ VGND VPWR VPWR _01397_ sky130_fd_sc_hd__mux2_1
XFILLER_179_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15618_ _12672_ _12673_ VGND VGND VPWR VPWR _12674_ sky130_fd_sc_hd__and2_1
XFILLER_195_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19386_ _06374_ _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__xnor2_1
X_16598_ systolic_inst.B_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[1\] systolic_inst.A_outs\[11\]\[2\]
+ systolic_inst.B_outs\[11\]\[0\] VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a22oi_1
XFILLER_124_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18337_ _05490_ _05497_ _05498_ net60 VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__a31o_1
X_15549_ _12570_ _12571_ _12569_ VGND VGND VPWR VPWR _12607_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18268_ _05414_ _05417_ _05420_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__a211o_1
X_17219_ _04473_ _04475_ _04479_ _04480_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__nor4_1
XFILLER_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18199_ systolic_inst.row_loop\[2\].col_loop\[1\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[9\]\[0\]
+ _05379_ _05380_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__a22o_1
XFILLER_239_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20230_ systolic_inst.A_outs\[5\]\[7\] systolic_inst.A_outs\[4\]\[7\] net117 VGND
+ VGND VPWR VPWR _01593_ sky130_fd_sc_hd__mux2_1
XFILLER_190_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20161_ _07130_ _07131_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__and2_1
XFILLER_226_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20092_ _07049_ _07072_ _07062_ _07071_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_205_clk clknet_5_27__leaf_clk VGND VGND VPWR VPWR clknet_leaf_205_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_163_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23920_ systolic_inst.B_shift\[22\]\[4\] B_in\[84\] net59 VGND VGND VPWR VPWR _10493_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23851_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[24\]
+ VGND VGND VPWR VPWR _10444_ sky130_fd_sc_hd__and2_1
XFILLER_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22802_ _09479_ _09483_ VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26570_ clknet_leaf_24_A_in_serial_clk _00373_ net134 VGND VGND VPWR VPWR deser_A.shift_reg\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_232_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23782_ _11713_ _10385_ VGND VGND VPWR VPWR _10386_ sky130_fd_sc_hd__nor2_1
X_20994_ _07834_ _07867_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__and2b_1
XFILLER_77_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_225_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_241_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25521_ systolic_inst.cycle_cnt\[31\] _11279_ VGND VGND VPWR VPWR _11243_ sky130_fd_sc_hd__nand2_1
XFILLER_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22733_ _09395_ _09398_ _09416_ _09417_ VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__a211o_1
XFILLER_38_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28240_ clknet_leaf_130_clk _02038_ VGND VGND VPWR VPWR systolic_inst.B_shift\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22664_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[30\]
+ VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__or2_1
X_25452_ systolic_inst.cycle_cnt\[6\] _11306_ _11195_ systolic_inst.cycle_cnt\[7\]
+ VGND VGND VPWR VPWR _11198_ sky130_fd_sc_hd__a31o_1
XFILLER_55_1320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_240_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24403_ C_out\[28\] _11302_ net81 ser_C.shift_reg\[28\] _10671_ VGND VGND VPWR VPWR
+ _02278_ sky130_fd_sc_hd__a221o_1
X_21615_ _08417_ _08423_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28171_ clknet_leaf_80_clk _01969_ VGND VGND VPWR VPWR systolic_inst.B_shift\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22595_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[19\]
+ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25383_ systolic_inst.B_shift\[18\]\[7\] B_in\[55\] net59 VGND VGND VPWR VPWR _11161_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27122_ clknet_leaf_14_A_in_serial_clk _00920_ net143 VGND VGND VPWR VPWR deser_A.shift_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_205_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21546_ _08356_ _08357_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__and2b_1
X_24334_ _10640_ systolic_inst.A_shift\[9\]\[6\] net70 VGND VGND VPWR VPWR _02240_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Left_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24265_ systolic_inst.B_shift\[17\]\[0\] net72 _11333_ B_in\[104\] VGND VGND VPWR
+ VPWR _02202_ sky130_fd_sc_hd__a22o_1
X_27053_ clknet_leaf_27_B_in_serial_clk _00851_ net153 VGND VGND VPWR VPWR deser_B.shift_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_107_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21477_ systolic_inst.B_outs\[2\]\[5\] systolic_inst.B_shift\[2\]\[5\] systolic_inst.ce_local
+ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23216_ _09865_ _09866_ VGND VGND VPWR VPWR _09867_ sky130_fd_sc_hd__and2_1
X_26004_ systolic_inst.acc_wires\[15\]\[0\] ser_C.parallel_data\[480\] net23 VGND
+ VGND VPWR VPWR _03306_ sky130_fd_sc_hd__mux2_1
X_20428_ systolic_inst.B_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[7\] VGND VGND VPWR
+ VPWR _07364_ sky130_fd_sc_hd__nand2_4
XFILLER_175_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24196_ systolic_inst.B_shift\[22\]\[3\] net71 _11333_ B_in\[115\] VGND VGND VPWR
+ VPWR _02157_ sky130_fd_sc_hd__a22o_1
XFILLER_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_218_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_21_A_in_serial_clk clknet_2_1__leaf_A_in_serial_clk VGND VGND VPWR VPWR
+ clknet_leaf_21_A_in_serial_clk sky130_fd_sc_hd__clkbuf_8
X_23147_ _09784_ _09807_ _09797_ _09806_ VGND VGND VPWR VPWR _09808_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_136_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20359_ systolic_inst.A_outs\[5\]\[2\] systolic_inst.A_outs\[5\]\[3\] systolic_inst.B_outs\[5\]\[4\]
+ systolic_inst.B_outs\[5\]\[5\] VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__and4_1
XFILLER_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23078_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[1\]\[2\]
+ VGND VGND VPWR VPWR _09749_ sky130_fd_sc_hd__nand2_1
X_27955_ clknet_leaf_169_clk _01753_ net148 VGND VGND VPWR VPWR systolic_inst.acc_wires\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_153_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22029_ systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[3\]\[24\]
+ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_125_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ systolic_inst.A_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[2\] systolic_inst.B_outs\[14\]\[6\]
+ systolic_inst.B_outs\[14\]\[7\] VGND VGND VPWR VPWR _12042_ sky130_fd_sc_hd__and4b_1
X_26906_ clknet_leaf_17_A_in_serial_clk _00704_ net143 VGND VGND VPWR VPWR deser_A.serial_word\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27886_ clknet_leaf_309_clk _01684_ net142 VGND VGND VPWR VPWR systolic_inst.acc_wires\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_212_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29625_ clknet_leaf_8_B_in_serial_clk _03420_ net5 VGND VGND VPWR VPWR deser_B.serial_word\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26837_ clknet_leaf_88_clk _00639_ net153 VGND VGND VPWR VPWR B_in\[109\] sky130_fd_sc_hd__dfrtp_1
XFILLER_48_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14851_ systolic_inst.A_outs\[14\]\[1\] systolic_inst.B_outs\[14\]\[6\] VGND VGND
+ VPWR VPWR _11975_ sky130_fd_sc_hd__nand2_1
XFILLER_76_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13802_ B_in\[109\] deser_B.word_buffer\[109\] net88 VGND VGND VPWR VPWR _00639_
+ sky130_fd_sc_hd__mux2_1
XFILLER_112_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29556_ clknet_leaf_18_B_in_serial_clk _03351_ net144 VGND VGND VPWR VPWR deser_B.serial_word\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _04739_ _04799_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__xnor2_1
X_26768_ clknet_leaf_95_clk _00570_ net5 VGND VGND VPWR VPWR B_in\[40\] sky130_fd_sc_hd__dfrtp_1
X_14782_ _11901_ _11907_ VGND VGND VPWR VPWR _11909_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28507_ clknet_leaf_110_clk _02305_ net151 VGND VGND VPWR VPWR ser_C.shift_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16521_ _03872_ _03873_ _03874_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__or3_1
XFILLER_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_231_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13733_ B_in\[40\] deser_B.word_buffer\[40\] net90 VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25719_ systolic_inst.acc_wires\[6\]\[3\] C_out\[195\] net47 VGND VGND VPWR VPWR
+ _03021_ sky130_fd_sc_hd__mux2_1
XFILLER_72_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_231_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29487_ clknet_leaf_280_clk _03285_ net139 VGND VGND VPWR VPWR ser_C.parallel_data\[459\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_231_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26699_ clknet_leaf_6_B_in_serial_clk _00502_ net153 VGND VGND VPWR VPWR deser_B.word_buffer\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19240_ _06302_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__nor2_1
X_16452_ _03811_ _03815_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__and2_1
X_28438_ clknet_leaf_35_clk _02236_ VGND VGND VPWR VPWR systolic_inst.A_shift\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13664_ deser_B.word_buffer\[100\] deser_B.serial_word\[100\] net123 VGND VGND VPWR
+ VPWR _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_223_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15403_ systolic_inst.A_outs\[13\]\[1\] systolic_inst.B_outs\[13\]\[3\] systolic_inst.B_outs\[13\]\[4\]
+ systolic_inst.A_outs\[13\]\[0\] VGND VGND VPWR VPWR _12465_ sky130_fd_sc_hd__a22o_1
XFILLER_213_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19171_ _06208_ _06210_ _06209_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__o21bai_1
XFILLER_223_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16383_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__inv_2
X_28369_ clknet_leaf_4_clk _02167_ VGND VGND VPWR VPWR systolic_inst.A_shift\[20\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_225_Right_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13595_ deser_B.word_buffer\[31\] deser_B.serial_word\[31\] net124 VGND VGND VPWR
+ VPWR _00432_ sky130_fd_sc_hd__mux2_1
XFILLER_169_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18122_ _05257_ _05309_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_26_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15334_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[28\]
+ VGND VGND VPWR VPWR _12420_ sky130_fd_sc_hd__or2_1
XFILLER_223_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18053_ _05241_ _05242_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_229_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15265_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[16\]
+ _12358_ VGND VGND VPWR VPWR _12362_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _10520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17004_ _04308_ _04309_ _04310_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14216_ _11387_ _11389_ _11388_ VGND VGND VPWR VPWR _11404_ sky130_fd_sc_hd__o21bai_1
X_15196_ _12298_ _12301_ VGND VGND VPWR VPWR _12302_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14147_ systolic_inst.A_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[1\] systolic_inst.B_outs\[15\]\[2\]
+ systolic_inst.A_outs\[15\]\[0\] VGND VGND VPWR VPWR _11339_ sky130_fd_sc_hd__a22o_1
XFILLER_158_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14078_ deser_B.shift_reg\[112\] deser_B.shift_reg\[113\] deser_B.receiving VGND
+ VGND VPWR VPWR _00904_ sky130_fd_sc_hd__mux2_1
X_18955_ net66 _06052_ _06053_ systolic_inst.acc_wires\[8\]\[22\] net108 VGND VGND
+ VPWR VPWR _01448_ sky130_fd_sc_hd__a32o_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17906_ _05055_ _05057_ _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__a21oi_1
X_18886_ systolic_inst.row_loop\[2\].col_loop\[0\].pe_i.prod_reg\[13\] systolic_inst.acc_wires\[8\]\[13\]
+ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__nand2_1
XFILLER_6_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17837_ _05033_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_176_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17768_ systolic_inst.row_loop\[2\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[10\]\[29\]
+ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__xor2_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_235_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19507_ _06546_ _06547_ _06540_ _06544_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__o211ai_1
XFILLER_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16719_ _04003_ _04039_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__and2_1
X_17699_ _04928_ _04929_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__nand2_1
XFILLER_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19438_ _06489_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__inv_2
XFILLER_165_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19369_ _06396_ _06401_ _06427_ net119 VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__o31a_1
XFILLER_37_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21400_ _08243_ _08242_ systolic_inst.acc_wires\[4\]\[21\] _11258_ VGND VGND VPWR
+ VPWR _01703_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22380_ net122 systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[11\] _09119_
+ _09121_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__o22a_1
XFILLER_109_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21331_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[10\] systolic_inst.acc_wires\[4\]\[10\]
+ _08175_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__and3_1
XFILLER_11_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24050_ _10542_ systolic_inst.B_shift\[0\]\[4\] _11332_ VGND VGND VPWR VPWR _02054_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_867 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21262_ systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[2\] systolic_inst.acc_wires\[4\]\[2\]
+ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__and2_1
XFILLER_144_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23001_ _09676_ _09677_ VGND VGND VPWR VPWR _09678_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_165_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20213_ systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[6\]\[30\]
+ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__nand2_1
XFILLER_11_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21193_ systolic_inst.A_outs\[4\]\[6\] _07852_ _08060_ VGND VGND VPWR VPWR _08061_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_104_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20144_ net106 systolic_inst.acc_wires\[6\]\[19\] net62 _07117_ VGND VGND VPWR VPWR
+ _01573_ sky130_fd_sc_hd__a22o_1
XFILLER_172_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27740_ clknet_leaf_208_clk _01538_ net147 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[2\].pe_i.prod_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_20075_ _07054_ _07056_ _07058_ systolic_inst.acc_wires\[6\]\[9\] net106 VGND VGND
+ VPWR VPWR _01563_ sky130_fd_sc_hd__a32o_1
X_24952_ net111 ser_C.shift_reg\[304\] VGND VGND VPWR VPWR _10946_ sky130_fd_sc_hd__and2_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23903_ _10484_ systolic_inst.B_shift\[13\]\[3\] net72 VGND VGND VPWR VPWR _01965_
+ sky130_fd_sc_hd__mux2_1
X_27671_ clknet_leaf_147_clk _01469_ net149 VGND VGND VPWR VPWR systolic_inst.B_outs\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24883_ C_out\[268\] net101 net75 ser_C.shift_reg\[268\] _10911_ VGND VGND VPWR VPWR
+ _02518_ sky130_fd_sc_hd__a221o_1
XFILLER_218_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29410_ clknet_leaf_236_clk _03208_ net145 VGND VGND VPWR VPWR C_out\[382\] sky130_fd_sc_hd__dfrtp_1
X_26622_ clknet_leaf_22_B_in_serial_clk _00425_ net137 VGND VGND VPWR VPWR deser_B.word_buffer\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23834_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[0\]\[22\]
+ VGND VGND VPWR VPWR _10429_ sky130_fd_sc_hd__nand2_1
XFILLER_22_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29341_ clknet_leaf_223_clk _03139_ net149 VGND VGND VPWR VPWR C_out\[313\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26553_ clknet_leaf_26_A_in_serial_clk _00356_ net133 VGND VGND VPWR VPWR deser_A.shift_reg\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_23765_ _10363_ _10365_ _10361_ VGND VGND VPWR VPWR _10371_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_159_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ systolic_inst.A_outs\[4\]\[0\] systolic_inst.B_outs\[4\]\[7\] VGND VGND VPWR
+ VPWR _07851_ sky130_fd_sc_hd__and2b_1
XFILLER_122_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25504_ _11231_ _11232_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__nor2_1
XFILLER_207_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22716_ _11258_ systolic_inst.row_loop\[0\].col_loop\[1\].pe_i.prod_reg\[3\] VGND
+ VGND VPWR VPWR _09402_ sky130_fd_sc_hd__nand2_1
X_29272_ clknet_leaf_193_clk _03070_ net146 VGND VGND VPWR VPWR C_out\[244\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26484_ clknet_leaf_9_A_in_serial_clk _00287_ net135 VGND VGND VPWR VPWR deser_A.shift_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_214_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23696_ systolic_inst.row_loop\[0\].col_loop\[0\].pe_i.prod_reg\[1\] systolic_inst.acc_wires\[0\]\[1\]
+ VGND VGND VPWR VPWR _10312_ sky130_fd_sc_hd__or2_1
XFILLER_144_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28223_ clknet_leaf_99_clk _02021_ VGND VGND VPWR VPWR systolic_inst.B_shift\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25435_ systolic_inst.cycle_cnt\[1\] systolic_inst.cycle_cnt\[0\] VGND VGND VPWR
+ VPWR _11187_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22647_ net109 systolic_inst.acc_wires\[2\]\[27\] net65 _09356_ VGND VGND VPWR VPWR
+ _01837_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28154_ clknet_leaf_102_clk _01952_ net151 VGND VGND VPWR VPWR systolic_inst.acc_wires\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_220_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13380_ A_in\[89\] deser_A.word_buffer\[89\] net95 VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__mux2_1
X_22578_ systolic_inst.row_loop\[0\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[2\]\[16\]
+ VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__xnor2_1
X_25366_ net112 ser_C.shift_reg\[511\] VGND VGND VPWR VPWR _11153_ sky130_fd_sc_hd__and2_1
XFILLER_222_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27105_ clknet_leaf_10_B_in_serial_clk _00903_ net144 VGND VGND VPWR VPWR deser_B.shift_reg\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24317_ systolic_inst.A_shift\[11\]\[6\] A_in\[46\] net59 VGND VGND VPWR VPWR _10632_
+ sky130_fd_sc_hd__mux2_1
X_28085_ clknet_leaf_120_clk _01883_ net149 VGND VGND VPWR VPWR systolic_inst.acc_wires\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_21529_ _08322_ _08338_ _08340_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__and3_1
XFILLER_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25297_ ser_C.parallel_data\[475\] net102 net74 ser_C.shift_reg\[475\] _11118_ VGND
+ VGND VPWR VPWR _02725_ sky130_fd_sc_hd__a221o_1
XFILLER_182_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27036_ clknet_leaf_14_B_in_serial_clk _00834_ net5 VGND VGND VPWR VPWR deser_B.shift_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15050_ _12167_ _12168_ VGND VGND VPWR VPWR _12169_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24248_ _10609_ systolic_inst.A_shift\[18\]\[7\] net70 VGND VGND VPWR VPWR _02185_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_224_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14001_ deser_B.shift_reg\[35\] deser_B.shift_reg\[36\] deser_B.receiving VGND VGND
+ VPWR VPWR _00827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_224_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24179_ systolic_inst.A_shift\[25\]\[2\] net70 _10505_ systolic_inst.A_shift\[26\]\[2\]
+ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__a22o_1
XFILLER_107_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28987_ clknet_leaf_24_clk _02785_ VGND VGND VPWR VPWR systolic_inst.A_shift\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_231_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18740_ systolic_inst.B_outs\[8\]\[6\] systolic_inst.A_outs\[8\]\[7\] VGND VGND VPWR
+ VPWR _05864_ sky130_fd_sc_hd__nand2_1
X_27938_ clknet_leaf_171_clk _01736_ net148 VGND VGND VPWR VPWR systolic_inst.row_loop\[0\].col_loop\[3\].pe_i.prod_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15952_ _12968_ _12971_ VGND VGND VPWR VPWR _12972_ sky130_fd_sc_hd__nand2_1
XFILLER_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14903_ _11985_ _11988_ _12024_ net118 VGND VGND VPWR VPWR _12026_ sky130_fd_sc_hd__o31a_1
XFILLER_62_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18671_ _05794_ _05795_ _05796_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__and3_1
X_15883_ systolic_inst.row_loop\[3\].col_loop\[1\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[13\]\[20\]
+ VGND VGND VPWR VPWR _12913_ sky130_fd_sc_hd__nand2_1
X_27869_ clknet_leaf_310_clk _01667_ net137 VGND VGND VPWR VPWR systolic_inst.row_loop\[1\].col_loop\[0\].pe_i.prod_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_236_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17622_ _04857_ _04858_ _04856_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__a21bo_1
X_29608_ clknet_leaf_24_B_in_serial_clk _03403_ net143 VGND VGND VPWR VPWR deser_B.serial_word\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14834_ _11958_ _11957_ VGND VGND VPWR VPWR _11959_ sky130_fd_sc_hd__nand2b_1
XFILLER_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29539_ clknet_leaf_246_clk _03337_ net145 VGND VGND VPWR VPWR ser_C.parallel_data\[511\]
+ sky130_fd_sc_hd__dfrtp_1
X_17553_ _04802_ _04803_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_218_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ systolic_inst.B_outs\[14\]\[0\] systolic_inst.B_outs\[14\]\[1\] systolic_inst.A_outs\[14\]\[1\]
+ systolic_inst.A_outs\[14\]\[2\] VGND VGND VPWR VPWR _11893_ sky130_fd_sc_hd__and4_1
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16504_ _03852_ _03857_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__nor2_1
X_13716_ B_in\[23\] deser_B.word_buffer\[23\] net86 VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17484_ net105 _04736_ _04737_ _04707_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__o31a_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14696_ _11843_ _11845_ _11848_ VGND VGND VPWR VPWR _11850_ sky130_fd_sc_hd__a21oi_2
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19223_ _06248_ _06250_ _06249_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__o21ba_1
XFILLER_176_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16435_ systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[11\] systolic_inst.acc_wires\[12\]\[11\]
+ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__or2_1
XFILLER_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13647_ deser_B.word_buffer\[83\] deser_B.serial_word\[83\] net124 VGND VGND VPWR
+ VPWR _00484_ sky130_fd_sc_hd__mux2_1
XFILLER_220_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19154_ _06212_ _06218_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_15_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16366_ net115 systolic_inst.row_loop\[3\].col_loop\[0\].pe_i.prod_reg\[0\] systolic_inst.acc_wires\[12\]\[0\]
+ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__a21oi_1
X_13578_ deser_B.word_buffer\[14\] deser_B.serial_word\[14\] net124 VGND VGND VPWR
+ VPWR _00415_ sky130_fd_sc_hd__mux2_1
XFILLER_121_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18105_ systolic_inst.A_outs\[9\]\[5\] systolic_inst.B_outs\[9\]\[6\] systolic_inst.A_outs\[9\]\[6\]
+ systolic_inst.B_outs\[9\]\[7\] VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__and4b_1
X_15317_ _12401_ _12403_ _12405_ VGND VGND VPWR VPWR _12406_ sky130_fd_sc_hd__or3_1
X_19085_ systolic_inst.A_outs\[7\]\[2\] systolic_inst.B_outs\[7\]\[3\] systolic_inst.B_outs\[7\]\[4\]
+ systolic_inst.A_outs\[7\]\[1\] VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__a22o_1
XFILLER_185_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16297_ _03627_ _03677_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__and2b_1
XFILLER_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18036_ systolic_inst.B_outs\[9\]\[5\] systolic_inst.A_outs\[9\]\[5\] VGND VGND VPWR
+ VPWR _05227_ sky130_fd_sc_hd__nand2_1
X_15248_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[15\] systolic_inst.acc_wires\[14\]\[15\]
+ VGND VGND VPWR VPWR _12347_ sky130_fd_sc_hd__nor2_1
XFILLER_172_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15179_ systolic_inst.row_loop\[3\].col_loop\[2\].pe_i.prod_reg\[5\] systolic_inst.acc_wires\[14\]\[5\]
+ VGND VGND VPWR VPWR _12288_ sky130_fd_sc_hd__or2_1
XFILLER_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19987_ _06895_ _06980_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__nand2_1
XFILLER_141_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18938_ _06014_ _06038_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__nor2_1
XFILLER_80_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

