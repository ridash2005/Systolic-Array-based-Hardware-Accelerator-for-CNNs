module Systolic4x4_serial_io (A_in_frame_sync,
    A_in_serial_clk,
    A_in_serial_data,
    B_in_frame_sync,
    B_in_serial_clk,
    B_in_serial_data,
    C_out_frame_sync,
    C_out_serial_clk,
    C_out_serial_data,
    clk,
    done,
    rst_n,
    start);
 input A_in_frame_sync;
 input A_in_serial_clk;
 input A_in_serial_data;
 input B_in_frame_sync;
 input B_in_serial_clk;
 input B_in_serial_data;
 output C_out_frame_sync;
 output C_out_serial_clk;
 output C_out_serial_data;
 input clk;
 output done;
 input rst_n;
 input start;

 wire \A_in[0] ;
 wire \A_in[100] ;
 wire \A_in[101] ;
 wire \A_in[102] ;
 wire \A_in[103] ;
 wire \A_in[104] ;
 wire \A_in[105] ;
 wire \A_in[106] ;
 wire \A_in[107] ;
 wire \A_in[108] ;
 wire \A_in[109] ;
 wire \A_in[10] ;
 wire \A_in[110] ;
 wire \A_in[111] ;
 wire \A_in[112] ;
 wire \A_in[113] ;
 wire \A_in[114] ;
 wire \A_in[115] ;
 wire \A_in[116] ;
 wire \A_in[117] ;
 wire \A_in[118] ;
 wire \A_in[119] ;
 wire \A_in[11] ;
 wire \A_in[120] ;
 wire \A_in[121] ;
 wire \A_in[122] ;
 wire \A_in[123] ;
 wire \A_in[124] ;
 wire \A_in[125] ;
 wire \A_in[126] ;
 wire \A_in[127] ;
 wire \A_in[12] ;
 wire \A_in[13] ;
 wire \A_in[14] ;
 wire \A_in[15] ;
 wire \A_in[16] ;
 wire \A_in[17] ;
 wire \A_in[18] ;
 wire \A_in[19] ;
 wire \A_in[1] ;
 wire \A_in[20] ;
 wire \A_in[21] ;
 wire \A_in[22] ;
 wire \A_in[23] ;
 wire \A_in[24] ;
 wire \A_in[25] ;
 wire \A_in[26] ;
 wire \A_in[27] ;
 wire \A_in[28] ;
 wire \A_in[29] ;
 wire \A_in[2] ;
 wire \A_in[30] ;
 wire \A_in[31] ;
 wire \A_in[32] ;
 wire \A_in[33] ;
 wire \A_in[34] ;
 wire \A_in[35] ;
 wire \A_in[36] ;
 wire \A_in[37] ;
 wire \A_in[38] ;
 wire \A_in[39] ;
 wire \A_in[3] ;
 wire \A_in[40] ;
 wire \A_in[41] ;
 wire \A_in[42] ;
 wire \A_in[43] ;
 wire \A_in[44] ;
 wire \A_in[45] ;
 wire \A_in[46] ;
 wire \A_in[47] ;
 wire \A_in[48] ;
 wire \A_in[49] ;
 wire \A_in[4] ;
 wire \A_in[50] ;
 wire \A_in[51] ;
 wire \A_in[52] ;
 wire \A_in[53] ;
 wire \A_in[54] ;
 wire \A_in[55] ;
 wire \A_in[56] ;
 wire \A_in[57] ;
 wire \A_in[58] ;
 wire \A_in[59] ;
 wire \A_in[5] ;
 wire \A_in[60] ;
 wire \A_in[61] ;
 wire \A_in[62] ;
 wire \A_in[63] ;
 wire \A_in[64] ;
 wire \A_in[65] ;
 wire \A_in[66] ;
 wire \A_in[67] ;
 wire \A_in[68] ;
 wire \A_in[69] ;
 wire \A_in[6] ;
 wire \A_in[70] ;
 wire \A_in[71] ;
 wire \A_in[72] ;
 wire \A_in[73] ;
 wire \A_in[74] ;
 wire \A_in[75] ;
 wire \A_in[76] ;
 wire \A_in[77] ;
 wire \A_in[78] ;
 wire \A_in[79] ;
 wire \A_in[7] ;
 wire \A_in[80] ;
 wire \A_in[81] ;
 wire \A_in[82] ;
 wire \A_in[83] ;
 wire \A_in[84] ;
 wire \A_in[85] ;
 wire \A_in[86] ;
 wire \A_in[87] ;
 wire \A_in[88] ;
 wire \A_in[89] ;
 wire \A_in[8] ;
 wire \A_in[90] ;
 wire \A_in[91] ;
 wire \A_in[92] ;
 wire \A_in[93] ;
 wire \A_in[94] ;
 wire \A_in[95] ;
 wire \A_in[96] ;
 wire \A_in[97] ;
 wire \A_in[98] ;
 wire \A_in[99] ;
 wire \A_in[9] ;
 wire A_in_valid;
 wire \B_in[0] ;
 wire \B_in[100] ;
 wire \B_in[101] ;
 wire \B_in[102] ;
 wire \B_in[103] ;
 wire \B_in[104] ;
 wire \B_in[105] ;
 wire \B_in[106] ;
 wire \B_in[107] ;
 wire \B_in[108] ;
 wire \B_in[109] ;
 wire \B_in[10] ;
 wire \B_in[110] ;
 wire \B_in[111] ;
 wire \B_in[112] ;
 wire \B_in[113] ;
 wire \B_in[114] ;
 wire \B_in[115] ;
 wire \B_in[116] ;
 wire \B_in[117] ;
 wire \B_in[118] ;
 wire \B_in[119] ;
 wire \B_in[11] ;
 wire \B_in[120] ;
 wire \B_in[121] ;
 wire \B_in[122] ;
 wire \B_in[123] ;
 wire \B_in[124] ;
 wire \B_in[125] ;
 wire \B_in[126] ;
 wire \B_in[127] ;
 wire \B_in[12] ;
 wire \B_in[13] ;
 wire \B_in[14] ;
 wire \B_in[15] ;
 wire \B_in[16] ;
 wire \B_in[17] ;
 wire \B_in[18] ;
 wire \B_in[19] ;
 wire \B_in[1] ;
 wire \B_in[20] ;
 wire \B_in[21] ;
 wire \B_in[22] ;
 wire \B_in[23] ;
 wire \B_in[24] ;
 wire \B_in[25] ;
 wire \B_in[26] ;
 wire \B_in[27] ;
 wire \B_in[28] ;
 wire \B_in[29] ;
 wire \B_in[2] ;
 wire \B_in[30] ;
 wire \B_in[31] ;
 wire \B_in[32] ;
 wire \B_in[33] ;
 wire \B_in[34] ;
 wire \B_in[35] ;
 wire \B_in[36] ;
 wire \B_in[37] ;
 wire \B_in[38] ;
 wire \B_in[39] ;
 wire \B_in[3] ;
 wire \B_in[40] ;
 wire \B_in[41] ;
 wire \B_in[42] ;
 wire \B_in[43] ;
 wire \B_in[44] ;
 wire \B_in[45] ;
 wire \B_in[46] ;
 wire \B_in[47] ;
 wire \B_in[48] ;
 wire \B_in[49] ;
 wire \B_in[4] ;
 wire \B_in[50] ;
 wire \B_in[51] ;
 wire \B_in[52] ;
 wire \B_in[53] ;
 wire \B_in[54] ;
 wire \B_in[55] ;
 wire \B_in[56] ;
 wire \B_in[57] ;
 wire \B_in[58] ;
 wire \B_in[59] ;
 wire \B_in[5] ;
 wire \B_in[60] ;
 wire \B_in[61] ;
 wire \B_in[62] ;
 wire \B_in[63] ;
 wire \B_in[64] ;
 wire \B_in[65] ;
 wire \B_in[66] ;
 wire \B_in[67] ;
 wire \B_in[68] ;
 wire \B_in[69] ;
 wire \B_in[6] ;
 wire \B_in[70] ;
 wire \B_in[71] ;
 wire \B_in[72] ;
 wire \B_in[73] ;
 wire \B_in[74] ;
 wire \B_in[75] ;
 wire \B_in[76] ;
 wire \B_in[77] ;
 wire \B_in[78] ;
 wire \B_in[79] ;
 wire \B_in[7] ;
 wire \B_in[80] ;
 wire \B_in[81] ;
 wire \B_in[82] ;
 wire \B_in[83] ;
 wire \B_in[84] ;
 wire \B_in[85] ;
 wire \B_in[86] ;
 wire \B_in[87] ;
 wire \B_in[88] ;
 wire \B_in[89] ;
 wire \B_in[8] ;
 wire \B_in[90] ;
 wire \B_in[91] ;
 wire \B_in[92] ;
 wire \B_in[93] ;
 wire \B_in[94] ;
 wire \B_in[95] ;
 wire \B_in[96] ;
 wire \B_in[97] ;
 wire \B_in[98] ;
 wire \B_in[99] ;
 wire \B_in[9] ;
 wire B_in_valid;
 wire \C_out[0] ;
 wire \C_out[100] ;
 wire \C_out[101] ;
 wire \C_out[102] ;
 wire \C_out[103] ;
 wire \C_out[104] ;
 wire \C_out[105] ;
 wire \C_out[106] ;
 wire \C_out[107] ;
 wire \C_out[108] ;
 wire \C_out[109] ;
 wire \C_out[10] ;
 wire \C_out[110] ;
 wire \C_out[111] ;
 wire \C_out[112] ;
 wire \C_out[113] ;
 wire \C_out[114] ;
 wire \C_out[115] ;
 wire \C_out[116] ;
 wire \C_out[117] ;
 wire \C_out[118] ;
 wire \C_out[119] ;
 wire \C_out[11] ;
 wire \C_out[120] ;
 wire \C_out[121] ;
 wire \C_out[122] ;
 wire \C_out[123] ;
 wire \C_out[124] ;
 wire \C_out[125] ;
 wire \C_out[126] ;
 wire \C_out[127] ;
 wire \C_out[128] ;
 wire \C_out[129] ;
 wire \C_out[12] ;
 wire \C_out[130] ;
 wire \C_out[131] ;
 wire \C_out[132] ;
 wire \C_out[133] ;
 wire \C_out[134] ;
 wire \C_out[135] ;
 wire \C_out[136] ;
 wire \C_out[137] ;
 wire \C_out[138] ;
 wire \C_out[139] ;
 wire \C_out[13] ;
 wire \C_out[140] ;
 wire \C_out[141] ;
 wire \C_out[142] ;
 wire \C_out[143] ;
 wire \C_out[144] ;
 wire \C_out[145] ;
 wire \C_out[146] ;
 wire \C_out[147] ;
 wire \C_out[148] ;
 wire \C_out[149] ;
 wire \C_out[14] ;
 wire \C_out[150] ;
 wire \C_out[151] ;
 wire \C_out[152] ;
 wire \C_out[153] ;
 wire \C_out[154] ;
 wire \C_out[155] ;
 wire \C_out[156] ;
 wire \C_out[157] ;
 wire \C_out[158] ;
 wire \C_out[159] ;
 wire \C_out[15] ;
 wire \C_out[160] ;
 wire \C_out[161] ;
 wire \C_out[162] ;
 wire \C_out[163] ;
 wire \C_out[164] ;
 wire \C_out[165] ;
 wire \C_out[166] ;
 wire \C_out[167] ;
 wire \C_out[168] ;
 wire \C_out[169] ;
 wire \C_out[16] ;
 wire \C_out[170] ;
 wire \C_out[171] ;
 wire \C_out[172] ;
 wire \C_out[173] ;
 wire \C_out[174] ;
 wire \C_out[175] ;
 wire \C_out[176] ;
 wire \C_out[177] ;
 wire \C_out[178] ;
 wire \C_out[179] ;
 wire \C_out[17] ;
 wire \C_out[180] ;
 wire \C_out[181] ;
 wire \C_out[182] ;
 wire \C_out[183] ;
 wire \C_out[184] ;
 wire \C_out[185] ;
 wire \C_out[186] ;
 wire \C_out[187] ;
 wire \C_out[188] ;
 wire \C_out[189] ;
 wire \C_out[18] ;
 wire \C_out[190] ;
 wire \C_out[191] ;
 wire \C_out[192] ;
 wire \C_out[193] ;
 wire \C_out[194] ;
 wire \C_out[195] ;
 wire \C_out[196] ;
 wire \C_out[197] ;
 wire \C_out[198] ;
 wire \C_out[199] ;
 wire \C_out[19] ;
 wire \C_out[1] ;
 wire \C_out[200] ;
 wire \C_out[201] ;
 wire \C_out[202] ;
 wire \C_out[203] ;
 wire \C_out[204] ;
 wire \C_out[205] ;
 wire \C_out[206] ;
 wire \C_out[207] ;
 wire \C_out[208] ;
 wire \C_out[209] ;
 wire \C_out[20] ;
 wire \C_out[210] ;
 wire \C_out[211] ;
 wire \C_out[212] ;
 wire \C_out[213] ;
 wire \C_out[214] ;
 wire \C_out[215] ;
 wire \C_out[216] ;
 wire \C_out[217] ;
 wire \C_out[218] ;
 wire \C_out[219] ;
 wire \C_out[21] ;
 wire \C_out[220] ;
 wire \C_out[221] ;
 wire \C_out[222] ;
 wire \C_out[223] ;
 wire \C_out[224] ;
 wire \C_out[225] ;
 wire \C_out[226] ;
 wire \C_out[227] ;
 wire \C_out[228] ;
 wire \C_out[229] ;
 wire \C_out[22] ;
 wire \C_out[230] ;
 wire \C_out[231] ;
 wire \C_out[232] ;
 wire \C_out[233] ;
 wire \C_out[234] ;
 wire \C_out[235] ;
 wire \C_out[236] ;
 wire \C_out[237] ;
 wire \C_out[238] ;
 wire \C_out[239] ;
 wire \C_out[23] ;
 wire \C_out[240] ;
 wire \C_out[241] ;
 wire \C_out[242] ;
 wire \C_out[243] ;
 wire \C_out[244] ;
 wire \C_out[245] ;
 wire \C_out[246] ;
 wire \C_out[247] ;
 wire \C_out[248] ;
 wire \C_out[249] ;
 wire \C_out[24] ;
 wire \C_out[250] ;
 wire \C_out[251] ;
 wire \C_out[252] ;
 wire \C_out[253] ;
 wire \C_out[254] ;
 wire \C_out[255] ;
 wire \C_out[256] ;
 wire \C_out[257] ;
 wire \C_out[258] ;
 wire \C_out[259] ;
 wire \C_out[25] ;
 wire \C_out[260] ;
 wire \C_out[261] ;
 wire \C_out[262] ;
 wire \C_out[263] ;
 wire \C_out[264] ;
 wire \C_out[265] ;
 wire \C_out[266] ;
 wire \C_out[267] ;
 wire \C_out[268] ;
 wire \C_out[269] ;
 wire \C_out[26] ;
 wire \C_out[270] ;
 wire \C_out[271] ;
 wire \C_out[272] ;
 wire \C_out[273] ;
 wire \C_out[274] ;
 wire \C_out[275] ;
 wire \C_out[276] ;
 wire \C_out[277] ;
 wire \C_out[278] ;
 wire \C_out[279] ;
 wire \C_out[27] ;
 wire \C_out[280] ;
 wire \C_out[281] ;
 wire \C_out[282] ;
 wire \C_out[283] ;
 wire \C_out[284] ;
 wire \C_out[285] ;
 wire \C_out[286] ;
 wire \C_out[287] ;
 wire \C_out[288] ;
 wire \C_out[289] ;
 wire \C_out[28] ;
 wire \C_out[290] ;
 wire \C_out[291] ;
 wire \C_out[292] ;
 wire \C_out[293] ;
 wire \C_out[294] ;
 wire \C_out[295] ;
 wire \C_out[296] ;
 wire \C_out[297] ;
 wire \C_out[298] ;
 wire \C_out[299] ;
 wire \C_out[29] ;
 wire \C_out[2] ;
 wire \C_out[300] ;
 wire \C_out[301] ;
 wire \C_out[302] ;
 wire \C_out[303] ;
 wire \C_out[304] ;
 wire \C_out[305] ;
 wire \C_out[306] ;
 wire \C_out[307] ;
 wire \C_out[308] ;
 wire \C_out[309] ;
 wire \C_out[30] ;
 wire \C_out[310] ;
 wire \C_out[311] ;
 wire \C_out[312] ;
 wire \C_out[313] ;
 wire \C_out[314] ;
 wire \C_out[315] ;
 wire \C_out[316] ;
 wire \C_out[317] ;
 wire \C_out[318] ;
 wire \C_out[319] ;
 wire \C_out[31] ;
 wire \C_out[320] ;
 wire \C_out[321] ;
 wire \C_out[322] ;
 wire \C_out[323] ;
 wire \C_out[324] ;
 wire \C_out[325] ;
 wire \C_out[326] ;
 wire \C_out[327] ;
 wire \C_out[328] ;
 wire \C_out[329] ;
 wire \C_out[32] ;
 wire \C_out[330] ;
 wire \C_out[331] ;
 wire \C_out[332] ;
 wire \C_out[333] ;
 wire \C_out[334] ;
 wire \C_out[335] ;
 wire \C_out[336] ;
 wire \C_out[337] ;
 wire \C_out[338] ;
 wire \C_out[339] ;
 wire \C_out[33] ;
 wire \C_out[340] ;
 wire \C_out[341] ;
 wire \C_out[342] ;
 wire \C_out[343] ;
 wire \C_out[344] ;
 wire \C_out[345] ;
 wire \C_out[346] ;
 wire \C_out[347] ;
 wire \C_out[348] ;
 wire \C_out[349] ;
 wire \C_out[34] ;
 wire \C_out[350] ;
 wire \C_out[351] ;
 wire \C_out[352] ;
 wire \C_out[353] ;
 wire \C_out[354] ;
 wire \C_out[355] ;
 wire \C_out[356] ;
 wire \C_out[357] ;
 wire \C_out[358] ;
 wire \C_out[359] ;
 wire \C_out[35] ;
 wire \C_out[360] ;
 wire \C_out[361] ;
 wire \C_out[362] ;
 wire \C_out[363] ;
 wire \C_out[364] ;
 wire \C_out[365] ;
 wire \C_out[366] ;
 wire \C_out[367] ;
 wire \C_out[368] ;
 wire \C_out[369] ;
 wire \C_out[36] ;
 wire \C_out[370] ;
 wire \C_out[371] ;
 wire \C_out[372] ;
 wire \C_out[373] ;
 wire \C_out[374] ;
 wire \C_out[375] ;
 wire \C_out[376] ;
 wire \C_out[377] ;
 wire \C_out[378] ;
 wire \C_out[379] ;
 wire \C_out[37] ;
 wire \C_out[380] ;
 wire \C_out[381] ;
 wire \C_out[382] ;
 wire \C_out[383] ;
 wire \C_out[384] ;
 wire \C_out[385] ;
 wire \C_out[386] ;
 wire \C_out[387] ;
 wire \C_out[388] ;
 wire \C_out[389] ;
 wire \C_out[38] ;
 wire \C_out[390] ;
 wire \C_out[391] ;
 wire \C_out[392] ;
 wire \C_out[393] ;
 wire \C_out[394] ;
 wire \C_out[395] ;
 wire \C_out[396] ;
 wire \C_out[397] ;
 wire \C_out[398] ;
 wire \C_out[399] ;
 wire \C_out[39] ;
 wire \C_out[3] ;
 wire \C_out[400] ;
 wire \C_out[401] ;
 wire \C_out[402] ;
 wire \C_out[403] ;
 wire \C_out[404] ;
 wire \C_out[405] ;
 wire \C_out[406] ;
 wire \C_out[407] ;
 wire \C_out[408] ;
 wire \C_out[409] ;
 wire \C_out[40] ;
 wire \C_out[410] ;
 wire \C_out[411] ;
 wire \C_out[412] ;
 wire \C_out[413] ;
 wire \C_out[414] ;
 wire \C_out[415] ;
 wire \C_out[416] ;
 wire \C_out[417] ;
 wire \C_out[418] ;
 wire \C_out[419] ;
 wire \C_out[41] ;
 wire \C_out[420] ;
 wire \C_out[421] ;
 wire \C_out[422] ;
 wire \C_out[423] ;
 wire \C_out[424] ;
 wire \C_out[425] ;
 wire \C_out[426] ;
 wire \C_out[427] ;
 wire \C_out[428] ;
 wire \C_out[429] ;
 wire \C_out[42] ;
 wire \C_out[430] ;
 wire \C_out[431] ;
 wire \C_out[432] ;
 wire \C_out[433] ;
 wire \C_out[434] ;
 wire \C_out[435] ;
 wire \C_out[436] ;
 wire \C_out[437] ;
 wire \C_out[438] ;
 wire \C_out[439] ;
 wire \C_out[43] ;
 wire \C_out[44] ;
 wire \C_out[45] ;
 wire \C_out[46] ;
 wire \C_out[47] ;
 wire \C_out[48] ;
 wire \C_out[49] ;
 wire \C_out[4] ;
 wire \C_out[50] ;
 wire \C_out[51] ;
 wire \C_out[52] ;
 wire \C_out[53] ;
 wire \C_out[54] ;
 wire \C_out[55] ;
 wire \C_out[56] ;
 wire \C_out[57] ;
 wire \C_out[58] ;
 wire \C_out[59] ;
 wire \C_out[5] ;
 wire \C_out[60] ;
 wire \C_out[61] ;
 wire \C_out[62] ;
 wire \C_out[63] ;
 wire \C_out[64] ;
 wire \C_out[65] ;
 wire \C_out[66] ;
 wire \C_out[67] ;
 wire \C_out[68] ;
 wire \C_out[69] ;
 wire \C_out[6] ;
 wire \C_out[70] ;
 wire \C_out[71] ;
 wire \C_out[72] ;
 wire \C_out[73] ;
 wire \C_out[74] ;
 wire \C_out[75] ;
 wire \C_out[76] ;
 wire \C_out[77] ;
 wire \C_out[78] ;
 wire \C_out[79] ;
 wire \C_out[7] ;
 wire \C_out[80] ;
 wire \C_out[81] ;
 wire \C_out[82] ;
 wire \C_out[83] ;
 wire \C_out[84] ;
 wire \C_out[85] ;
 wire \C_out[86] ;
 wire \C_out[87] ;
 wire \C_out[88] ;
 wire \C_out[89] ;
 wire \C_out[8] ;
 wire \C_out[90] ;
 wire \C_out[91] ;
 wire \C_out[92] ;
 wire \C_out[93] ;
 wire \C_out[94] ;
 wire \C_out[95] ;
 wire \C_out[96] ;
 wire \C_out[97] ;
 wire \C_out[98] ;
 wire \C_out[99] ;
 wire \C_out[9] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire \deser_A.bit_idx[0] ;
 wire \deser_A.bit_idx[1] ;
 wire \deser_A.bit_idx[2] ;
 wire \deser_A.bit_idx[3] ;
 wire \deser_A.bit_idx[4] ;
 wire \deser_A.bit_idx[5] ;
 wire \deser_A.bit_idx[6] ;
 wire \deser_A.receiving ;
 wire \deser_A.serial_toggle ;
 wire \deser_A.serial_toggle_sync1 ;
 wire \deser_A.serial_toggle_sync2 ;
 wire \deser_A.serial_word[0] ;
 wire \deser_A.serial_word[100] ;
 wire \deser_A.serial_word[101] ;
 wire \deser_A.serial_word[102] ;
 wire \deser_A.serial_word[103] ;
 wire \deser_A.serial_word[104] ;
 wire \deser_A.serial_word[105] ;
 wire \deser_A.serial_word[106] ;
 wire \deser_A.serial_word[107] ;
 wire \deser_A.serial_word[108] ;
 wire \deser_A.serial_word[109] ;
 wire \deser_A.serial_word[10] ;
 wire \deser_A.serial_word[110] ;
 wire \deser_A.serial_word[111] ;
 wire \deser_A.serial_word[112] ;
 wire \deser_A.serial_word[113] ;
 wire \deser_A.serial_word[114] ;
 wire \deser_A.serial_word[115] ;
 wire \deser_A.serial_word[116] ;
 wire \deser_A.serial_word[117] ;
 wire \deser_A.serial_word[118] ;
 wire \deser_A.serial_word[119] ;
 wire \deser_A.serial_word[11] ;
 wire \deser_A.serial_word[120] ;
 wire \deser_A.serial_word[121] ;
 wire \deser_A.serial_word[122] ;
 wire \deser_A.serial_word[123] ;
 wire \deser_A.serial_word[124] ;
 wire \deser_A.serial_word[125] ;
 wire \deser_A.serial_word[126] ;
 wire \deser_A.serial_word[127] ;
 wire \deser_A.serial_word[12] ;
 wire \deser_A.serial_word[13] ;
 wire \deser_A.serial_word[14] ;
 wire \deser_A.serial_word[15] ;
 wire \deser_A.serial_word[16] ;
 wire \deser_A.serial_word[17] ;
 wire \deser_A.serial_word[18] ;
 wire \deser_A.serial_word[19] ;
 wire \deser_A.serial_word[1] ;
 wire \deser_A.serial_word[20] ;
 wire \deser_A.serial_word[21] ;
 wire \deser_A.serial_word[22] ;
 wire \deser_A.serial_word[23] ;
 wire \deser_A.serial_word[24] ;
 wire \deser_A.serial_word[25] ;
 wire \deser_A.serial_word[26] ;
 wire \deser_A.serial_word[27] ;
 wire \deser_A.serial_word[28] ;
 wire \deser_A.serial_word[29] ;
 wire \deser_A.serial_word[2] ;
 wire \deser_A.serial_word[30] ;
 wire \deser_A.serial_word[31] ;
 wire \deser_A.serial_word[32] ;
 wire \deser_A.serial_word[33] ;
 wire \deser_A.serial_word[34] ;
 wire \deser_A.serial_word[35] ;
 wire \deser_A.serial_word[36] ;
 wire \deser_A.serial_word[37] ;
 wire \deser_A.serial_word[38] ;
 wire \deser_A.serial_word[39] ;
 wire \deser_A.serial_word[3] ;
 wire \deser_A.serial_word[40] ;
 wire \deser_A.serial_word[41] ;
 wire \deser_A.serial_word[42] ;
 wire \deser_A.serial_word[43] ;
 wire \deser_A.serial_word[44] ;
 wire \deser_A.serial_word[45] ;
 wire \deser_A.serial_word[46] ;
 wire \deser_A.serial_word[47] ;
 wire \deser_A.serial_word[48] ;
 wire \deser_A.serial_word[49] ;
 wire \deser_A.serial_word[4] ;
 wire \deser_A.serial_word[50] ;
 wire \deser_A.serial_word[51] ;
 wire \deser_A.serial_word[52] ;
 wire \deser_A.serial_word[53] ;
 wire \deser_A.serial_word[54] ;
 wire \deser_A.serial_word[55] ;
 wire \deser_A.serial_word[56] ;
 wire \deser_A.serial_word[57] ;
 wire \deser_A.serial_word[58] ;
 wire \deser_A.serial_word[59] ;
 wire \deser_A.serial_word[5] ;
 wire \deser_A.serial_word[60] ;
 wire \deser_A.serial_word[61] ;
 wire \deser_A.serial_word[62] ;
 wire \deser_A.serial_word[63] ;
 wire \deser_A.serial_word[64] ;
 wire \deser_A.serial_word[65] ;
 wire \deser_A.serial_word[66] ;
 wire \deser_A.serial_word[67] ;
 wire \deser_A.serial_word[68] ;
 wire \deser_A.serial_word[69] ;
 wire \deser_A.serial_word[6] ;
 wire \deser_A.serial_word[70] ;
 wire \deser_A.serial_word[71] ;
 wire \deser_A.serial_word[72] ;
 wire \deser_A.serial_word[73] ;
 wire \deser_A.serial_word[74] ;
 wire \deser_A.serial_word[75] ;
 wire \deser_A.serial_word[76] ;
 wire \deser_A.serial_word[77] ;
 wire \deser_A.serial_word[78] ;
 wire \deser_A.serial_word[79] ;
 wire \deser_A.serial_word[7] ;
 wire \deser_A.serial_word[80] ;
 wire \deser_A.serial_word[81] ;
 wire \deser_A.serial_word[82] ;
 wire \deser_A.serial_word[83] ;
 wire \deser_A.serial_word[84] ;
 wire \deser_A.serial_word[85] ;
 wire \deser_A.serial_word[86] ;
 wire \deser_A.serial_word[87] ;
 wire \deser_A.serial_word[88] ;
 wire \deser_A.serial_word[89] ;
 wire \deser_A.serial_word[8] ;
 wire \deser_A.serial_word[90] ;
 wire \deser_A.serial_word[91] ;
 wire \deser_A.serial_word[92] ;
 wire \deser_A.serial_word[93] ;
 wire \deser_A.serial_word[94] ;
 wire \deser_A.serial_word[95] ;
 wire \deser_A.serial_word[96] ;
 wire \deser_A.serial_word[97] ;
 wire \deser_A.serial_word[98] ;
 wire \deser_A.serial_word[99] ;
 wire \deser_A.serial_word[9] ;
 wire \deser_A.serial_word_ready ;
 wire \deser_A.shift_reg[0] ;
 wire \deser_A.shift_reg[100] ;
 wire \deser_A.shift_reg[101] ;
 wire \deser_A.shift_reg[102] ;
 wire \deser_A.shift_reg[103] ;
 wire \deser_A.shift_reg[104] ;
 wire \deser_A.shift_reg[105] ;
 wire \deser_A.shift_reg[106] ;
 wire \deser_A.shift_reg[107] ;
 wire \deser_A.shift_reg[108] ;
 wire \deser_A.shift_reg[109] ;
 wire \deser_A.shift_reg[10] ;
 wire \deser_A.shift_reg[110] ;
 wire \deser_A.shift_reg[111] ;
 wire \deser_A.shift_reg[112] ;
 wire \deser_A.shift_reg[113] ;
 wire \deser_A.shift_reg[114] ;
 wire \deser_A.shift_reg[115] ;
 wire \deser_A.shift_reg[116] ;
 wire \deser_A.shift_reg[117] ;
 wire \deser_A.shift_reg[118] ;
 wire \deser_A.shift_reg[119] ;
 wire \deser_A.shift_reg[11] ;
 wire \deser_A.shift_reg[120] ;
 wire \deser_A.shift_reg[121] ;
 wire \deser_A.shift_reg[122] ;
 wire \deser_A.shift_reg[123] ;
 wire \deser_A.shift_reg[124] ;
 wire \deser_A.shift_reg[125] ;
 wire \deser_A.shift_reg[126] ;
 wire \deser_A.shift_reg[127] ;
 wire \deser_A.shift_reg[12] ;
 wire \deser_A.shift_reg[13] ;
 wire \deser_A.shift_reg[14] ;
 wire \deser_A.shift_reg[15] ;
 wire \deser_A.shift_reg[16] ;
 wire \deser_A.shift_reg[17] ;
 wire \deser_A.shift_reg[18] ;
 wire \deser_A.shift_reg[19] ;
 wire \deser_A.shift_reg[1] ;
 wire \deser_A.shift_reg[20] ;
 wire \deser_A.shift_reg[21] ;
 wire \deser_A.shift_reg[22] ;
 wire \deser_A.shift_reg[23] ;
 wire \deser_A.shift_reg[24] ;
 wire \deser_A.shift_reg[25] ;
 wire \deser_A.shift_reg[26] ;
 wire \deser_A.shift_reg[27] ;
 wire \deser_A.shift_reg[28] ;
 wire \deser_A.shift_reg[29] ;
 wire \deser_A.shift_reg[2] ;
 wire \deser_A.shift_reg[30] ;
 wire \deser_A.shift_reg[31] ;
 wire \deser_A.shift_reg[32] ;
 wire \deser_A.shift_reg[33] ;
 wire \deser_A.shift_reg[34] ;
 wire \deser_A.shift_reg[35] ;
 wire \deser_A.shift_reg[36] ;
 wire \deser_A.shift_reg[37] ;
 wire \deser_A.shift_reg[38] ;
 wire \deser_A.shift_reg[39] ;
 wire \deser_A.shift_reg[3] ;
 wire \deser_A.shift_reg[40] ;
 wire \deser_A.shift_reg[41] ;
 wire \deser_A.shift_reg[42] ;
 wire \deser_A.shift_reg[43] ;
 wire \deser_A.shift_reg[44] ;
 wire \deser_A.shift_reg[45] ;
 wire \deser_A.shift_reg[46] ;
 wire \deser_A.shift_reg[47] ;
 wire \deser_A.shift_reg[48] ;
 wire \deser_A.shift_reg[49] ;
 wire \deser_A.shift_reg[4] ;
 wire \deser_A.shift_reg[50] ;
 wire \deser_A.shift_reg[51] ;
 wire \deser_A.shift_reg[52] ;
 wire \deser_A.shift_reg[53] ;
 wire \deser_A.shift_reg[54] ;
 wire \deser_A.shift_reg[55] ;
 wire \deser_A.shift_reg[56] ;
 wire \deser_A.shift_reg[57] ;
 wire \deser_A.shift_reg[58] ;
 wire \deser_A.shift_reg[59] ;
 wire \deser_A.shift_reg[5] ;
 wire \deser_A.shift_reg[60] ;
 wire \deser_A.shift_reg[61] ;
 wire \deser_A.shift_reg[62] ;
 wire \deser_A.shift_reg[63] ;
 wire \deser_A.shift_reg[64] ;
 wire \deser_A.shift_reg[65] ;
 wire \deser_A.shift_reg[66] ;
 wire \deser_A.shift_reg[67] ;
 wire \deser_A.shift_reg[68] ;
 wire \deser_A.shift_reg[69] ;
 wire \deser_A.shift_reg[6] ;
 wire \deser_A.shift_reg[70] ;
 wire \deser_A.shift_reg[71] ;
 wire \deser_A.shift_reg[72] ;
 wire \deser_A.shift_reg[73] ;
 wire \deser_A.shift_reg[74] ;
 wire \deser_A.shift_reg[75] ;
 wire \deser_A.shift_reg[76] ;
 wire \deser_A.shift_reg[77] ;
 wire \deser_A.shift_reg[78] ;
 wire \deser_A.shift_reg[79] ;
 wire \deser_A.shift_reg[7] ;
 wire \deser_A.shift_reg[80] ;
 wire \deser_A.shift_reg[81] ;
 wire \deser_A.shift_reg[82] ;
 wire \deser_A.shift_reg[83] ;
 wire \deser_A.shift_reg[84] ;
 wire \deser_A.shift_reg[85] ;
 wire \deser_A.shift_reg[86] ;
 wire \deser_A.shift_reg[87] ;
 wire \deser_A.shift_reg[88] ;
 wire \deser_A.shift_reg[89] ;
 wire \deser_A.shift_reg[8] ;
 wire \deser_A.shift_reg[90] ;
 wire \deser_A.shift_reg[91] ;
 wire \deser_A.shift_reg[92] ;
 wire \deser_A.shift_reg[93] ;
 wire \deser_A.shift_reg[94] ;
 wire \deser_A.shift_reg[95] ;
 wire \deser_A.shift_reg[96] ;
 wire \deser_A.shift_reg[97] ;
 wire \deser_A.shift_reg[98] ;
 wire \deser_A.shift_reg[99] ;
 wire \deser_A.shift_reg[9] ;
 wire \deser_A.word_buffer[0] ;
 wire \deser_A.word_buffer[100] ;
 wire \deser_A.word_buffer[101] ;
 wire \deser_A.word_buffer[102] ;
 wire \deser_A.word_buffer[103] ;
 wire \deser_A.word_buffer[104] ;
 wire \deser_A.word_buffer[105] ;
 wire \deser_A.word_buffer[106] ;
 wire \deser_A.word_buffer[107] ;
 wire \deser_A.word_buffer[108] ;
 wire \deser_A.word_buffer[109] ;
 wire \deser_A.word_buffer[10] ;
 wire \deser_A.word_buffer[110] ;
 wire \deser_A.word_buffer[111] ;
 wire \deser_A.word_buffer[112] ;
 wire \deser_A.word_buffer[113] ;
 wire \deser_A.word_buffer[114] ;
 wire \deser_A.word_buffer[115] ;
 wire \deser_A.word_buffer[116] ;
 wire \deser_A.word_buffer[117] ;
 wire \deser_A.word_buffer[118] ;
 wire \deser_A.word_buffer[119] ;
 wire \deser_A.word_buffer[11] ;
 wire \deser_A.word_buffer[120] ;
 wire \deser_A.word_buffer[121] ;
 wire \deser_A.word_buffer[122] ;
 wire \deser_A.word_buffer[123] ;
 wire \deser_A.word_buffer[124] ;
 wire \deser_A.word_buffer[125] ;
 wire \deser_A.word_buffer[126] ;
 wire \deser_A.word_buffer[127] ;
 wire \deser_A.word_buffer[12] ;
 wire \deser_A.word_buffer[13] ;
 wire \deser_A.word_buffer[14] ;
 wire \deser_A.word_buffer[15] ;
 wire \deser_A.word_buffer[16] ;
 wire \deser_A.word_buffer[17] ;
 wire \deser_A.word_buffer[18] ;
 wire \deser_A.word_buffer[19] ;
 wire \deser_A.word_buffer[1] ;
 wire \deser_A.word_buffer[20] ;
 wire \deser_A.word_buffer[21] ;
 wire \deser_A.word_buffer[22] ;
 wire \deser_A.word_buffer[23] ;
 wire \deser_A.word_buffer[24] ;
 wire \deser_A.word_buffer[25] ;
 wire \deser_A.word_buffer[26] ;
 wire \deser_A.word_buffer[27] ;
 wire \deser_A.word_buffer[28] ;
 wire \deser_A.word_buffer[29] ;
 wire \deser_A.word_buffer[2] ;
 wire \deser_A.word_buffer[30] ;
 wire \deser_A.word_buffer[31] ;
 wire \deser_A.word_buffer[32] ;
 wire \deser_A.word_buffer[33] ;
 wire \deser_A.word_buffer[34] ;
 wire \deser_A.word_buffer[35] ;
 wire \deser_A.word_buffer[36] ;
 wire \deser_A.word_buffer[37] ;
 wire \deser_A.word_buffer[38] ;
 wire \deser_A.word_buffer[39] ;
 wire \deser_A.word_buffer[3] ;
 wire \deser_A.word_buffer[40] ;
 wire \deser_A.word_buffer[41] ;
 wire \deser_A.word_buffer[42] ;
 wire \deser_A.word_buffer[43] ;
 wire \deser_A.word_buffer[44] ;
 wire \deser_A.word_buffer[45] ;
 wire \deser_A.word_buffer[46] ;
 wire \deser_A.word_buffer[47] ;
 wire \deser_A.word_buffer[48] ;
 wire \deser_A.word_buffer[49] ;
 wire \deser_A.word_buffer[4] ;
 wire \deser_A.word_buffer[50] ;
 wire \deser_A.word_buffer[51] ;
 wire \deser_A.word_buffer[52] ;
 wire \deser_A.word_buffer[53] ;
 wire \deser_A.word_buffer[54] ;
 wire \deser_A.word_buffer[55] ;
 wire \deser_A.word_buffer[56] ;
 wire \deser_A.word_buffer[57] ;
 wire \deser_A.word_buffer[58] ;
 wire \deser_A.word_buffer[59] ;
 wire \deser_A.word_buffer[5] ;
 wire \deser_A.word_buffer[60] ;
 wire \deser_A.word_buffer[61] ;
 wire \deser_A.word_buffer[62] ;
 wire \deser_A.word_buffer[63] ;
 wire \deser_A.word_buffer[64] ;
 wire \deser_A.word_buffer[65] ;
 wire \deser_A.word_buffer[66] ;
 wire \deser_A.word_buffer[67] ;
 wire \deser_A.word_buffer[68] ;
 wire \deser_A.word_buffer[69] ;
 wire \deser_A.word_buffer[6] ;
 wire \deser_A.word_buffer[70] ;
 wire \deser_A.word_buffer[71] ;
 wire \deser_A.word_buffer[72] ;
 wire \deser_A.word_buffer[73] ;
 wire \deser_A.word_buffer[74] ;
 wire \deser_A.word_buffer[75] ;
 wire \deser_A.word_buffer[76] ;
 wire \deser_A.word_buffer[77] ;
 wire \deser_A.word_buffer[78] ;
 wire \deser_A.word_buffer[79] ;
 wire \deser_A.word_buffer[7] ;
 wire \deser_A.word_buffer[80] ;
 wire \deser_A.word_buffer[81] ;
 wire \deser_A.word_buffer[82] ;
 wire \deser_A.word_buffer[83] ;
 wire \deser_A.word_buffer[84] ;
 wire \deser_A.word_buffer[85] ;
 wire \deser_A.word_buffer[86] ;
 wire \deser_A.word_buffer[87] ;
 wire \deser_A.word_buffer[88] ;
 wire \deser_A.word_buffer[89] ;
 wire \deser_A.word_buffer[8] ;
 wire \deser_A.word_buffer[90] ;
 wire \deser_A.word_buffer[91] ;
 wire \deser_A.word_buffer[92] ;
 wire \deser_A.word_buffer[93] ;
 wire \deser_A.word_buffer[94] ;
 wire \deser_A.word_buffer[95] ;
 wire \deser_A.word_buffer[96] ;
 wire \deser_A.word_buffer[97] ;
 wire \deser_A.word_buffer[98] ;
 wire \deser_A.word_buffer[99] ;
 wire \deser_A.word_buffer[9] ;
 wire \deser_B.bit_idx[0] ;
 wire \deser_B.bit_idx[1] ;
 wire \deser_B.bit_idx[2] ;
 wire \deser_B.bit_idx[3] ;
 wire \deser_B.bit_idx[4] ;
 wire \deser_B.bit_idx[5] ;
 wire \deser_B.bit_idx[6] ;
 wire \deser_B.receiving ;
 wire \deser_B.serial_toggle ;
 wire \deser_B.serial_toggle_sync1 ;
 wire \deser_B.serial_toggle_sync2 ;
 wire \deser_B.serial_word[0] ;
 wire \deser_B.serial_word[100] ;
 wire \deser_B.serial_word[101] ;
 wire \deser_B.serial_word[102] ;
 wire \deser_B.serial_word[103] ;
 wire \deser_B.serial_word[104] ;
 wire \deser_B.serial_word[105] ;
 wire \deser_B.serial_word[106] ;
 wire \deser_B.serial_word[107] ;
 wire \deser_B.serial_word[108] ;
 wire \deser_B.serial_word[109] ;
 wire \deser_B.serial_word[10] ;
 wire \deser_B.serial_word[110] ;
 wire \deser_B.serial_word[111] ;
 wire \deser_B.serial_word[112] ;
 wire \deser_B.serial_word[113] ;
 wire \deser_B.serial_word[114] ;
 wire \deser_B.serial_word[115] ;
 wire \deser_B.serial_word[116] ;
 wire \deser_B.serial_word[117] ;
 wire \deser_B.serial_word[118] ;
 wire \deser_B.serial_word[119] ;
 wire \deser_B.serial_word[11] ;
 wire \deser_B.serial_word[120] ;
 wire \deser_B.serial_word[121] ;
 wire \deser_B.serial_word[122] ;
 wire \deser_B.serial_word[123] ;
 wire \deser_B.serial_word[124] ;
 wire \deser_B.serial_word[125] ;
 wire \deser_B.serial_word[126] ;
 wire \deser_B.serial_word[127] ;
 wire \deser_B.serial_word[12] ;
 wire \deser_B.serial_word[13] ;
 wire \deser_B.serial_word[14] ;
 wire \deser_B.serial_word[15] ;
 wire \deser_B.serial_word[16] ;
 wire \deser_B.serial_word[17] ;
 wire \deser_B.serial_word[18] ;
 wire \deser_B.serial_word[19] ;
 wire \deser_B.serial_word[1] ;
 wire \deser_B.serial_word[20] ;
 wire \deser_B.serial_word[21] ;
 wire \deser_B.serial_word[22] ;
 wire \deser_B.serial_word[23] ;
 wire \deser_B.serial_word[24] ;
 wire \deser_B.serial_word[25] ;
 wire \deser_B.serial_word[26] ;
 wire \deser_B.serial_word[27] ;
 wire \deser_B.serial_word[28] ;
 wire \deser_B.serial_word[29] ;
 wire \deser_B.serial_word[2] ;
 wire \deser_B.serial_word[30] ;
 wire \deser_B.serial_word[31] ;
 wire \deser_B.serial_word[32] ;
 wire \deser_B.serial_word[33] ;
 wire \deser_B.serial_word[34] ;
 wire \deser_B.serial_word[35] ;
 wire \deser_B.serial_word[36] ;
 wire \deser_B.serial_word[37] ;
 wire \deser_B.serial_word[38] ;
 wire \deser_B.serial_word[39] ;
 wire \deser_B.serial_word[3] ;
 wire \deser_B.serial_word[40] ;
 wire \deser_B.serial_word[41] ;
 wire \deser_B.serial_word[42] ;
 wire \deser_B.serial_word[43] ;
 wire \deser_B.serial_word[44] ;
 wire \deser_B.serial_word[45] ;
 wire \deser_B.serial_word[46] ;
 wire \deser_B.serial_word[47] ;
 wire \deser_B.serial_word[48] ;
 wire \deser_B.serial_word[49] ;
 wire \deser_B.serial_word[4] ;
 wire \deser_B.serial_word[50] ;
 wire \deser_B.serial_word[51] ;
 wire \deser_B.serial_word[52] ;
 wire \deser_B.serial_word[53] ;
 wire \deser_B.serial_word[54] ;
 wire \deser_B.serial_word[55] ;
 wire \deser_B.serial_word[56] ;
 wire \deser_B.serial_word[57] ;
 wire \deser_B.serial_word[58] ;
 wire \deser_B.serial_word[59] ;
 wire \deser_B.serial_word[5] ;
 wire \deser_B.serial_word[60] ;
 wire \deser_B.serial_word[61] ;
 wire \deser_B.serial_word[62] ;
 wire \deser_B.serial_word[63] ;
 wire \deser_B.serial_word[64] ;
 wire \deser_B.serial_word[65] ;
 wire \deser_B.serial_word[66] ;
 wire \deser_B.serial_word[67] ;
 wire \deser_B.serial_word[68] ;
 wire \deser_B.serial_word[69] ;
 wire \deser_B.serial_word[6] ;
 wire \deser_B.serial_word[70] ;
 wire \deser_B.serial_word[71] ;
 wire \deser_B.serial_word[72] ;
 wire \deser_B.serial_word[73] ;
 wire \deser_B.serial_word[74] ;
 wire \deser_B.serial_word[75] ;
 wire \deser_B.serial_word[76] ;
 wire \deser_B.serial_word[77] ;
 wire \deser_B.serial_word[78] ;
 wire \deser_B.serial_word[79] ;
 wire \deser_B.serial_word[7] ;
 wire \deser_B.serial_word[80] ;
 wire \deser_B.serial_word[81] ;
 wire \deser_B.serial_word[82] ;
 wire \deser_B.serial_word[83] ;
 wire \deser_B.serial_word[84] ;
 wire \deser_B.serial_word[85] ;
 wire \deser_B.serial_word[86] ;
 wire \deser_B.serial_word[87] ;
 wire \deser_B.serial_word[88] ;
 wire \deser_B.serial_word[89] ;
 wire \deser_B.serial_word[8] ;
 wire \deser_B.serial_word[90] ;
 wire \deser_B.serial_word[91] ;
 wire \deser_B.serial_word[92] ;
 wire \deser_B.serial_word[93] ;
 wire \deser_B.serial_word[94] ;
 wire \deser_B.serial_word[95] ;
 wire \deser_B.serial_word[96] ;
 wire \deser_B.serial_word[97] ;
 wire \deser_B.serial_word[98] ;
 wire \deser_B.serial_word[99] ;
 wire \deser_B.serial_word[9] ;
 wire \deser_B.serial_word_ready ;
 wire \deser_B.shift_reg[0] ;
 wire \deser_B.shift_reg[100] ;
 wire \deser_B.shift_reg[101] ;
 wire \deser_B.shift_reg[102] ;
 wire \deser_B.shift_reg[103] ;
 wire \deser_B.shift_reg[104] ;
 wire \deser_B.shift_reg[105] ;
 wire \deser_B.shift_reg[106] ;
 wire \deser_B.shift_reg[107] ;
 wire \deser_B.shift_reg[108] ;
 wire \deser_B.shift_reg[109] ;
 wire \deser_B.shift_reg[10] ;
 wire \deser_B.shift_reg[110] ;
 wire \deser_B.shift_reg[111] ;
 wire \deser_B.shift_reg[112] ;
 wire \deser_B.shift_reg[113] ;
 wire \deser_B.shift_reg[114] ;
 wire \deser_B.shift_reg[115] ;
 wire \deser_B.shift_reg[116] ;
 wire \deser_B.shift_reg[117] ;
 wire \deser_B.shift_reg[118] ;
 wire \deser_B.shift_reg[119] ;
 wire \deser_B.shift_reg[11] ;
 wire \deser_B.shift_reg[120] ;
 wire \deser_B.shift_reg[121] ;
 wire \deser_B.shift_reg[122] ;
 wire \deser_B.shift_reg[123] ;
 wire \deser_B.shift_reg[124] ;
 wire \deser_B.shift_reg[125] ;
 wire \deser_B.shift_reg[126] ;
 wire \deser_B.shift_reg[127] ;
 wire \deser_B.shift_reg[12] ;
 wire \deser_B.shift_reg[13] ;
 wire \deser_B.shift_reg[14] ;
 wire \deser_B.shift_reg[15] ;
 wire \deser_B.shift_reg[16] ;
 wire \deser_B.shift_reg[17] ;
 wire \deser_B.shift_reg[18] ;
 wire \deser_B.shift_reg[19] ;
 wire \deser_B.shift_reg[1] ;
 wire \deser_B.shift_reg[20] ;
 wire \deser_B.shift_reg[21] ;
 wire \deser_B.shift_reg[22] ;
 wire \deser_B.shift_reg[23] ;
 wire \deser_B.shift_reg[24] ;
 wire \deser_B.shift_reg[25] ;
 wire \deser_B.shift_reg[26] ;
 wire \deser_B.shift_reg[27] ;
 wire \deser_B.shift_reg[28] ;
 wire \deser_B.shift_reg[29] ;
 wire \deser_B.shift_reg[2] ;
 wire \deser_B.shift_reg[30] ;
 wire \deser_B.shift_reg[31] ;
 wire \deser_B.shift_reg[32] ;
 wire \deser_B.shift_reg[33] ;
 wire \deser_B.shift_reg[34] ;
 wire \deser_B.shift_reg[35] ;
 wire \deser_B.shift_reg[36] ;
 wire \deser_B.shift_reg[37] ;
 wire \deser_B.shift_reg[38] ;
 wire \deser_B.shift_reg[39] ;
 wire \deser_B.shift_reg[3] ;
 wire \deser_B.shift_reg[40] ;
 wire \deser_B.shift_reg[41] ;
 wire \deser_B.shift_reg[42] ;
 wire \deser_B.shift_reg[43] ;
 wire \deser_B.shift_reg[44] ;
 wire \deser_B.shift_reg[45] ;
 wire \deser_B.shift_reg[46] ;
 wire \deser_B.shift_reg[47] ;
 wire \deser_B.shift_reg[48] ;
 wire \deser_B.shift_reg[49] ;
 wire \deser_B.shift_reg[4] ;
 wire \deser_B.shift_reg[50] ;
 wire \deser_B.shift_reg[51] ;
 wire \deser_B.shift_reg[52] ;
 wire \deser_B.shift_reg[53] ;
 wire \deser_B.shift_reg[54] ;
 wire \deser_B.shift_reg[55] ;
 wire \deser_B.shift_reg[56] ;
 wire \deser_B.shift_reg[57] ;
 wire \deser_B.shift_reg[58] ;
 wire \deser_B.shift_reg[59] ;
 wire \deser_B.shift_reg[5] ;
 wire \deser_B.shift_reg[60] ;
 wire \deser_B.shift_reg[61] ;
 wire \deser_B.shift_reg[62] ;
 wire \deser_B.shift_reg[63] ;
 wire \deser_B.shift_reg[64] ;
 wire \deser_B.shift_reg[65] ;
 wire \deser_B.shift_reg[66] ;
 wire \deser_B.shift_reg[67] ;
 wire \deser_B.shift_reg[68] ;
 wire \deser_B.shift_reg[69] ;
 wire \deser_B.shift_reg[6] ;
 wire \deser_B.shift_reg[70] ;
 wire \deser_B.shift_reg[71] ;
 wire \deser_B.shift_reg[72] ;
 wire \deser_B.shift_reg[73] ;
 wire \deser_B.shift_reg[74] ;
 wire \deser_B.shift_reg[75] ;
 wire \deser_B.shift_reg[76] ;
 wire \deser_B.shift_reg[77] ;
 wire \deser_B.shift_reg[78] ;
 wire \deser_B.shift_reg[79] ;
 wire \deser_B.shift_reg[7] ;
 wire \deser_B.shift_reg[80] ;
 wire \deser_B.shift_reg[81] ;
 wire \deser_B.shift_reg[82] ;
 wire \deser_B.shift_reg[83] ;
 wire \deser_B.shift_reg[84] ;
 wire \deser_B.shift_reg[85] ;
 wire \deser_B.shift_reg[86] ;
 wire \deser_B.shift_reg[87] ;
 wire \deser_B.shift_reg[88] ;
 wire \deser_B.shift_reg[89] ;
 wire \deser_B.shift_reg[8] ;
 wire \deser_B.shift_reg[90] ;
 wire \deser_B.shift_reg[91] ;
 wire \deser_B.shift_reg[92] ;
 wire \deser_B.shift_reg[93] ;
 wire \deser_B.shift_reg[94] ;
 wire \deser_B.shift_reg[95] ;
 wire \deser_B.shift_reg[96] ;
 wire \deser_B.shift_reg[97] ;
 wire \deser_B.shift_reg[98] ;
 wire \deser_B.shift_reg[99] ;
 wire \deser_B.shift_reg[9] ;
 wire \deser_B.word_buffer[0] ;
 wire \deser_B.word_buffer[100] ;
 wire \deser_B.word_buffer[101] ;
 wire \deser_B.word_buffer[102] ;
 wire \deser_B.word_buffer[103] ;
 wire \deser_B.word_buffer[104] ;
 wire \deser_B.word_buffer[105] ;
 wire \deser_B.word_buffer[106] ;
 wire \deser_B.word_buffer[107] ;
 wire \deser_B.word_buffer[108] ;
 wire \deser_B.word_buffer[109] ;
 wire \deser_B.word_buffer[10] ;
 wire \deser_B.word_buffer[110] ;
 wire \deser_B.word_buffer[111] ;
 wire \deser_B.word_buffer[112] ;
 wire \deser_B.word_buffer[113] ;
 wire \deser_B.word_buffer[114] ;
 wire \deser_B.word_buffer[115] ;
 wire \deser_B.word_buffer[116] ;
 wire \deser_B.word_buffer[117] ;
 wire \deser_B.word_buffer[118] ;
 wire \deser_B.word_buffer[119] ;
 wire \deser_B.word_buffer[11] ;
 wire \deser_B.word_buffer[120] ;
 wire \deser_B.word_buffer[121] ;
 wire \deser_B.word_buffer[122] ;
 wire \deser_B.word_buffer[123] ;
 wire \deser_B.word_buffer[124] ;
 wire \deser_B.word_buffer[125] ;
 wire \deser_B.word_buffer[126] ;
 wire \deser_B.word_buffer[127] ;
 wire \deser_B.word_buffer[12] ;
 wire \deser_B.word_buffer[13] ;
 wire \deser_B.word_buffer[14] ;
 wire \deser_B.word_buffer[15] ;
 wire \deser_B.word_buffer[16] ;
 wire \deser_B.word_buffer[17] ;
 wire \deser_B.word_buffer[18] ;
 wire \deser_B.word_buffer[19] ;
 wire \deser_B.word_buffer[1] ;
 wire \deser_B.word_buffer[20] ;
 wire \deser_B.word_buffer[21] ;
 wire \deser_B.word_buffer[22] ;
 wire \deser_B.word_buffer[23] ;
 wire \deser_B.word_buffer[24] ;
 wire \deser_B.word_buffer[25] ;
 wire \deser_B.word_buffer[26] ;
 wire \deser_B.word_buffer[27] ;
 wire \deser_B.word_buffer[28] ;
 wire \deser_B.word_buffer[29] ;
 wire \deser_B.word_buffer[2] ;
 wire \deser_B.word_buffer[30] ;
 wire \deser_B.word_buffer[31] ;
 wire \deser_B.word_buffer[32] ;
 wire \deser_B.word_buffer[33] ;
 wire \deser_B.word_buffer[34] ;
 wire \deser_B.word_buffer[35] ;
 wire \deser_B.word_buffer[36] ;
 wire \deser_B.word_buffer[37] ;
 wire \deser_B.word_buffer[38] ;
 wire \deser_B.word_buffer[39] ;
 wire \deser_B.word_buffer[3] ;
 wire \deser_B.word_buffer[40] ;
 wire \deser_B.word_buffer[41] ;
 wire \deser_B.word_buffer[42] ;
 wire \deser_B.word_buffer[43] ;
 wire \deser_B.word_buffer[44] ;
 wire \deser_B.word_buffer[45] ;
 wire \deser_B.word_buffer[46] ;
 wire \deser_B.word_buffer[47] ;
 wire \deser_B.word_buffer[48] ;
 wire \deser_B.word_buffer[49] ;
 wire \deser_B.word_buffer[4] ;
 wire \deser_B.word_buffer[50] ;
 wire \deser_B.word_buffer[51] ;
 wire \deser_B.word_buffer[52] ;
 wire \deser_B.word_buffer[53] ;
 wire \deser_B.word_buffer[54] ;
 wire \deser_B.word_buffer[55] ;
 wire \deser_B.word_buffer[56] ;
 wire \deser_B.word_buffer[57] ;
 wire \deser_B.word_buffer[58] ;
 wire \deser_B.word_buffer[59] ;
 wire \deser_B.word_buffer[5] ;
 wire \deser_B.word_buffer[60] ;
 wire \deser_B.word_buffer[61] ;
 wire \deser_B.word_buffer[62] ;
 wire \deser_B.word_buffer[63] ;
 wire \deser_B.word_buffer[64] ;
 wire \deser_B.word_buffer[65] ;
 wire \deser_B.word_buffer[66] ;
 wire \deser_B.word_buffer[67] ;
 wire \deser_B.word_buffer[68] ;
 wire \deser_B.word_buffer[69] ;
 wire \deser_B.word_buffer[6] ;
 wire \deser_B.word_buffer[70] ;
 wire \deser_B.word_buffer[71] ;
 wire \deser_B.word_buffer[72] ;
 wire \deser_B.word_buffer[73] ;
 wire \deser_B.word_buffer[74] ;
 wire \deser_B.word_buffer[75] ;
 wire \deser_B.word_buffer[76] ;
 wire \deser_B.word_buffer[77] ;
 wire \deser_B.word_buffer[78] ;
 wire \deser_B.word_buffer[79] ;
 wire \deser_B.word_buffer[7] ;
 wire \deser_B.word_buffer[80] ;
 wire \deser_B.word_buffer[81] ;
 wire \deser_B.word_buffer[82] ;
 wire \deser_B.word_buffer[83] ;
 wire \deser_B.word_buffer[84] ;
 wire \deser_B.word_buffer[85] ;
 wire \deser_B.word_buffer[86] ;
 wire \deser_B.word_buffer[87] ;
 wire \deser_B.word_buffer[88] ;
 wire \deser_B.word_buffer[89] ;
 wire \deser_B.word_buffer[8] ;
 wire \deser_B.word_buffer[90] ;
 wire \deser_B.word_buffer[91] ;
 wire \deser_B.word_buffer[92] ;
 wire \deser_B.word_buffer[93] ;
 wire \deser_B.word_buffer[94] ;
 wire \deser_B.word_buffer[95] ;
 wire \deser_B.word_buffer[96] ;
 wire \deser_B.word_buffer[97] ;
 wire \deser_B.word_buffer[98] ;
 wire \deser_B.word_buffer[99] ;
 wire \deser_B.word_buffer[9] ;
 wire \ser_C.bit_idx[0] ;
 wire \ser_C.bit_idx[1] ;
 wire \ser_C.bit_idx[2] ;
 wire \ser_C.bit_idx[3] ;
 wire \ser_C.bit_idx[4] ;
 wire \ser_C.bit_idx[5] ;
 wire \ser_C.bit_idx[6] ;
 wire \ser_C.bit_idx[7] ;
 wire \ser_C.bit_idx[8] ;
 wire \ser_C.parallel_data[440] ;
 wire \ser_C.parallel_data[441] ;
 wire \ser_C.parallel_data[442] ;
 wire \ser_C.parallel_data[443] ;
 wire \ser_C.parallel_data[444] ;
 wire \ser_C.parallel_data[445] ;
 wire \ser_C.parallel_data[446] ;
 wire \ser_C.parallel_data[447] ;
 wire \ser_C.parallel_data[448] ;
 wire \ser_C.parallel_data[449] ;
 wire \ser_C.parallel_data[450] ;
 wire \ser_C.parallel_data[451] ;
 wire \ser_C.parallel_data[452] ;
 wire \ser_C.parallel_data[453] ;
 wire \ser_C.parallel_data[454] ;
 wire \ser_C.parallel_data[455] ;
 wire \ser_C.parallel_data[456] ;
 wire \ser_C.parallel_data[457] ;
 wire \ser_C.parallel_data[458] ;
 wire \ser_C.parallel_data[459] ;
 wire \ser_C.parallel_data[460] ;
 wire \ser_C.parallel_data[461] ;
 wire \ser_C.parallel_data[462] ;
 wire \ser_C.parallel_data[463] ;
 wire \ser_C.parallel_data[464] ;
 wire \ser_C.parallel_data[465] ;
 wire \ser_C.parallel_data[466] ;
 wire \ser_C.parallel_data[467] ;
 wire \ser_C.parallel_data[468] ;
 wire \ser_C.parallel_data[469] ;
 wire \ser_C.parallel_data[470] ;
 wire \ser_C.parallel_data[471] ;
 wire \ser_C.parallel_data[472] ;
 wire \ser_C.parallel_data[473] ;
 wire \ser_C.parallel_data[474] ;
 wire \ser_C.parallel_data[475] ;
 wire \ser_C.parallel_data[476] ;
 wire \ser_C.parallel_data[477] ;
 wire \ser_C.parallel_data[478] ;
 wire \ser_C.parallel_data[479] ;
 wire \ser_C.parallel_data[480] ;
 wire \ser_C.parallel_data[481] ;
 wire \ser_C.parallel_data[482] ;
 wire \ser_C.parallel_data[483] ;
 wire \ser_C.parallel_data[484] ;
 wire \ser_C.parallel_data[485] ;
 wire \ser_C.parallel_data[486] ;
 wire \ser_C.parallel_data[487] ;
 wire \ser_C.parallel_data[488] ;
 wire \ser_C.parallel_data[489] ;
 wire \ser_C.parallel_data[490] ;
 wire \ser_C.parallel_data[491] ;
 wire \ser_C.parallel_data[492] ;
 wire \ser_C.parallel_data[493] ;
 wire \ser_C.parallel_data[494] ;
 wire \ser_C.parallel_data[495] ;
 wire \ser_C.parallel_data[496] ;
 wire \ser_C.parallel_data[497] ;
 wire \ser_C.parallel_data[498] ;
 wire \ser_C.parallel_data[499] ;
 wire \ser_C.parallel_data[500] ;
 wire \ser_C.parallel_data[501] ;
 wire \ser_C.parallel_data[502] ;
 wire \ser_C.parallel_data[503] ;
 wire \ser_C.parallel_data[504] ;
 wire \ser_C.parallel_data[505] ;
 wire \ser_C.parallel_data[506] ;
 wire \ser_C.parallel_data[507] ;
 wire \ser_C.parallel_data[508] ;
 wire \ser_C.parallel_data[509] ;
 wire \ser_C.parallel_data[510] ;
 wire \ser_C.parallel_data[511] ;
 wire \ser_C.shift_reg[0] ;
 wire \ser_C.shift_reg[100] ;
 wire \ser_C.shift_reg[101] ;
 wire \ser_C.shift_reg[102] ;
 wire \ser_C.shift_reg[103] ;
 wire \ser_C.shift_reg[104] ;
 wire \ser_C.shift_reg[105] ;
 wire \ser_C.shift_reg[106] ;
 wire \ser_C.shift_reg[107] ;
 wire \ser_C.shift_reg[108] ;
 wire \ser_C.shift_reg[109] ;
 wire \ser_C.shift_reg[10] ;
 wire \ser_C.shift_reg[110] ;
 wire \ser_C.shift_reg[111] ;
 wire \ser_C.shift_reg[112] ;
 wire \ser_C.shift_reg[113] ;
 wire \ser_C.shift_reg[114] ;
 wire \ser_C.shift_reg[115] ;
 wire \ser_C.shift_reg[116] ;
 wire \ser_C.shift_reg[117] ;
 wire \ser_C.shift_reg[118] ;
 wire \ser_C.shift_reg[119] ;
 wire \ser_C.shift_reg[11] ;
 wire \ser_C.shift_reg[120] ;
 wire \ser_C.shift_reg[121] ;
 wire \ser_C.shift_reg[122] ;
 wire \ser_C.shift_reg[123] ;
 wire \ser_C.shift_reg[124] ;
 wire \ser_C.shift_reg[125] ;
 wire \ser_C.shift_reg[126] ;
 wire \ser_C.shift_reg[127] ;
 wire \ser_C.shift_reg[128] ;
 wire \ser_C.shift_reg[129] ;
 wire \ser_C.shift_reg[12] ;
 wire \ser_C.shift_reg[130] ;
 wire \ser_C.shift_reg[131] ;
 wire \ser_C.shift_reg[132] ;
 wire \ser_C.shift_reg[133] ;
 wire \ser_C.shift_reg[134] ;
 wire \ser_C.shift_reg[135] ;
 wire \ser_C.shift_reg[136] ;
 wire \ser_C.shift_reg[137] ;
 wire \ser_C.shift_reg[138] ;
 wire \ser_C.shift_reg[139] ;
 wire \ser_C.shift_reg[13] ;
 wire \ser_C.shift_reg[140] ;
 wire \ser_C.shift_reg[141] ;
 wire \ser_C.shift_reg[142] ;
 wire \ser_C.shift_reg[143] ;
 wire \ser_C.shift_reg[144] ;
 wire \ser_C.shift_reg[145] ;
 wire \ser_C.shift_reg[146] ;
 wire \ser_C.shift_reg[147] ;
 wire \ser_C.shift_reg[148] ;
 wire \ser_C.shift_reg[149] ;
 wire \ser_C.shift_reg[14] ;
 wire \ser_C.shift_reg[150] ;
 wire \ser_C.shift_reg[151] ;
 wire \ser_C.shift_reg[152] ;
 wire \ser_C.shift_reg[153] ;
 wire \ser_C.shift_reg[154] ;
 wire \ser_C.shift_reg[155] ;
 wire \ser_C.shift_reg[156] ;
 wire \ser_C.shift_reg[157] ;
 wire \ser_C.shift_reg[158] ;
 wire \ser_C.shift_reg[159] ;
 wire \ser_C.shift_reg[15] ;
 wire \ser_C.shift_reg[160] ;
 wire \ser_C.shift_reg[161] ;
 wire \ser_C.shift_reg[162] ;
 wire \ser_C.shift_reg[163] ;
 wire \ser_C.shift_reg[164] ;
 wire \ser_C.shift_reg[165] ;
 wire \ser_C.shift_reg[166] ;
 wire \ser_C.shift_reg[167] ;
 wire \ser_C.shift_reg[168] ;
 wire \ser_C.shift_reg[169] ;
 wire \ser_C.shift_reg[16] ;
 wire \ser_C.shift_reg[170] ;
 wire \ser_C.shift_reg[171] ;
 wire \ser_C.shift_reg[172] ;
 wire \ser_C.shift_reg[173] ;
 wire \ser_C.shift_reg[174] ;
 wire \ser_C.shift_reg[175] ;
 wire \ser_C.shift_reg[176] ;
 wire \ser_C.shift_reg[177] ;
 wire \ser_C.shift_reg[178] ;
 wire \ser_C.shift_reg[179] ;
 wire \ser_C.shift_reg[17] ;
 wire \ser_C.shift_reg[180] ;
 wire \ser_C.shift_reg[181] ;
 wire \ser_C.shift_reg[182] ;
 wire \ser_C.shift_reg[183] ;
 wire \ser_C.shift_reg[184] ;
 wire \ser_C.shift_reg[185] ;
 wire \ser_C.shift_reg[186] ;
 wire \ser_C.shift_reg[187] ;
 wire \ser_C.shift_reg[188] ;
 wire \ser_C.shift_reg[189] ;
 wire \ser_C.shift_reg[18] ;
 wire \ser_C.shift_reg[190] ;
 wire \ser_C.shift_reg[191] ;
 wire \ser_C.shift_reg[192] ;
 wire \ser_C.shift_reg[193] ;
 wire \ser_C.shift_reg[194] ;
 wire \ser_C.shift_reg[195] ;
 wire \ser_C.shift_reg[196] ;
 wire \ser_C.shift_reg[197] ;
 wire \ser_C.shift_reg[198] ;
 wire \ser_C.shift_reg[199] ;
 wire \ser_C.shift_reg[19] ;
 wire \ser_C.shift_reg[1] ;
 wire \ser_C.shift_reg[200] ;
 wire \ser_C.shift_reg[201] ;
 wire \ser_C.shift_reg[202] ;
 wire \ser_C.shift_reg[203] ;
 wire \ser_C.shift_reg[204] ;
 wire \ser_C.shift_reg[205] ;
 wire \ser_C.shift_reg[206] ;
 wire \ser_C.shift_reg[207] ;
 wire \ser_C.shift_reg[208] ;
 wire \ser_C.shift_reg[209] ;
 wire \ser_C.shift_reg[20] ;
 wire \ser_C.shift_reg[210] ;
 wire \ser_C.shift_reg[211] ;
 wire \ser_C.shift_reg[212] ;
 wire \ser_C.shift_reg[213] ;
 wire \ser_C.shift_reg[214] ;
 wire \ser_C.shift_reg[215] ;
 wire \ser_C.shift_reg[216] ;
 wire \ser_C.shift_reg[217] ;
 wire \ser_C.shift_reg[218] ;
 wire \ser_C.shift_reg[219] ;
 wire \ser_C.shift_reg[21] ;
 wire \ser_C.shift_reg[220] ;
 wire \ser_C.shift_reg[221] ;
 wire \ser_C.shift_reg[222] ;
 wire \ser_C.shift_reg[223] ;
 wire \ser_C.shift_reg[224] ;
 wire \ser_C.shift_reg[225] ;
 wire \ser_C.shift_reg[226] ;
 wire \ser_C.shift_reg[227] ;
 wire \ser_C.shift_reg[228] ;
 wire \ser_C.shift_reg[229] ;
 wire \ser_C.shift_reg[22] ;
 wire \ser_C.shift_reg[230] ;
 wire \ser_C.shift_reg[231] ;
 wire \ser_C.shift_reg[232] ;
 wire \ser_C.shift_reg[233] ;
 wire \ser_C.shift_reg[234] ;
 wire \ser_C.shift_reg[235] ;
 wire \ser_C.shift_reg[236] ;
 wire \ser_C.shift_reg[237] ;
 wire \ser_C.shift_reg[238] ;
 wire \ser_C.shift_reg[239] ;
 wire \ser_C.shift_reg[23] ;
 wire \ser_C.shift_reg[240] ;
 wire \ser_C.shift_reg[241] ;
 wire \ser_C.shift_reg[242] ;
 wire \ser_C.shift_reg[243] ;
 wire \ser_C.shift_reg[244] ;
 wire \ser_C.shift_reg[245] ;
 wire \ser_C.shift_reg[246] ;
 wire \ser_C.shift_reg[247] ;
 wire \ser_C.shift_reg[248] ;
 wire \ser_C.shift_reg[249] ;
 wire \ser_C.shift_reg[24] ;
 wire \ser_C.shift_reg[250] ;
 wire \ser_C.shift_reg[251] ;
 wire \ser_C.shift_reg[252] ;
 wire \ser_C.shift_reg[253] ;
 wire \ser_C.shift_reg[254] ;
 wire \ser_C.shift_reg[255] ;
 wire \ser_C.shift_reg[256] ;
 wire \ser_C.shift_reg[257] ;
 wire \ser_C.shift_reg[258] ;
 wire \ser_C.shift_reg[259] ;
 wire \ser_C.shift_reg[25] ;
 wire \ser_C.shift_reg[260] ;
 wire \ser_C.shift_reg[261] ;
 wire \ser_C.shift_reg[262] ;
 wire \ser_C.shift_reg[263] ;
 wire \ser_C.shift_reg[264] ;
 wire \ser_C.shift_reg[265] ;
 wire \ser_C.shift_reg[266] ;
 wire \ser_C.shift_reg[267] ;
 wire \ser_C.shift_reg[268] ;
 wire \ser_C.shift_reg[269] ;
 wire \ser_C.shift_reg[26] ;
 wire \ser_C.shift_reg[270] ;
 wire \ser_C.shift_reg[271] ;
 wire \ser_C.shift_reg[272] ;
 wire \ser_C.shift_reg[273] ;
 wire \ser_C.shift_reg[274] ;
 wire \ser_C.shift_reg[275] ;
 wire \ser_C.shift_reg[276] ;
 wire \ser_C.shift_reg[277] ;
 wire \ser_C.shift_reg[278] ;
 wire \ser_C.shift_reg[279] ;
 wire \ser_C.shift_reg[27] ;
 wire \ser_C.shift_reg[280] ;
 wire \ser_C.shift_reg[281] ;
 wire \ser_C.shift_reg[282] ;
 wire \ser_C.shift_reg[283] ;
 wire \ser_C.shift_reg[284] ;
 wire \ser_C.shift_reg[285] ;
 wire \ser_C.shift_reg[286] ;
 wire \ser_C.shift_reg[287] ;
 wire \ser_C.shift_reg[288] ;
 wire \ser_C.shift_reg[289] ;
 wire \ser_C.shift_reg[28] ;
 wire \ser_C.shift_reg[290] ;
 wire \ser_C.shift_reg[291] ;
 wire \ser_C.shift_reg[292] ;
 wire \ser_C.shift_reg[293] ;
 wire \ser_C.shift_reg[294] ;
 wire \ser_C.shift_reg[295] ;
 wire \ser_C.shift_reg[296] ;
 wire \ser_C.shift_reg[297] ;
 wire \ser_C.shift_reg[298] ;
 wire \ser_C.shift_reg[299] ;
 wire \ser_C.shift_reg[29] ;
 wire \ser_C.shift_reg[2] ;
 wire \ser_C.shift_reg[300] ;
 wire \ser_C.shift_reg[301] ;
 wire \ser_C.shift_reg[302] ;
 wire \ser_C.shift_reg[303] ;
 wire \ser_C.shift_reg[304] ;
 wire \ser_C.shift_reg[305] ;
 wire \ser_C.shift_reg[306] ;
 wire \ser_C.shift_reg[307] ;
 wire \ser_C.shift_reg[308] ;
 wire \ser_C.shift_reg[309] ;
 wire \ser_C.shift_reg[30] ;
 wire \ser_C.shift_reg[310] ;
 wire \ser_C.shift_reg[311] ;
 wire \ser_C.shift_reg[312] ;
 wire \ser_C.shift_reg[313] ;
 wire \ser_C.shift_reg[314] ;
 wire \ser_C.shift_reg[315] ;
 wire \ser_C.shift_reg[316] ;
 wire \ser_C.shift_reg[317] ;
 wire \ser_C.shift_reg[318] ;
 wire \ser_C.shift_reg[319] ;
 wire \ser_C.shift_reg[31] ;
 wire \ser_C.shift_reg[320] ;
 wire \ser_C.shift_reg[321] ;
 wire \ser_C.shift_reg[322] ;
 wire \ser_C.shift_reg[323] ;
 wire \ser_C.shift_reg[324] ;
 wire \ser_C.shift_reg[325] ;
 wire \ser_C.shift_reg[326] ;
 wire \ser_C.shift_reg[327] ;
 wire \ser_C.shift_reg[328] ;
 wire \ser_C.shift_reg[329] ;
 wire \ser_C.shift_reg[32] ;
 wire \ser_C.shift_reg[330] ;
 wire \ser_C.shift_reg[331] ;
 wire \ser_C.shift_reg[332] ;
 wire \ser_C.shift_reg[333] ;
 wire \ser_C.shift_reg[334] ;
 wire \ser_C.shift_reg[335] ;
 wire \ser_C.shift_reg[336] ;
 wire \ser_C.shift_reg[337] ;
 wire \ser_C.shift_reg[338] ;
 wire \ser_C.shift_reg[339] ;
 wire \ser_C.shift_reg[33] ;
 wire \ser_C.shift_reg[340] ;
 wire \ser_C.shift_reg[341] ;
 wire \ser_C.shift_reg[342] ;
 wire \ser_C.shift_reg[343] ;
 wire \ser_C.shift_reg[344] ;
 wire \ser_C.shift_reg[345] ;
 wire \ser_C.shift_reg[346] ;
 wire \ser_C.shift_reg[347] ;
 wire \ser_C.shift_reg[348] ;
 wire \ser_C.shift_reg[349] ;
 wire \ser_C.shift_reg[34] ;
 wire \ser_C.shift_reg[350] ;
 wire \ser_C.shift_reg[351] ;
 wire \ser_C.shift_reg[352] ;
 wire \ser_C.shift_reg[353] ;
 wire \ser_C.shift_reg[354] ;
 wire \ser_C.shift_reg[355] ;
 wire \ser_C.shift_reg[356] ;
 wire \ser_C.shift_reg[357] ;
 wire \ser_C.shift_reg[358] ;
 wire \ser_C.shift_reg[359] ;
 wire \ser_C.shift_reg[35] ;
 wire \ser_C.shift_reg[360] ;
 wire \ser_C.shift_reg[361] ;
 wire \ser_C.shift_reg[362] ;
 wire \ser_C.shift_reg[363] ;
 wire \ser_C.shift_reg[364] ;
 wire \ser_C.shift_reg[365] ;
 wire \ser_C.shift_reg[366] ;
 wire \ser_C.shift_reg[367] ;
 wire \ser_C.shift_reg[368] ;
 wire \ser_C.shift_reg[369] ;
 wire \ser_C.shift_reg[36] ;
 wire \ser_C.shift_reg[370] ;
 wire \ser_C.shift_reg[371] ;
 wire \ser_C.shift_reg[372] ;
 wire \ser_C.shift_reg[373] ;
 wire \ser_C.shift_reg[374] ;
 wire \ser_C.shift_reg[375] ;
 wire \ser_C.shift_reg[376] ;
 wire \ser_C.shift_reg[377] ;
 wire \ser_C.shift_reg[378] ;
 wire \ser_C.shift_reg[379] ;
 wire \ser_C.shift_reg[37] ;
 wire \ser_C.shift_reg[380] ;
 wire \ser_C.shift_reg[381] ;
 wire \ser_C.shift_reg[382] ;
 wire \ser_C.shift_reg[383] ;
 wire \ser_C.shift_reg[384] ;
 wire \ser_C.shift_reg[385] ;
 wire \ser_C.shift_reg[386] ;
 wire \ser_C.shift_reg[387] ;
 wire \ser_C.shift_reg[388] ;
 wire \ser_C.shift_reg[389] ;
 wire \ser_C.shift_reg[38] ;
 wire \ser_C.shift_reg[390] ;
 wire \ser_C.shift_reg[391] ;
 wire \ser_C.shift_reg[392] ;
 wire \ser_C.shift_reg[393] ;
 wire \ser_C.shift_reg[394] ;
 wire \ser_C.shift_reg[395] ;
 wire \ser_C.shift_reg[396] ;
 wire \ser_C.shift_reg[397] ;
 wire \ser_C.shift_reg[398] ;
 wire \ser_C.shift_reg[399] ;
 wire \ser_C.shift_reg[39] ;
 wire \ser_C.shift_reg[3] ;
 wire \ser_C.shift_reg[400] ;
 wire \ser_C.shift_reg[401] ;
 wire \ser_C.shift_reg[402] ;
 wire \ser_C.shift_reg[403] ;
 wire \ser_C.shift_reg[404] ;
 wire \ser_C.shift_reg[405] ;
 wire \ser_C.shift_reg[406] ;
 wire \ser_C.shift_reg[407] ;
 wire \ser_C.shift_reg[408] ;
 wire \ser_C.shift_reg[409] ;
 wire \ser_C.shift_reg[40] ;
 wire \ser_C.shift_reg[410] ;
 wire \ser_C.shift_reg[411] ;
 wire \ser_C.shift_reg[412] ;
 wire \ser_C.shift_reg[413] ;
 wire \ser_C.shift_reg[414] ;
 wire \ser_C.shift_reg[415] ;
 wire \ser_C.shift_reg[416] ;
 wire \ser_C.shift_reg[417] ;
 wire \ser_C.shift_reg[418] ;
 wire \ser_C.shift_reg[419] ;
 wire \ser_C.shift_reg[41] ;
 wire \ser_C.shift_reg[420] ;
 wire \ser_C.shift_reg[421] ;
 wire \ser_C.shift_reg[422] ;
 wire \ser_C.shift_reg[423] ;
 wire \ser_C.shift_reg[424] ;
 wire \ser_C.shift_reg[425] ;
 wire \ser_C.shift_reg[426] ;
 wire \ser_C.shift_reg[427] ;
 wire \ser_C.shift_reg[428] ;
 wire \ser_C.shift_reg[429] ;
 wire \ser_C.shift_reg[42] ;
 wire \ser_C.shift_reg[430] ;
 wire \ser_C.shift_reg[431] ;
 wire \ser_C.shift_reg[432] ;
 wire \ser_C.shift_reg[433] ;
 wire \ser_C.shift_reg[434] ;
 wire \ser_C.shift_reg[435] ;
 wire \ser_C.shift_reg[436] ;
 wire \ser_C.shift_reg[437] ;
 wire \ser_C.shift_reg[438] ;
 wire \ser_C.shift_reg[439] ;
 wire \ser_C.shift_reg[43] ;
 wire \ser_C.shift_reg[440] ;
 wire \ser_C.shift_reg[441] ;
 wire \ser_C.shift_reg[442] ;
 wire \ser_C.shift_reg[443] ;
 wire \ser_C.shift_reg[444] ;
 wire \ser_C.shift_reg[445] ;
 wire \ser_C.shift_reg[446] ;
 wire \ser_C.shift_reg[447] ;
 wire \ser_C.shift_reg[448] ;
 wire \ser_C.shift_reg[449] ;
 wire \ser_C.shift_reg[44] ;
 wire \ser_C.shift_reg[450] ;
 wire \ser_C.shift_reg[451] ;
 wire \ser_C.shift_reg[452] ;
 wire \ser_C.shift_reg[453] ;
 wire \ser_C.shift_reg[454] ;
 wire \ser_C.shift_reg[455] ;
 wire \ser_C.shift_reg[456] ;
 wire \ser_C.shift_reg[457] ;
 wire \ser_C.shift_reg[458] ;
 wire \ser_C.shift_reg[459] ;
 wire \ser_C.shift_reg[45] ;
 wire \ser_C.shift_reg[460] ;
 wire \ser_C.shift_reg[461] ;
 wire \ser_C.shift_reg[462] ;
 wire \ser_C.shift_reg[463] ;
 wire \ser_C.shift_reg[464] ;
 wire \ser_C.shift_reg[465] ;
 wire \ser_C.shift_reg[466] ;
 wire \ser_C.shift_reg[467] ;
 wire \ser_C.shift_reg[468] ;
 wire \ser_C.shift_reg[469] ;
 wire \ser_C.shift_reg[46] ;
 wire \ser_C.shift_reg[470] ;
 wire \ser_C.shift_reg[471] ;
 wire \ser_C.shift_reg[472] ;
 wire \ser_C.shift_reg[473] ;
 wire \ser_C.shift_reg[474] ;
 wire \ser_C.shift_reg[475] ;
 wire \ser_C.shift_reg[476] ;
 wire \ser_C.shift_reg[477] ;
 wire \ser_C.shift_reg[478] ;
 wire \ser_C.shift_reg[479] ;
 wire \ser_C.shift_reg[47] ;
 wire \ser_C.shift_reg[480] ;
 wire \ser_C.shift_reg[481] ;
 wire \ser_C.shift_reg[482] ;
 wire \ser_C.shift_reg[483] ;
 wire \ser_C.shift_reg[484] ;
 wire \ser_C.shift_reg[485] ;
 wire \ser_C.shift_reg[486] ;
 wire \ser_C.shift_reg[487] ;
 wire \ser_C.shift_reg[488] ;
 wire \ser_C.shift_reg[489] ;
 wire \ser_C.shift_reg[48] ;
 wire \ser_C.shift_reg[490] ;
 wire \ser_C.shift_reg[491] ;
 wire \ser_C.shift_reg[492] ;
 wire \ser_C.shift_reg[493] ;
 wire \ser_C.shift_reg[494] ;
 wire \ser_C.shift_reg[495] ;
 wire \ser_C.shift_reg[496] ;
 wire \ser_C.shift_reg[497] ;
 wire \ser_C.shift_reg[498] ;
 wire \ser_C.shift_reg[499] ;
 wire \ser_C.shift_reg[49] ;
 wire \ser_C.shift_reg[4] ;
 wire \ser_C.shift_reg[500] ;
 wire \ser_C.shift_reg[501] ;
 wire \ser_C.shift_reg[502] ;
 wire \ser_C.shift_reg[503] ;
 wire \ser_C.shift_reg[504] ;
 wire \ser_C.shift_reg[505] ;
 wire \ser_C.shift_reg[506] ;
 wire \ser_C.shift_reg[507] ;
 wire \ser_C.shift_reg[508] ;
 wire \ser_C.shift_reg[509] ;
 wire \ser_C.shift_reg[50] ;
 wire \ser_C.shift_reg[510] ;
 wire \ser_C.shift_reg[511] ;
 wire \ser_C.shift_reg[51] ;
 wire \ser_C.shift_reg[52] ;
 wire \ser_C.shift_reg[53] ;
 wire \ser_C.shift_reg[54] ;
 wire \ser_C.shift_reg[55] ;
 wire \ser_C.shift_reg[56] ;
 wire \ser_C.shift_reg[57] ;
 wire \ser_C.shift_reg[58] ;
 wire \ser_C.shift_reg[59] ;
 wire \ser_C.shift_reg[5] ;
 wire \ser_C.shift_reg[60] ;
 wire \ser_C.shift_reg[61] ;
 wire \ser_C.shift_reg[62] ;
 wire \ser_C.shift_reg[63] ;
 wire \ser_C.shift_reg[64] ;
 wire \ser_C.shift_reg[65] ;
 wire \ser_C.shift_reg[66] ;
 wire \ser_C.shift_reg[67] ;
 wire \ser_C.shift_reg[68] ;
 wire \ser_C.shift_reg[69] ;
 wire \ser_C.shift_reg[6] ;
 wire \ser_C.shift_reg[70] ;
 wire \ser_C.shift_reg[71] ;
 wire \ser_C.shift_reg[72] ;
 wire \ser_C.shift_reg[73] ;
 wire \ser_C.shift_reg[74] ;
 wire \ser_C.shift_reg[75] ;
 wire \ser_C.shift_reg[76] ;
 wire \ser_C.shift_reg[77] ;
 wire \ser_C.shift_reg[78] ;
 wire \ser_C.shift_reg[79] ;
 wire \ser_C.shift_reg[7] ;
 wire \ser_C.shift_reg[80] ;
 wire \ser_C.shift_reg[81] ;
 wire \ser_C.shift_reg[82] ;
 wire \ser_C.shift_reg[83] ;
 wire \ser_C.shift_reg[84] ;
 wire \ser_C.shift_reg[85] ;
 wire \ser_C.shift_reg[86] ;
 wire \ser_C.shift_reg[87] ;
 wire \ser_C.shift_reg[88] ;
 wire \ser_C.shift_reg[89] ;
 wire \ser_C.shift_reg[8] ;
 wire \ser_C.shift_reg[90] ;
 wire \ser_C.shift_reg[91] ;
 wire \ser_C.shift_reg[92] ;
 wire \ser_C.shift_reg[93] ;
 wire \ser_C.shift_reg[94] ;
 wire \ser_C.shift_reg[95] ;
 wire \ser_C.shift_reg[96] ;
 wire \ser_C.shift_reg[97] ;
 wire \ser_C.shift_reg[98] ;
 wire \ser_C.shift_reg[99] ;
 wire \ser_C.shift_reg[9] ;
 wire \systolic_inst.A_outs[0][0] ;
 wire \systolic_inst.A_outs[0][1] ;
 wire \systolic_inst.A_outs[0][2] ;
 wire \systolic_inst.A_outs[0][3] ;
 wire \systolic_inst.A_outs[0][4] ;
 wire \systolic_inst.A_outs[0][5] ;
 wire \systolic_inst.A_outs[0][6] ;
 wire \systolic_inst.A_outs[0][7] ;
 wire \systolic_inst.A_outs[10][0] ;
 wire \systolic_inst.A_outs[10][1] ;
 wire \systolic_inst.A_outs[10][2] ;
 wire \systolic_inst.A_outs[10][3] ;
 wire \systolic_inst.A_outs[10][4] ;
 wire \systolic_inst.A_outs[10][5] ;
 wire \systolic_inst.A_outs[10][6] ;
 wire \systolic_inst.A_outs[10][7] ;
 wire \systolic_inst.A_outs[11][0] ;
 wire \systolic_inst.A_outs[11][1] ;
 wire \systolic_inst.A_outs[11][2] ;
 wire \systolic_inst.A_outs[11][3] ;
 wire \systolic_inst.A_outs[11][4] ;
 wire \systolic_inst.A_outs[11][5] ;
 wire \systolic_inst.A_outs[11][6] ;
 wire \systolic_inst.A_outs[11][7] ;
 wire \systolic_inst.A_outs[12][0] ;
 wire \systolic_inst.A_outs[12][1] ;
 wire \systolic_inst.A_outs[12][2] ;
 wire \systolic_inst.A_outs[12][3] ;
 wire \systolic_inst.A_outs[12][4] ;
 wire \systolic_inst.A_outs[12][5] ;
 wire \systolic_inst.A_outs[12][6] ;
 wire \systolic_inst.A_outs[12][7] ;
 wire \systolic_inst.A_outs[13][0] ;
 wire \systolic_inst.A_outs[13][1] ;
 wire \systolic_inst.A_outs[13][2] ;
 wire \systolic_inst.A_outs[13][3] ;
 wire \systolic_inst.A_outs[13][4] ;
 wire \systolic_inst.A_outs[13][5] ;
 wire \systolic_inst.A_outs[13][6] ;
 wire \systolic_inst.A_outs[13][7] ;
 wire \systolic_inst.A_outs[14][0] ;
 wire \systolic_inst.A_outs[14][1] ;
 wire \systolic_inst.A_outs[14][2] ;
 wire \systolic_inst.A_outs[14][3] ;
 wire \systolic_inst.A_outs[14][4] ;
 wire \systolic_inst.A_outs[14][5] ;
 wire \systolic_inst.A_outs[14][6] ;
 wire \systolic_inst.A_outs[14][7] ;
 wire \systolic_inst.A_outs[15][0] ;
 wire \systolic_inst.A_outs[15][1] ;
 wire \systolic_inst.A_outs[15][2] ;
 wire \systolic_inst.A_outs[15][3] ;
 wire \systolic_inst.A_outs[15][4] ;
 wire \systolic_inst.A_outs[15][5] ;
 wire \systolic_inst.A_outs[15][6] ;
 wire \systolic_inst.A_outs[15][7] ;
 wire \systolic_inst.A_outs[1][0] ;
 wire \systolic_inst.A_outs[1][1] ;
 wire \systolic_inst.A_outs[1][2] ;
 wire \systolic_inst.A_outs[1][3] ;
 wire \systolic_inst.A_outs[1][4] ;
 wire \systolic_inst.A_outs[1][5] ;
 wire \systolic_inst.A_outs[1][6] ;
 wire \systolic_inst.A_outs[1][7] ;
 wire \systolic_inst.A_outs[2][0] ;
 wire \systolic_inst.A_outs[2][1] ;
 wire \systolic_inst.A_outs[2][2] ;
 wire \systolic_inst.A_outs[2][3] ;
 wire \systolic_inst.A_outs[2][4] ;
 wire \systolic_inst.A_outs[2][5] ;
 wire \systolic_inst.A_outs[2][6] ;
 wire \systolic_inst.A_outs[2][7] ;
 wire \systolic_inst.A_outs[3][0] ;
 wire \systolic_inst.A_outs[3][1] ;
 wire \systolic_inst.A_outs[3][2] ;
 wire \systolic_inst.A_outs[3][3] ;
 wire \systolic_inst.A_outs[3][4] ;
 wire \systolic_inst.A_outs[3][5] ;
 wire \systolic_inst.A_outs[3][6] ;
 wire \systolic_inst.A_outs[3][7] ;
 wire \systolic_inst.A_outs[4][0] ;
 wire \systolic_inst.A_outs[4][1] ;
 wire \systolic_inst.A_outs[4][2] ;
 wire \systolic_inst.A_outs[4][3] ;
 wire \systolic_inst.A_outs[4][4] ;
 wire \systolic_inst.A_outs[4][5] ;
 wire \systolic_inst.A_outs[4][6] ;
 wire \systolic_inst.A_outs[4][7] ;
 wire \systolic_inst.A_outs[5][0] ;
 wire \systolic_inst.A_outs[5][1] ;
 wire \systolic_inst.A_outs[5][2] ;
 wire \systolic_inst.A_outs[5][3] ;
 wire \systolic_inst.A_outs[5][4] ;
 wire \systolic_inst.A_outs[5][5] ;
 wire \systolic_inst.A_outs[5][6] ;
 wire \systolic_inst.A_outs[5][7] ;
 wire \systolic_inst.A_outs[6][0] ;
 wire \systolic_inst.A_outs[6][1] ;
 wire \systolic_inst.A_outs[6][2] ;
 wire \systolic_inst.A_outs[6][3] ;
 wire \systolic_inst.A_outs[6][4] ;
 wire \systolic_inst.A_outs[6][5] ;
 wire \systolic_inst.A_outs[6][6] ;
 wire \systolic_inst.A_outs[6][7] ;
 wire \systolic_inst.A_outs[7][0] ;
 wire \systolic_inst.A_outs[7][1] ;
 wire \systolic_inst.A_outs[7][2] ;
 wire \systolic_inst.A_outs[7][3] ;
 wire \systolic_inst.A_outs[7][4] ;
 wire \systolic_inst.A_outs[7][5] ;
 wire \systolic_inst.A_outs[7][6] ;
 wire \systolic_inst.A_outs[7][7] ;
 wire \systolic_inst.A_outs[8][0] ;
 wire \systolic_inst.A_outs[8][1] ;
 wire \systolic_inst.A_outs[8][2] ;
 wire \systolic_inst.A_outs[8][3] ;
 wire \systolic_inst.A_outs[8][4] ;
 wire \systolic_inst.A_outs[8][5] ;
 wire \systolic_inst.A_outs[8][6] ;
 wire \systolic_inst.A_outs[8][7] ;
 wire \systolic_inst.A_outs[9][0] ;
 wire \systolic_inst.A_outs[9][1] ;
 wire \systolic_inst.A_outs[9][2] ;
 wire \systolic_inst.A_outs[9][3] ;
 wire \systolic_inst.A_outs[9][4] ;
 wire \systolic_inst.A_outs[9][5] ;
 wire \systolic_inst.A_outs[9][6] ;
 wire \systolic_inst.A_outs[9][7] ;
 wire \systolic_inst.A_shift[0][0] ;
 wire \systolic_inst.A_shift[0][1] ;
 wire \systolic_inst.A_shift[0][2] ;
 wire \systolic_inst.A_shift[0][3] ;
 wire \systolic_inst.A_shift[0][4] ;
 wire \systolic_inst.A_shift[0][5] ;
 wire \systolic_inst.A_shift[0][6] ;
 wire \systolic_inst.A_shift[0][7] ;
 wire \systolic_inst.A_shift[10][0] ;
 wire \systolic_inst.A_shift[10][1] ;
 wire \systolic_inst.A_shift[10][2] ;
 wire \systolic_inst.A_shift[10][3] ;
 wire \systolic_inst.A_shift[10][4] ;
 wire \systolic_inst.A_shift[10][5] ;
 wire \systolic_inst.A_shift[10][6] ;
 wire \systolic_inst.A_shift[10][7] ;
 wire \systolic_inst.A_shift[11][0] ;
 wire \systolic_inst.A_shift[11][1] ;
 wire \systolic_inst.A_shift[11][2] ;
 wire \systolic_inst.A_shift[11][3] ;
 wire \systolic_inst.A_shift[11][4] ;
 wire \systolic_inst.A_shift[11][5] ;
 wire \systolic_inst.A_shift[11][6] ;
 wire \systolic_inst.A_shift[11][7] ;
 wire \systolic_inst.A_shift[12][0] ;
 wire \systolic_inst.A_shift[12][1] ;
 wire \systolic_inst.A_shift[12][2] ;
 wire \systolic_inst.A_shift[12][3] ;
 wire \systolic_inst.A_shift[12][4] ;
 wire \systolic_inst.A_shift[12][5] ;
 wire \systolic_inst.A_shift[12][6] ;
 wire \systolic_inst.A_shift[12][7] ;
 wire \systolic_inst.A_shift[16][0] ;
 wire \systolic_inst.A_shift[16][1] ;
 wire \systolic_inst.A_shift[16][2] ;
 wire \systolic_inst.A_shift[16][3] ;
 wire \systolic_inst.A_shift[16][4] ;
 wire \systolic_inst.A_shift[16][5] ;
 wire \systolic_inst.A_shift[16][6] ;
 wire \systolic_inst.A_shift[16][7] ;
 wire \systolic_inst.A_shift[17][0] ;
 wire \systolic_inst.A_shift[17][1] ;
 wire \systolic_inst.A_shift[17][2] ;
 wire \systolic_inst.A_shift[17][3] ;
 wire \systolic_inst.A_shift[17][4] ;
 wire \systolic_inst.A_shift[17][5] ;
 wire \systolic_inst.A_shift[17][6] ;
 wire \systolic_inst.A_shift[17][7] ;
 wire \systolic_inst.A_shift[18][0] ;
 wire \systolic_inst.A_shift[18][1] ;
 wire \systolic_inst.A_shift[18][2] ;
 wire \systolic_inst.A_shift[18][3] ;
 wire \systolic_inst.A_shift[18][4] ;
 wire \systolic_inst.A_shift[18][5] ;
 wire \systolic_inst.A_shift[18][6] ;
 wire \systolic_inst.A_shift[18][7] ;
 wire \systolic_inst.A_shift[19][0] ;
 wire \systolic_inst.A_shift[19][1] ;
 wire \systolic_inst.A_shift[19][2] ;
 wire \systolic_inst.A_shift[19][3] ;
 wire \systolic_inst.A_shift[19][4] ;
 wire \systolic_inst.A_shift[19][5] ;
 wire \systolic_inst.A_shift[19][6] ;
 wire \systolic_inst.A_shift[19][7] ;
 wire \systolic_inst.A_shift[1][0] ;
 wire \systolic_inst.A_shift[1][1] ;
 wire \systolic_inst.A_shift[1][2] ;
 wire \systolic_inst.A_shift[1][3] ;
 wire \systolic_inst.A_shift[1][4] ;
 wire \systolic_inst.A_shift[1][5] ;
 wire \systolic_inst.A_shift[1][6] ;
 wire \systolic_inst.A_shift[1][7] ;
 wire \systolic_inst.A_shift[20][0] ;
 wire \systolic_inst.A_shift[20][1] ;
 wire \systolic_inst.A_shift[20][2] ;
 wire \systolic_inst.A_shift[20][3] ;
 wire \systolic_inst.A_shift[20][4] ;
 wire \systolic_inst.A_shift[20][5] ;
 wire \systolic_inst.A_shift[20][6] ;
 wire \systolic_inst.A_shift[20][7] ;
 wire \systolic_inst.A_shift[21][0] ;
 wire \systolic_inst.A_shift[21][1] ;
 wire \systolic_inst.A_shift[21][2] ;
 wire \systolic_inst.A_shift[21][3] ;
 wire \systolic_inst.A_shift[21][4] ;
 wire \systolic_inst.A_shift[21][5] ;
 wire \systolic_inst.A_shift[21][6] ;
 wire \systolic_inst.A_shift[21][7] ;
 wire \systolic_inst.A_shift[24][0] ;
 wire \systolic_inst.A_shift[24][1] ;
 wire \systolic_inst.A_shift[24][2] ;
 wire \systolic_inst.A_shift[24][3] ;
 wire \systolic_inst.A_shift[24][4] ;
 wire \systolic_inst.A_shift[24][5] ;
 wire \systolic_inst.A_shift[24][6] ;
 wire \systolic_inst.A_shift[24][7] ;
 wire \systolic_inst.A_shift[25][0] ;
 wire \systolic_inst.A_shift[25][1] ;
 wire \systolic_inst.A_shift[25][2] ;
 wire \systolic_inst.A_shift[25][3] ;
 wire \systolic_inst.A_shift[25][4] ;
 wire \systolic_inst.A_shift[25][5] ;
 wire \systolic_inst.A_shift[25][6] ;
 wire \systolic_inst.A_shift[25][7] ;
 wire \systolic_inst.A_shift[26][0] ;
 wire \systolic_inst.A_shift[26][1] ;
 wire \systolic_inst.A_shift[26][2] ;
 wire \systolic_inst.A_shift[26][3] ;
 wire \systolic_inst.A_shift[26][4] ;
 wire \systolic_inst.A_shift[26][5] ;
 wire \systolic_inst.A_shift[26][6] ;
 wire \systolic_inst.A_shift[26][7] ;
 wire \systolic_inst.A_shift[27][0] ;
 wire \systolic_inst.A_shift[27][1] ;
 wire \systolic_inst.A_shift[27][2] ;
 wire \systolic_inst.A_shift[27][3] ;
 wire \systolic_inst.A_shift[27][4] ;
 wire \systolic_inst.A_shift[27][5] ;
 wire \systolic_inst.A_shift[27][6] ;
 wire \systolic_inst.A_shift[27][7] ;
 wire \systolic_inst.A_shift[28][0] ;
 wire \systolic_inst.A_shift[28][1] ;
 wire \systolic_inst.A_shift[28][2] ;
 wire \systolic_inst.A_shift[28][3] ;
 wire \systolic_inst.A_shift[28][4] ;
 wire \systolic_inst.A_shift[28][5] ;
 wire \systolic_inst.A_shift[28][6] ;
 wire \systolic_inst.A_shift[28][7] ;
 wire \systolic_inst.A_shift[29][0] ;
 wire \systolic_inst.A_shift[29][1] ;
 wire \systolic_inst.A_shift[29][2] ;
 wire \systolic_inst.A_shift[29][3] ;
 wire \systolic_inst.A_shift[29][4] ;
 wire \systolic_inst.A_shift[29][5] ;
 wire \systolic_inst.A_shift[29][6] ;
 wire \systolic_inst.A_shift[29][7] ;
 wire \systolic_inst.A_shift[2][0] ;
 wire \systolic_inst.A_shift[2][1] ;
 wire \systolic_inst.A_shift[2][2] ;
 wire \systolic_inst.A_shift[2][3] ;
 wire \systolic_inst.A_shift[2][4] ;
 wire \systolic_inst.A_shift[2][5] ;
 wire \systolic_inst.A_shift[2][6] ;
 wire \systolic_inst.A_shift[2][7] ;
 wire \systolic_inst.A_shift[30][0] ;
 wire \systolic_inst.A_shift[30][1] ;
 wire \systolic_inst.A_shift[30][2] ;
 wire \systolic_inst.A_shift[30][3] ;
 wire \systolic_inst.A_shift[30][4] ;
 wire \systolic_inst.A_shift[30][5] ;
 wire \systolic_inst.A_shift[30][6] ;
 wire \systolic_inst.A_shift[30][7] ;
 wire \systolic_inst.A_shift[3][0] ;
 wire \systolic_inst.A_shift[3][1] ;
 wire \systolic_inst.A_shift[3][2] ;
 wire \systolic_inst.A_shift[3][3] ;
 wire \systolic_inst.A_shift[3][4] ;
 wire \systolic_inst.A_shift[3][5] ;
 wire \systolic_inst.A_shift[3][6] ;
 wire \systolic_inst.A_shift[3][7] ;
 wire \systolic_inst.A_shift[8][0] ;
 wire \systolic_inst.A_shift[8][1] ;
 wire \systolic_inst.A_shift[8][2] ;
 wire \systolic_inst.A_shift[8][3] ;
 wire \systolic_inst.A_shift[8][4] ;
 wire \systolic_inst.A_shift[8][5] ;
 wire \systolic_inst.A_shift[8][6] ;
 wire \systolic_inst.A_shift[8][7] ;
 wire \systolic_inst.A_shift[9][0] ;
 wire \systolic_inst.A_shift[9][1] ;
 wire \systolic_inst.A_shift[9][2] ;
 wire \systolic_inst.A_shift[9][3] ;
 wire \systolic_inst.A_shift[9][4] ;
 wire \systolic_inst.A_shift[9][5] ;
 wire \systolic_inst.A_shift[9][6] ;
 wire \systolic_inst.A_shift[9][7] ;
 wire \systolic_inst.B_outs[0][0] ;
 wire \systolic_inst.B_outs[0][1] ;
 wire \systolic_inst.B_outs[0][2] ;
 wire \systolic_inst.B_outs[0][3] ;
 wire \systolic_inst.B_outs[0][4] ;
 wire \systolic_inst.B_outs[0][5] ;
 wire \systolic_inst.B_outs[0][6] ;
 wire \systolic_inst.B_outs[0][7] ;
 wire \systolic_inst.B_outs[10][0] ;
 wire \systolic_inst.B_outs[10][1] ;
 wire \systolic_inst.B_outs[10][2] ;
 wire \systolic_inst.B_outs[10][3] ;
 wire \systolic_inst.B_outs[10][4] ;
 wire \systolic_inst.B_outs[10][5] ;
 wire \systolic_inst.B_outs[10][6] ;
 wire \systolic_inst.B_outs[10][7] ;
 wire \systolic_inst.B_outs[11][0] ;
 wire \systolic_inst.B_outs[11][1] ;
 wire \systolic_inst.B_outs[11][2] ;
 wire \systolic_inst.B_outs[11][3] ;
 wire \systolic_inst.B_outs[11][4] ;
 wire \systolic_inst.B_outs[11][5] ;
 wire \systolic_inst.B_outs[11][6] ;
 wire \systolic_inst.B_outs[11][7] ;
 wire \systolic_inst.B_outs[12][0] ;
 wire \systolic_inst.B_outs[12][1] ;
 wire \systolic_inst.B_outs[12][2] ;
 wire \systolic_inst.B_outs[12][3] ;
 wire \systolic_inst.B_outs[12][4] ;
 wire \systolic_inst.B_outs[12][5] ;
 wire \systolic_inst.B_outs[12][6] ;
 wire \systolic_inst.B_outs[12][7] ;
 wire \systolic_inst.B_outs[13][0] ;
 wire \systolic_inst.B_outs[13][1] ;
 wire \systolic_inst.B_outs[13][2] ;
 wire \systolic_inst.B_outs[13][3] ;
 wire \systolic_inst.B_outs[13][4] ;
 wire \systolic_inst.B_outs[13][5] ;
 wire \systolic_inst.B_outs[13][6] ;
 wire \systolic_inst.B_outs[13][7] ;
 wire \systolic_inst.B_outs[14][0] ;
 wire \systolic_inst.B_outs[14][1] ;
 wire \systolic_inst.B_outs[14][2] ;
 wire \systolic_inst.B_outs[14][3] ;
 wire \systolic_inst.B_outs[14][4] ;
 wire \systolic_inst.B_outs[14][5] ;
 wire \systolic_inst.B_outs[14][6] ;
 wire \systolic_inst.B_outs[14][7] ;
 wire \systolic_inst.B_outs[15][0] ;
 wire \systolic_inst.B_outs[15][1] ;
 wire \systolic_inst.B_outs[15][2] ;
 wire \systolic_inst.B_outs[15][3] ;
 wire \systolic_inst.B_outs[15][4] ;
 wire \systolic_inst.B_outs[15][5] ;
 wire \systolic_inst.B_outs[15][6] ;
 wire \systolic_inst.B_outs[15][7] ;
 wire \systolic_inst.B_outs[1][0] ;
 wire \systolic_inst.B_outs[1][1] ;
 wire \systolic_inst.B_outs[1][2] ;
 wire \systolic_inst.B_outs[1][3] ;
 wire \systolic_inst.B_outs[1][4] ;
 wire \systolic_inst.B_outs[1][5] ;
 wire \systolic_inst.B_outs[1][6] ;
 wire \systolic_inst.B_outs[1][7] ;
 wire \systolic_inst.B_outs[2][0] ;
 wire \systolic_inst.B_outs[2][1] ;
 wire \systolic_inst.B_outs[2][2] ;
 wire \systolic_inst.B_outs[2][3] ;
 wire \systolic_inst.B_outs[2][4] ;
 wire \systolic_inst.B_outs[2][5] ;
 wire \systolic_inst.B_outs[2][6] ;
 wire \systolic_inst.B_outs[2][7] ;
 wire \systolic_inst.B_outs[3][0] ;
 wire \systolic_inst.B_outs[3][1] ;
 wire \systolic_inst.B_outs[3][2] ;
 wire \systolic_inst.B_outs[3][3] ;
 wire \systolic_inst.B_outs[3][4] ;
 wire \systolic_inst.B_outs[3][5] ;
 wire \systolic_inst.B_outs[3][6] ;
 wire \systolic_inst.B_outs[3][7] ;
 wire \systolic_inst.B_outs[4][0] ;
 wire \systolic_inst.B_outs[4][1] ;
 wire \systolic_inst.B_outs[4][2] ;
 wire \systolic_inst.B_outs[4][3] ;
 wire \systolic_inst.B_outs[4][4] ;
 wire \systolic_inst.B_outs[4][5] ;
 wire \systolic_inst.B_outs[4][6] ;
 wire \systolic_inst.B_outs[4][7] ;
 wire \systolic_inst.B_outs[5][0] ;
 wire \systolic_inst.B_outs[5][1] ;
 wire \systolic_inst.B_outs[5][2] ;
 wire \systolic_inst.B_outs[5][3] ;
 wire \systolic_inst.B_outs[5][4] ;
 wire \systolic_inst.B_outs[5][5] ;
 wire \systolic_inst.B_outs[5][6] ;
 wire \systolic_inst.B_outs[5][7] ;
 wire \systolic_inst.B_outs[6][0] ;
 wire \systolic_inst.B_outs[6][1] ;
 wire \systolic_inst.B_outs[6][2] ;
 wire \systolic_inst.B_outs[6][3] ;
 wire \systolic_inst.B_outs[6][4] ;
 wire \systolic_inst.B_outs[6][5] ;
 wire \systolic_inst.B_outs[6][6] ;
 wire \systolic_inst.B_outs[6][7] ;
 wire \systolic_inst.B_outs[7][0] ;
 wire \systolic_inst.B_outs[7][1] ;
 wire \systolic_inst.B_outs[7][2] ;
 wire \systolic_inst.B_outs[7][3] ;
 wire \systolic_inst.B_outs[7][4] ;
 wire \systolic_inst.B_outs[7][5] ;
 wire \systolic_inst.B_outs[7][6] ;
 wire \systolic_inst.B_outs[7][7] ;
 wire \systolic_inst.B_outs[8][0] ;
 wire \systolic_inst.B_outs[8][1] ;
 wire \systolic_inst.B_outs[8][2] ;
 wire \systolic_inst.B_outs[8][3] ;
 wire \systolic_inst.B_outs[8][4] ;
 wire \systolic_inst.B_outs[8][5] ;
 wire \systolic_inst.B_outs[8][6] ;
 wire \systolic_inst.B_outs[8][7] ;
 wire \systolic_inst.B_outs[9][0] ;
 wire \systolic_inst.B_outs[9][1] ;
 wire \systolic_inst.B_outs[9][2] ;
 wire \systolic_inst.B_outs[9][3] ;
 wire \systolic_inst.B_outs[9][4] ;
 wire \systolic_inst.B_outs[9][5] ;
 wire \systolic_inst.B_outs[9][6] ;
 wire \systolic_inst.B_outs[9][7] ;
 wire \systolic_inst.B_shift[0][0] ;
 wire \systolic_inst.B_shift[0][1] ;
 wire \systolic_inst.B_shift[0][2] ;
 wire \systolic_inst.B_shift[0][3] ;
 wire \systolic_inst.B_shift[0][4] ;
 wire \systolic_inst.B_shift[0][5] ;
 wire \systolic_inst.B_shift[0][6] ;
 wire \systolic_inst.B_shift[0][7] ;
 wire \systolic_inst.B_shift[10][0] ;
 wire \systolic_inst.B_shift[10][1] ;
 wire \systolic_inst.B_shift[10][2] ;
 wire \systolic_inst.B_shift[10][3] ;
 wire \systolic_inst.B_shift[10][4] ;
 wire \systolic_inst.B_shift[10][5] ;
 wire \systolic_inst.B_shift[10][6] ;
 wire \systolic_inst.B_shift[10][7] ;
 wire \systolic_inst.B_shift[11][0] ;
 wire \systolic_inst.B_shift[11][1] ;
 wire \systolic_inst.B_shift[11][2] ;
 wire \systolic_inst.B_shift[11][3] ;
 wire \systolic_inst.B_shift[11][4] ;
 wire \systolic_inst.B_shift[11][5] ;
 wire \systolic_inst.B_shift[11][6] ;
 wire \systolic_inst.B_shift[11][7] ;
 wire \systolic_inst.B_shift[12][0] ;
 wire \systolic_inst.B_shift[12][1] ;
 wire \systolic_inst.B_shift[12][2] ;
 wire \systolic_inst.B_shift[12][3] ;
 wire \systolic_inst.B_shift[12][4] ;
 wire \systolic_inst.B_shift[12][5] ;
 wire \systolic_inst.B_shift[12][6] ;
 wire \systolic_inst.B_shift[12][7] ;
 wire \systolic_inst.B_shift[13][0] ;
 wire \systolic_inst.B_shift[13][1] ;
 wire \systolic_inst.B_shift[13][2] ;
 wire \systolic_inst.B_shift[13][3] ;
 wire \systolic_inst.B_shift[13][4] ;
 wire \systolic_inst.B_shift[13][5] ;
 wire \systolic_inst.B_shift[13][6] ;
 wire \systolic_inst.B_shift[13][7] ;
 wire \systolic_inst.B_shift[14][0] ;
 wire \systolic_inst.B_shift[14][1] ;
 wire \systolic_inst.B_shift[14][2] ;
 wire \systolic_inst.B_shift[14][3] ;
 wire \systolic_inst.B_shift[14][4] ;
 wire \systolic_inst.B_shift[14][5] ;
 wire \systolic_inst.B_shift[14][6] ;
 wire \systolic_inst.B_shift[14][7] ;
 wire \systolic_inst.B_shift[15][0] ;
 wire \systolic_inst.B_shift[15][1] ;
 wire \systolic_inst.B_shift[15][2] ;
 wire \systolic_inst.B_shift[15][3] ;
 wire \systolic_inst.B_shift[15][4] ;
 wire \systolic_inst.B_shift[15][5] ;
 wire \systolic_inst.B_shift[15][6] ;
 wire \systolic_inst.B_shift[15][7] ;
 wire \systolic_inst.B_shift[17][0] ;
 wire \systolic_inst.B_shift[17][1] ;
 wire \systolic_inst.B_shift[17][2] ;
 wire \systolic_inst.B_shift[17][3] ;
 wire \systolic_inst.B_shift[17][4] ;
 wire \systolic_inst.B_shift[17][5] ;
 wire \systolic_inst.B_shift[17][6] ;
 wire \systolic_inst.B_shift[17][7] ;
 wire \systolic_inst.B_shift[18][0] ;
 wire \systolic_inst.B_shift[18][1] ;
 wire \systolic_inst.B_shift[18][2] ;
 wire \systolic_inst.B_shift[18][3] ;
 wire \systolic_inst.B_shift[18][4] ;
 wire \systolic_inst.B_shift[18][5] ;
 wire \systolic_inst.B_shift[18][6] ;
 wire \systolic_inst.B_shift[18][7] ;
 wire \systolic_inst.B_shift[19][0] ;
 wire \systolic_inst.B_shift[19][1] ;
 wire \systolic_inst.B_shift[19][2] ;
 wire \systolic_inst.B_shift[19][3] ;
 wire \systolic_inst.B_shift[19][4] ;
 wire \systolic_inst.B_shift[19][5] ;
 wire \systolic_inst.B_shift[19][6] ;
 wire \systolic_inst.B_shift[19][7] ;
 wire \systolic_inst.B_shift[1][0] ;
 wire \systolic_inst.B_shift[1][1] ;
 wire \systolic_inst.B_shift[1][2] ;
 wire \systolic_inst.B_shift[1][3] ;
 wire \systolic_inst.B_shift[1][4] ;
 wire \systolic_inst.B_shift[1][5] ;
 wire \systolic_inst.B_shift[1][6] ;
 wire \systolic_inst.B_shift[1][7] ;
 wire \systolic_inst.B_shift[22][0] ;
 wire \systolic_inst.B_shift[22][1] ;
 wire \systolic_inst.B_shift[22][2] ;
 wire \systolic_inst.B_shift[22][3] ;
 wire \systolic_inst.B_shift[22][4] ;
 wire \systolic_inst.B_shift[22][5] ;
 wire \systolic_inst.B_shift[22][6] ;
 wire \systolic_inst.B_shift[22][7] ;
 wire \systolic_inst.B_shift[23][0] ;
 wire \systolic_inst.B_shift[23][1] ;
 wire \systolic_inst.B_shift[23][2] ;
 wire \systolic_inst.B_shift[23][3] ;
 wire \systolic_inst.B_shift[23][4] ;
 wire \systolic_inst.B_shift[23][5] ;
 wire \systolic_inst.B_shift[23][6] ;
 wire \systolic_inst.B_shift[23][7] ;
 wire \systolic_inst.B_shift[27][0] ;
 wire \systolic_inst.B_shift[27][1] ;
 wire \systolic_inst.B_shift[27][2] ;
 wire \systolic_inst.B_shift[27][3] ;
 wire \systolic_inst.B_shift[27][4] ;
 wire \systolic_inst.B_shift[27][5] ;
 wire \systolic_inst.B_shift[27][6] ;
 wire \systolic_inst.B_shift[27][7] ;
 wire \systolic_inst.B_shift[2][0] ;
 wire \systolic_inst.B_shift[2][1] ;
 wire \systolic_inst.B_shift[2][2] ;
 wire \systolic_inst.B_shift[2][3] ;
 wire \systolic_inst.B_shift[2][4] ;
 wire \systolic_inst.B_shift[2][5] ;
 wire \systolic_inst.B_shift[2][6] ;
 wire \systolic_inst.B_shift[2][7] ;
 wire \systolic_inst.B_shift[3][0] ;
 wire \systolic_inst.B_shift[3][1] ;
 wire \systolic_inst.B_shift[3][2] ;
 wire \systolic_inst.B_shift[3][3] ;
 wire \systolic_inst.B_shift[3][4] ;
 wire \systolic_inst.B_shift[3][5] ;
 wire \systolic_inst.B_shift[3][6] ;
 wire \systolic_inst.B_shift[3][7] ;
 wire \systolic_inst.B_shift[4][0] ;
 wire \systolic_inst.B_shift[4][1] ;
 wire \systolic_inst.B_shift[4][2] ;
 wire \systolic_inst.B_shift[4][3] ;
 wire \systolic_inst.B_shift[4][4] ;
 wire \systolic_inst.B_shift[4][5] ;
 wire \systolic_inst.B_shift[4][6] ;
 wire \systolic_inst.B_shift[4][7] ;
 wire \systolic_inst.B_shift[5][0] ;
 wire \systolic_inst.B_shift[5][1] ;
 wire \systolic_inst.B_shift[5][2] ;
 wire \systolic_inst.B_shift[5][3] ;
 wire \systolic_inst.B_shift[5][4] ;
 wire \systolic_inst.B_shift[5][5] ;
 wire \systolic_inst.B_shift[5][6] ;
 wire \systolic_inst.B_shift[5][7] ;
 wire \systolic_inst.B_shift[6][0] ;
 wire \systolic_inst.B_shift[6][1] ;
 wire \systolic_inst.B_shift[6][2] ;
 wire \systolic_inst.B_shift[6][3] ;
 wire \systolic_inst.B_shift[6][4] ;
 wire \systolic_inst.B_shift[6][5] ;
 wire \systolic_inst.B_shift[6][6] ;
 wire \systolic_inst.B_shift[6][7] ;
 wire \systolic_inst.B_shift[7][0] ;
 wire \systolic_inst.B_shift[7][1] ;
 wire \systolic_inst.B_shift[7][2] ;
 wire \systolic_inst.B_shift[7][3] ;
 wire \systolic_inst.B_shift[7][4] ;
 wire \systolic_inst.B_shift[7][5] ;
 wire \systolic_inst.B_shift[7][6] ;
 wire \systolic_inst.B_shift[7][7] ;
 wire \systolic_inst.B_shift[8][0] ;
 wire \systolic_inst.B_shift[8][1] ;
 wire \systolic_inst.B_shift[8][2] ;
 wire \systolic_inst.B_shift[8][3] ;
 wire \systolic_inst.B_shift[8][4] ;
 wire \systolic_inst.B_shift[8][5] ;
 wire \systolic_inst.B_shift[8][6] ;
 wire \systolic_inst.B_shift[8][7] ;
 wire \systolic_inst.B_shift[9][0] ;
 wire \systolic_inst.B_shift[9][1] ;
 wire \systolic_inst.B_shift[9][2] ;
 wire \systolic_inst.B_shift[9][3] ;
 wire \systolic_inst.B_shift[9][4] ;
 wire \systolic_inst.B_shift[9][5] ;
 wire \systolic_inst.B_shift[9][6] ;
 wire \systolic_inst.B_shift[9][7] ;
 wire \systolic_inst.acc_wires[0][0] ;
 wire \systolic_inst.acc_wires[0][10] ;
 wire \systolic_inst.acc_wires[0][11] ;
 wire \systolic_inst.acc_wires[0][12] ;
 wire \systolic_inst.acc_wires[0][13] ;
 wire \systolic_inst.acc_wires[0][14] ;
 wire \systolic_inst.acc_wires[0][15] ;
 wire \systolic_inst.acc_wires[0][16] ;
 wire \systolic_inst.acc_wires[0][17] ;
 wire \systolic_inst.acc_wires[0][18] ;
 wire \systolic_inst.acc_wires[0][19] ;
 wire \systolic_inst.acc_wires[0][1] ;
 wire \systolic_inst.acc_wires[0][20] ;
 wire \systolic_inst.acc_wires[0][21] ;
 wire \systolic_inst.acc_wires[0][22] ;
 wire \systolic_inst.acc_wires[0][23] ;
 wire \systolic_inst.acc_wires[0][24] ;
 wire \systolic_inst.acc_wires[0][25] ;
 wire \systolic_inst.acc_wires[0][26] ;
 wire \systolic_inst.acc_wires[0][27] ;
 wire \systolic_inst.acc_wires[0][28] ;
 wire \systolic_inst.acc_wires[0][29] ;
 wire \systolic_inst.acc_wires[0][2] ;
 wire \systolic_inst.acc_wires[0][30] ;
 wire \systolic_inst.acc_wires[0][31] ;
 wire \systolic_inst.acc_wires[0][3] ;
 wire \systolic_inst.acc_wires[0][4] ;
 wire \systolic_inst.acc_wires[0][5] ;
 wire \systolic_inst.acc_wires[0][6] ;
 wire \systolic_inst.acc_wires[0][7] ;
 wire \systolic_inst.acc_wires[0][8] ;
 wire \systolic_inst.acc_wires[0][9] ;
 wire \systolic_inst.acc_wires[10][0] ;
 wire \systolic_inst.acc_wires[10][10] ;
 wire \systolic_inst.acc_wires[10][11] ;
 wire \systolic_inst.acc_wires[10][12] ;
 wire \systolic_inst.acc_wires[10][13] ;
 wire \systolic_inst.acc_wires[10][14] ;
 wire \systolic_inst.acc_wires[10][15] ;
 wire \systolic_inst.acc_wires[10][16] ;
 wire \systolic_inst.acc_wires[10][17] ;
 wire \systolic_inst.acc_wires[10][18] ;
 wire \systolic_inst.acc_wires[10][19] ;
 wire \systolic_inst.acc_wires[10][1] ;
 wire \systolic_inst.acc_wires[10][20] ;
 wire \systolic_inst.acc_wires[10][21] ;
 wire \systolic_inst.acc_wires[10][22] ;
 wire \systolic_inst.acc_wires[10][23] ;
 wire \systolic_inst.acc_wires[10][24] ;
 wire \systolic_inst.acc_wires[10][25] ;
 wire \systolic_inst.acc_wires[10][26] ;
 wire \systolic_inst.acc_wires[10][27] ;
 wire \systolic_inst.acc_wires[10][28] ;
 wire \systolic_inst.acc_wires[10][29] ;
 wire \systolic_inst.acc_wires[10][2] ;
 wire \systolic_inst.acc_wires[10][30] ;
 wire \systolic_inst.acc_wires[10][31] ;
 wire \systolic_inst.acc_wires[10][3] ;
 wire \systolic_inst.acc_wires[10][4] ;
 wire \systolic_inst.acc_wires[10][5] ;
 wire \systolic_inst.acc_wires[10][6] ;
 wire \systolic_inst.acc_wires[10][7] ;
 wire \systolic_inst.acc_wires[10][8] ;
 wire \systolic_inst.acc_wires[10][9] ;
 wire \systolic_inst.acc_wires[11][0] ;
 wire \systolic_inst.acc_wires[11][10] ;
 wire \systolic_inst.acc_wires[11][11] ;
 wire \systolic_inst.acc_wires[11][12] ;
 wire \systolic_inst.acc_wires[11][13] ;
 wire \systolic_inst.acc_wires[11][14] ;
 wire \systolic_inst.acc_wires[11][15] ;
 wire \systolic_inst.acc_wires[11][16] ;
 wire \systolic_inst.acc_wires[11][17] ;
 wire \systolic_inst.acc_wires[11][18] ;
 wire \systolic_inst.acc_wires[11][19] ;
 wire \systolic_inst.acc_wires[11][1] ;
 wire \systolic_inst.acc_wires[11][20] ;
 wire \systolic_inst.acc_wires[11][21] ;
 wire \systolic_inst.acc_wires[11][22] ;
 wire \systolic_inst.acc_wires[11][23] ;
 wire \systolic_inst.acc_wires[11][24] ;
 wire \systolic_inst.acc_wires[11][25] ;
 wire \systolic_inst.acc_wires[11][26] ;
 wire \systolic_inst.acc_wires[11][27] ;
 wire \systolic_inst.acc_wires[11][28] ;
 wire \systolic_inst.acc_wires[11][29] ;
 wire \systolic_inst.acc_wires[11][2] ;
 wire \systolic_inst.acc_wires[11][30] ;
 wire \systolic_inst.acc_wires[11][31] ;
 wire \systolic_inst.acc_wires[11][3] ;
 wire \systolic_inst.acc_wires[11][4] ;
 wire \systolic_inst.acc_wires[11][5] ;
 wire \systolic_inst.acc_wires[11][6] ;
 wire \systolic_inst.acc_wires[11][7] ;
 wire \systolic_inst.acc_wires[11][8] ;
 wire \systolic_inst.acc_wires[11][9] ;
 wire \systolic_inst.acc_wires[12][0] ;
 wire \systolic_inst.acc_wires[12][10] ;
 wire \systolic_inst.acc_wires[12][11] ;
 wire \systolic_inst.acc_wires[12][12] ;
 wire \systolic_inst.acc_wires[12][13] ;
 wire \systolic_inst.acc_wires[12][14] ;
 wire \systolic_inst.acc_wires[12][15] ;
 wire \systolic_inst.acc_wires[12][16] ;
 wire \systolic_inst.acc_wires[12][17] ;
 wire \systolic_inst.acc_wires[12][18] ;
 wire \systolic_inst.acc_wires[12][19] ;
 wire \systolic_inst.acc_wires[12][1] ;
 wire \systolic_inst.acc_wires[12][20] ;
 wire \systolic_inst.acc_wires[12][21] ;
 wire \systolic_inst.acc_wires[12][22] ;
 wire \systolic_inst.acc_wires[12][23] ;
 wire \systolic_inst.acc_wires[12][24] ;
 wire \systolic_inst.acc_wires[12][25] ;
 wire \systolic_inst.acc_wires[12][26] ;
 wire \systolic_inst.acc_wires[12][27] ;
 wire \systolic_inst.acc_wires[12][28] ;
 wire \systolic_inst.acc_wires[12][29] ;
 wire \systolic_inst.acc_wires[12][2] ;
 wire \systolic_inst.acc_wires[12][30] ;
 wire \systolic_inst.acc_wires[12][31] ;
 wire \systolic_inst.acc_wires[12][3] ;
 wire \systolic_inst.acc_wires[12][4] ;
 wire \systolic_inst.acc_wires[12][5] ;
 wire \systolic_inst.acc_wires[12][6] ;
 wire \systolic_inst.acc_wires[12][7] ;
 wire \systolic_inst.acc_wires[12][8] ;
 wire \systolic_inst.acc_wires[12][9] ;
 wire \systolic_inst.acc_wires[13][0] ;
 wire \systolic_inst.acc_wires[13][10] ;
 wire \systolic_inst.acc_wires[13][11] ;
 wire \systolic_inst.acc_wires[13][12] ;
 wire \systolic_inst.acc_wires[13][13] ;
 wire \systolic_inst.acc_wires[13][14] ;
 wire \systolic_inst.acc_wires[13][15] ;
 wire \systolic_inst.acc_wires[13][16] ;
 wire \systolic_inst.acc_wires[13][17] ;
 wire \systolic_inst.acc_wires[13][18] ;
 wire \systolic_inst.acc_wires[13][19] ;
 wire \systolic_inst.acc_wires[13][1] ;
 wire \systolic_inst.acc_wires[13][20] ;
 wire \systolic_inst.acc_wires[13][21] ;
 wire \systolic_inst.acc_wires[13][22] ;
 wire \systolic_inst.acc_wires[13][23] ;
 wire \systolic_inst.acc_wires[13][24] ;
 wire \systolic_inst.acc_wires[13][25] ;
 wire \systolic_inst.acc_wires[13][26] ;
 wire \systolic_inst.acc_wires[13][27] ;
 wire \systolic_inst.acc_wires[13][28] ;
 wire \systolic_inst.acc_wires[13][29] ;
 wire \systolic_inst.acc_wires[13][2] ;
 wire \systolic_inst.acc_wires[13][30] ;
 wire \systolic_inst.acc_wires[13][31] ;
 wire \systolic_inst.acc_wires[13][3] ;
 wire \systolic_inst.acc_wires[13][4] ;
 wire \systolic_inst.acc_wires[13][5] ;
 wire \systolic_inst.acc_wires[13][6] ;
 wire \systolic_inst.acc_wires[13][7] ;
 wire \systolic_inst.acc_wires[13][8] ;
 wire \systolic_inst.acc_wires[13][9] ;
 wire \systolic_inst.acc_wires[14][0] ;
 wire \systolic_inst.acc_wires[14][10] ;
 wire \systolic_inst.acc_wires[14][11] ;
 wire \systolic_inst.acc_wires[14][12] ;
 wire \systolic_inst.acc_wires[14][13] ;
 wire \systolic_inst.acc_wires[14][14] ;
 wire \systolic_inst.acc_wires[14][15] ;
 wire \systolic_inst.acc_wires[14][16] ;
 wire \systolic_inst.acc_wires[14][17] ;
 wire \systolic_inst.acc_wires[14][18] ;
 wire \systolic_inst.acc_wires[14][19] ;
 wire \systolic_inst.acc_wires[14][1] ;
 wire \systolic_inst.acc_wires[14][20] ;
 wire \systolic_inst.acc_wires[14][21] ;
 wire \systolic_inst.acc_wires[14][22] ;
 wire \systolic_inst.acc_wires[14][23] ;
 wire \systolic_inst.acc_wires[14][24] ;
 wire \systolic_inst.acc_wires[14][25] ;
 wire \systolic_inst.acc_wires[14][26] ;
 wire \systolic_inst.acc_wires[14][27] ;
 wire \systolic_inst.acc_wires[14][28] ;
 wire \systolic_inst.acc_wires[14][29] ;
 wire \systolic_inst.acc_wires[14][2] ;
 wire \systolic_inst.acc_wires[14][30] ;
 wire \systolic_inst.acc_wires[14][31] ;
 wire \systolic_inst.acc_wires[14][3] ;
 wire \systolic_inst.acc_wires[14][4] ;
 wire \systolic_inst.acc_wires[14][5] ;
 wire \systolic_inst.acc_wires[14][6] ;
 wire \systolic_inst.acc_wires[14][7] ;
 wire \systolic_inst.acc_wires[14][8] ;
 wire \systolic_inst.acc_wires[14][9] ;
 wire \systolic_inst.acc_wires[15][0] ;
 wire \systolic_inst.acc_wires[15][10] ;
 wire \systolic_inst.acc_wires[15][11] ;
 wire \systolic_inst.acc_wires[15][12] ;
 wire \systolic_inst.acc_wires[15][13] ;
 wire \systolic_inst.acc_wires[15][14] ;
 wire \systolic_inst.acc_wires[15][15] ;
 wire \systolic_inst.acc_wires[15][16] ;
 wire \systolic_inst.acc_wires[15][17] ;
 wire \systolic_inst.acc_wires[15][18] ;
 wire \systolic_inst.acc_wires[15][19] ;
 wire \systolic_inst.acc_wires[15][1] ;
 wire \systolic_inst.acc_wires[15][20] ;
 wire \systolic_inst.acc_wires[15][21] ;
 wire \systolic_inst.acc_wires[15][22] ;
 wire \systolic_inst.acc_wires[15][23] ;
 wire \systolic_inst.acc_wires[15][24] ;
 wire \systolic_inst.acc_wires[15][25] ;
 wire \systolic_inst.acc_wires[15][26] ;
 wire \systolic_inst.acc_wires[15][27] ;
 wire \systolic_inst.acc_wires[15][28] ;
 wire \systolic_inst.acc_wires[15][29] ;
 wire \systolic_inst.acc_wires[15][2] ;
 wire \systolic_inst.acc_wires[15][30] ;
 wire \systolic_inst.acc_wires[15][31] ;
 wire \systolic_inst.acc_wires[15][3] ;
 wire \systolic_inst.acc_wires[15][4] ;
 wire \systolic_inst.acc_wires[15][5] ;
 wire \systolic_inst.acc_wires[15][6] ;
 wire \systolic_inst.acc_wires[15][7] ;
 wire \systolic_inst.acc_wires[15][8] ;
 wire \systolic_inst.acc_wires[15][9] ;
 wire \systolic_inst.acc_wires[1][0] ;
 wire \systolic_inst.acc_wires[1][10] ;
 wire \systolic_inst.acc_wires[1][11] ;
 wire \systolic_inst.acc_wires[1][12] ;
 wire \systolic_inst.acc_wires[1][13] ;
 wire \systolic_inst.acc_wires[1][14] ;
 wire \systolic_inst.acc_wires[1][15] ;
 wire \systolic_inst.acc_wires[1][16] ;
 wire \systolic_inst.acc_wires[1][17] ;
 wire \systolic_inst.acc_wires[1][18] ;
 wire \systolic_inst.acc_wires[1][19] ;
 wire \systolic_inst.acc_wires[1][1] ;
 wire \systolic_inst.acc_wires[1][20] ;
 wire \systolic_inst.acc_wires[1][21] ;
 wire \systolic_inst.acc_wires[1][22] ;
 wire \systolic_inst.acc_wires[1][23] ;
 wire \systolic_inst.acc_wires[1][24] ;
 wire \systolic_inst.acc_wires[1][25] ;
 wire \systolic_inst.acc_wires[1][26] ;
 wire \systolic_inst.acc_wires[1][27] ;
 wire \systolic_inst.acc_wires[1][28] ;
 wire \systolic_inst.acc_wires[1][29] ;
 wire \systolic_inst.acc_wires[1][2] ;
 wire \systolic_inst.acc_wires[1][30] ;
 wire \systolic_inst.acc_wires[1][31] ;
 wire \systolic_inst.acc_wires[1][3] ;
 wire \systolic_inst.acc_wires[1][4] ;
 wire \systolic_inst.acc_wires[1][5] ;
 wire \systolic_inst.acc_wires[1][6] ;
 wire \systolic_inst.acc_wires[1][7] ;
 wire \systolic_inst.acc_wires[1][8] ;
 wire \systolic_inst.acc_wires[1][9] ;
 wire \systolic_inst.acc_wires[2][0] ;
 wire \systolic_inst.acc_wires[2][10] ;
 wire \systolic_inst.acc_wires[2][11] ;
 wire \systolic_inst.acc_wires[2][12] ;
 wire \systolic_inst.acc_wires[2][13] ;
 wire \systolic_inst.acc_wires[2][14] ;
 wire \systolic_inst.acc_wires[2][15] ;
 wire \systolic_inst.acc_wires[2][16] ;
 wire \systolic_inst.acc_wires[2][17] ;
 wire \systolic_inst.acc_wires[2][18] ;
 wire \systolic_inst.acc_wires[2][19] ;
 wire \systolic_inst.acc_wires[2][1] ;
 wire \systolic_inst.acc_wires[2][20] ;
 wire \systolic_inst.acc_wires[2][21] ;
 wire \systolic_inst.acc_wires[2][22] ;
 wire \systolic_inst.acc_wires[2][23] ;
 wire \systolic_inst.acc_wires[2][24] ;
 wire \systolic_inst.acc_wires[2][25] ;
 wire \systolic_inst.acc_wires[2][26] ;
 wire \systolic_inst.acc_wires[2][27] ;
 wire \systolic_inst.acc_wires[2][28] ;
 wire \systolic_inst.acc_wires[2][29] ;
 wire \systolic_inst.acc_wires[2][2] ;
 wire \systolic_inst.acc_wires[2][30] ;
 wire \systolic_inst.acc_wires[2][31] ;
 wire \systolic_inst.acc_wires[2][3] ;
 wire \systolic_inst.acc_wires[2][4] ;
 wire \systolic_inst.acc_wires[2][5] ;
 wire \systolic_inst.acc_wires[2][6] ;
 wire \systolic_inst.acc_wires[2][7] ;
 wire \systolic_inst.acc_wires[2][8] ;
 wire \systolic_inst.acc_wires[2][9] ;
 wire \systolic_inst.acc_wires[3][0] ;
 wire \systolic_inst.acc_wires[3][10] ;
 wire \systolic_inst.acc_wires[3][11] ;
 wire \systolic_inst.acc_wires[3][12] ;
 wire \systolic_inst.acc_wires[3][13] ;
 wire \systolic_inst.acc_wires[3][14] ;
 wire \systolic_inst.acc_wires[3][15] ;
 wire \systolic_inst.acc_wires[3][16] ;
 wire \systolic_inst.acc_wires[3][17] ;
 wire \systolic_inst.acc_wires[3][18] ;
 wire \systolic_inst.acc_wires[3][19] ;
 wire \systolic_inst.acc_wires[3][1] ;
 wire \systolic_inst.acc_wires[3][20] ;
 wire \systolic_inst.acc_wires[3][21] ;
 wire \systolic_inst.acc_wires[3][22] ;
 wire \systolic_inst.acc_wires[3][23] ;
 wire \systolic_inst.acc_wires[3][24] ;
 wire \systolic_inst.acc_wires[3][25] ;
 wire \systolic_inst.acc_wires[3][26] ;
 wire \systolic_inst.acc_wires[3][27] ;
 wire \systolic_inst.acc_wires[3][28] ;
 wire \systolic_inst.acc_wires[3][29] ;
 wire \systolic_inst.acc_wires[3][2] ;
 wire \systolic_inst.acc_wires[3][30] ;
 wire \systolic_inst.acc_wires[3][31] ;
 wire \systolic_inst.acc_wires[3][3] ;
 wire \systolic_inst.acc_wires[3][4] ;
 wire \systolic_inst.acc_wires[3][5] ;
 wire \systolic_inst.acc_wires[3][6] ;
 wire \systolic_inst.acc_wires[3][7] ;
 wire \systolic_inst.acc_wires[3][8] ;
 wire \systolic_inst.acc_wires[3][9] ;
 wire \systolic_inst.acc_wires[4][0] ;
 wire \systolic_inst.acc_wires[4][10] ;
 wire \systolic_inst.acc_wires[4][11] ;
 wire \systolic_inst.acc_wires[4][12] ;
 wire \systolic_inst.acc_wires[4][13] ;
 wire \systolic_inst.acc_wires[4][14] ;
 wire \systolic_inst.acc_wires[4][15] ;
 wire \systolic_inst.acc_wires[4][16] ;
 wire \systolic_inst.acc_wires[4][17] ;
 wire \systolic_inst.acc_wires[4][18] ;
 wire \systolic_inst.acc_wires[4][19] ;
 wire \systolic_inst.acc_wires[4][1] ;
 wire \systolic_inst.acc_wires[4][20] ;
 wire \systolic_inst.acc_wires[4][21] ;
 wire \systolic_inst.acc_wires[4][22] ;
 wire \systolic_inst.acc_wires[4][23] ;
 wire \systolic_inst.acc_wires[4][24] ;
 wire \systolic_inst.acc_wires[4][25] ;
 wire \systolic_inst.acc_wires[4][26] ;
 wire \systolic_inst.acc_wires[4][27] ;
 wire \systolic_inst.acc_wires[4][28] ;
 wire \systolic_inst.acc_wires[4][29] ;
 wire \systolic_inst.acc_wires[4][2] ;
 wire \systolic_inst.acc_wires[4][30] ;
 wire \systolic_inst.acc_wires[4][31] ;
 wire \systolic_inst.acc_wires[4][3] ;
 wire \systolic_inst.acc_wires[4][4] ;
 wire \systolic_inst.acc_wires[4][5] ;
 wire \systolic_inst.acc_wires[4][6] ;
 wire \systolic_inst.acc_wires[4][7] ;
 wire \systolic_inst.acc_wires[4][8] ;
 wire \systolic_inst.acc_wires[4][9] ;
 wire \systolic_inst.acc_wires[5][0] ;
 wire \systolic_inst.acc_wires[5][10] ;
 wire \systolic_inst.acc_wires[5][11] ;
 wire \systolic_inst.acc_wires[5][12] ;
 wire \systolic_inst.acc_wires[5][13] ;
 wire \systolic_inst.acc_wires[5][14] ;
 wire \systolic_inst.acc_wires[5][15] ;
 wire \systolic_inst.acc_wires[5][16] ;
 wire \systolic_inst.acc_wires[5][17] ;
 wire \systolic_inst.acc_wires[5][18] ;
 wire \systolic_inst.acc_wires[5][19] ;
 wire \systolic_inst.acc_wires[5][1] ;
 wire \systolic_inst.acc_wires[5][20] ;
 wire \systolic_inst.acc_wires[5][21] ;
 wire \systolic_inst.acc_wires[5][22] ;
 wire \systolic_inst.acc_wires[5][23] ;
 wire \systolic_inst.acc_wires[5][24] ;
 wire \systolic_inst.acc_wires[5][25] ;
 wire \systolic_inst.acc_wires[5][26] ;
 wire \systolic_inst.acc_wires[5][27] ;
 wire \systolic_inst.acc_wires[5][28] ;
 wire \systolic_inst.acc_wires[5][29] ;
 wire \systolic_inst.acc_wires[5][2] ;
 wire \systolic_inst.acc_wires[5][30] ;
 wire \systolic_inst.acc_wires[5][31] ;
 wire \systolic_inst.acc_wires[5][3] ;
 wire \systolic_inst.acc_wires[5][4] ;
 wire \systolic_inst.acc_wires[5][5] ;
 wire \systolic_inst.acc_wires[5][6] ;
 wire \systolic_inst.acc_wires[5][7] ;
 wire \systolic_inst.acc_wires[5][8] ;
 wire \systolic_inst.acc_wires[5][9] ;
 wire \systolic_inst.acc_wires[6][0] ;
 wire \systolic_inst.acc_wires[6][10] ;
 wire \systolic_inst.acc_wires[6][11] ;
 wire \systolic_inst.acc_wires[6][12] ;
 wire \systolic_inst.acc_wires[6][13] ;
 wire \systolic_inst.acc_wires[6][14] ;
 wire \systolic_inst.acc_wires[6][15] ;
 wire \systolic_inst.acc_wires[6][16] ;
 wire \systolic_inst.acc_wires[6][17] ;
 wire \systolic_inst.acc_wires[6][18] ;
 wire \systolic_inst.acc_wires[6][19] ;
 wire \systolic_inst.acc_wires[6][1] ;
 wire \systolic_inst.acc_wires[6][20] ;
 wire \systolic_inst.acc_wires[6][21] ;
 wire \systolic_inst.acc_wires[6][22] ;
 wire \systolic_inst.acc_wires[6][23] ;
 wire \systolic_inst.acc_wires[6][24] ;
 wire \systolic_inst.acc_wires[6][25] ;
 wire \systolic_inst.acc_wires[6][26] ;
 wire \systolic_inst.acc_wires[6][27] ;
 wire \systolic_inst.acc_wires[6][28] ;
 wire \systolic_inst.acc_wires[6][29] ;
 wire \systolic_inst.acc_wires[6][2] ;
 wire \systolic_inst.acc_wires[6][30] ;
 wire \systolic_inst.acc_wires[6][31] ;
 wire \systolic_inst.acc_wires[6][3] ;
 wire \systolic_inst.acc_wires[6][4] ;
 wire \systolic_inst.acc_wires[6][5] ;
 wire \systolic_inst.acc_wires[6][6] ;
 wire \systolic_inst.acc_wires[6][7] ;
 wire \systolic_inst.acc_wires[6][8] ;
 wire \systolic_inst.acc_wires[6][9] ;
 wire \systolic_inst.acc_wires[7][0] ;
 wire \systolic_inst.acc_wires[7][10] ;
 wire \systolic_inst.acc_wires[7][11] ;
 wire \systolic_inst.acc_wires[7][12] ;
 wire \systolic_inst.acc_wires[7][13] ;
 wire \systolic_inst.acc_wires[7][14] ;
 wire \systolic_inst.acc_wires[7][15] ;
 wire \systolic_inst.acc_wires[7][16] ;
 wire \systolic_inst.acc_wires[7][17] ;
 wire \systolic_inst.acc_wires[7][18] ;
 wire \systolic_inst.acc_wires[7][19] ;
 wire \systolic_inst.acc_wires[7][1] ;
 wire \systolic_inst.acc_wires[7][20] ;
 wire \systolic_inst.acc_wires[7][21] ;
 wire \systolic_inst.acc_wires[7][22] ;
 wire \systolic_inst.acc_wires[7][23] ;
 wire \systolic_inst.acc_wires[7][24] ;
 wire \systolic_inst.acc_wires[7][25] ;
 wire \systolic_inst.acc_wires[7][26] ;
 wire \systolic_inst.acc_wires[7][27] ;
 wire \systolic_inst.acc_wires[7][28] ;
 wire \systolic_inst.acc_wires[7][29] ;
 wire \systolic_inst.acc_wires[7][2] ;
 wire \systolic_inst.acc_wires[7][30] ;
 wire \systolic_inst.acc_wires[7][31] ;
 wire \systolic_inst.acc_wires[7][3] ;
 wire \systolic_inst.acc_wires[7][4] ;
 wire \systolic_inst.acc_wires[7][5] ;
 wire \systolic_inst.acc_wires[7][6] ;
 wire \systolic_inst.acc_wires[7][7] ;
 wire \systolic_inst.acc_wires[7][8] ;
 wire \systolic_inst.acc_wires[7][9] ;
 wire \systolic_inst.acc_wires[8][0] ;
 wire \systolic_inst.acc_wires[8][10] ;
 wire \systolic_inst.acc_wires[8][11] ;
 wire \systolic_inst.acc_wires[8][12] ;
 wire \systolic_inst.acc_wires[8][13] ;
 wire \systolic_inst.acc_wires[8][14] ;
 wire \systolic_inst.acc_wires[8][15] ;
 wire \systolic_inst.acc_wires[8][16] ;
 wire \systolic_inst.acc_wires[8][17] ;
 wire \systolic_inst.acc_wires[8][18] ;
 wire \systolic_inst.acc_wires[8][19] ;
 wire \systolic_inst.acc_wires[8][1] ;
 wire \systolic_inst.acc_wires[8][20] ;
 wire \systolic_inst.acc_wires[8][21] ;
 wire \systolic_inst.acc_wires[8][22] ;
 wire \systolic_inst.acc_wires[8][23] ;
 wire \systolic_inst.acc_wires[8][24] ;
 wire \systolic_inst.acc_wires[8][25] ;
 wire \systolic_inst.acc_wires[8][26] ;
 wire \systolic_inst.acc_wires[8][27] ;
 wire \systolic_inst.acc_wires[8][28] ;
 wire \systolic_inst.acc_wires[8][29] ;
 wire \systolic_inst.acc_wires[8][2] ;
 wire \systolic_inst.acc_wires[8][30] ;
 wire \systolic_inst.acc_wires[8][31] ;
 wire \systolic_inst.acc_wires[8][3] ;
 wire \systolic_inst.acc_wires[8][4] ;
 wire \systolic_inst.acc_wires[8][5] ;
 wire \systolic_inst.acc_wires[8][6] ;
 wire \systolic_inst.acc_wires[8][7] ;
 wire \systolic_inst.acc_wires[8][8] ;
 wire \systolic_inst.acc_wires[8][9] ;
 wire \systolic_inst.acc_wires[9][0] ;
 wire \systolic_inst.acc_wires[9][10] ;
 wire \systolic_inst.acc_wires[9][11] ;
 wire \systolic_inst.acc_wires[9][12] ;
 wire \systolic_inst.acc_wires[9][13] ;
 wire \systolic_inst.acc_wires[9][14] ;
 wire \systolic_inst.acc_wires[9][15] ;
 wire \systolic_inst.acc_wires[9][16] ;
 wire \systolic_inst.acc_wires[9][17] ;
 wire \systolic_inst.acc_wires[9][18] ;
 wire \systolic_inst.acc_wires[9][19] ;
 wire \systolic_inst.acc_wires[9][1] ;
 wire \systolic_inst.acc_wires[9][20] ;
 wire \systolic_inst.acc_wires[9][21] ;
 wire \systolic_inst.acc_wires[9][22] ;
 wire \systolic_inst.acc_wires[9][23] ;
 wire \systolic_inst.acc_wires[9][24] ;
 wire \systolic_inst.acc_wires[9][25] ;
 wire \systolic_inst.acc_wires[9][26] ;
 wire \systolic_inst.acc_wires[9][27] ;
 wire \systolic_inst.acc_wires[9][28] ;
 wire \systolic_inst.acc_wires[9][29] ;
 wire \systolic_inst.acc_wires[9][2] ;
 wire \systolic_inst.acc_wires[9][30] ;
 wire \systolic_inst.acc_wires[9][31] ;
 wire \systolic_inst.acc_wires[9][3] ;
 wire \systolic_inst.acc_wires[9][4] ;
 wire \systolic_inst.acc_wires[9][5] ;
 wire \systolic_inst.acc_wires[9][6] ;
 wire \systolic_inst.acc_wires[9][7] ;
 wire \systolic_inst.acc_wires[9][8] ;
 wire \systolic_inst.acc_wires[9][9] ;
 wire \systolic_inst.ce_local ;
 wire \systolic_inst.cycle_cnt[0] ;
 wire \systolic_inst.cycle_cnt[10] ;
 wire \systolic_inst.cycle_cnt[11] ;
 wire \systolic_inst.cycle_cnt[12] ;
 wire \systolic_inst.cycle_cnt[13] ;
 wire \systolic_inst.cycle_cnt[14] ;
 wire \systolic_inst.cycle_cnt[15] ;
 wire \systolic_inst.cycle_cnt[16] ;
 wire \systolic_inst.cycle_cnt[17] ;
 wire \systolic_inst.cycle_cnt[18] ;
 wire \systolic_inst.cycle_cnt[19] ;
 wire \systolic_inst.cycle_cnt[1] ;
 wire \systolic_inst.cycle_cnt[20] ;
 wire \systolic_inst.cycle_cnt[21] ;
 wire \systolic_inst.cycle_cnt[22] ;
 wire \systolic_inst.cycle_cnt[23] ;
 wire \systolic_inst.cycle_cnt[24] ;
 wire \systolic_inst.cycle_cnt[25] ;
 wire \systolic_inst.cycle_cnt[26] ;
 wire \systolic_inst.cycle_cnt[27] ;
 wire \systolic_inst.cycle_cnt[28] ;
 wire \systolic_inst.cycle_cnt[29] ;
 wire \systolic_inst.cycle_cnt[2] ;
 wire \systolic_inst.cycle_cnt[30] ;
 wire \systolic_inst.cycle_cnt[31] ;
 wire \systolic_inst.cycle_cnt[3] ;
 wire \systolic_inst.cycle_cnt[4] ;
 wire \systolic_inst.cycle_cnt[5] ;
 wire \systolic_inst.cycle_cnt[6] ;
 wire \systolic_inst.cycle_cnt[7] ;
 wire \systolic_inst.cycle_cnt[8] ;
 wire \systolic_inst.cycle_cnt[9] ;
 wire \systolic_inst.load_acc ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[9] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[0] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[10] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[11] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[12] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[13] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[14] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[1] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[2] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[3] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[4] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[5] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[6] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[7] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[8] ;
 wire \systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[9] ;

 sky130_fd_sc_hd__inv_2 _13101_ (.A(\systolic_inst.cycle_cnt[2] ),
    .Y(_11257_));
 sky130_fd_sc_hd__inv_2 _13102_ (.A(\systolic_inst.ce_local ),
    .Y(_11258_));
 sky130_fd_sc_hd__inv_2 _13103_ (.A(\systolic_inst.B_outs[8][7] ),
    .Y(_11259_));
 sky130_fd_sc_hd__inv_2 _13104_ (.A(\systolic_inst.B_outs[12][7] ),
    .Y(_11260_));
 sky130_fd_sc_hd__inv_2 _13105_ (.A(\systolic_inst.B_outs[7][7] ),
    .Y(_11261_));
 sky130_fd_sc_hd__inv_2 _13106_ (.A(\systolic_inst.B_outs[11][7] ),
    .Y(_11262_));
 sky130_fd_sc_hd__inv_2 _13107_ (.A(\systolic_inst.B_outs[9][7] ),
    .Y(_11263_));
 sky130_fd_sc_hd__inv_2 _13108_ (.A(\systolic_inst.B_outs[14][7] ),
    .Y(_11264_));
 sky130_fd_sc_hd__inv_2 _13109_ (.A(\systolic_inst.B_outs[2][7] ),
    .Y(_11265_));
 sky130_fd_sc_hd__inv_2 _13110_ (.A(\systolic_inst.A_outs[0][2] ),
    .Y(_11266_));
 sky130_fd_sc_hd__inv_2 _13111_ (.A(\systolic_inst.A_outs[0][4] ),
    .Y(_11267_));
 sky130_fd_sc_hd__inv_2 _13112_ (.A(\systolic_inst.A_outs[0][5] ),
    .Y(_11268_));
 sky130_fd_sc_hd__inv_2 _13113_ (.A(\systolic_inst.A_outs[0][6] ),
    .Y(_11269_));
 sky130_fd_sc_hd__inv_2 _13114_ (.A(\systolic_inst.A_outs[0][7] ),
    .Y(_11270_));
 sky130_fd_sc_hd__inv_2 _13115_ (.A(\systolic_inst.B_outs[4][7] ),
    .Y(_11271_));
 sky130_fd_sc_hd__inv_2 _13116_ (.A(\systolic_inst.B_outs[13][7] ),
    .Y(_11272_));
 sky130_fd_sc_hd__inv_2 _13117_ (.A(\systolic_inst.B_outs[15][7] ),
    .Y(_11273_));
 sky130_fd_sc_hd__inv_2 _13118_ (.A(\systolic_inst.B_outs[3][7] ),
    .Y(_11274_));
 sky130_fd_sc_hd__inv_2 _13119_ (.A(\systolic_inst.B_outs[10][7] ),
    .Y(_11275_));
 sky130_fd_sc_hd__inv_2 _13120_ (.A(\systolic_inst.B_outs[5][7] ),
    .Y(_11276_));
 sky130_fd_sc_hd__inv_2 _13121_ (.A(\systolic_inst.B_outs[1][7] ),
    .Y(_11277_));
 sky130_fd_sc_hd__inv_2 _13122_ (.A(\systolic_inst.B_outs[6][7] ),
    .Y(_11278_));
 sky130_fd_sc_hd__nand4_2 _13123_ (.A(B_in_valid),
    .B(A_in_valid),
    .C(start),
    .D(_11258_),
    .Y(_11279_));
 sky130_fd_sc_hd__inv_2 _13124_ (.A(_11279_),
    .Y(_00008_));
 sky130_fd_sc_hd__and4_2 _13125_ (.A(\deser_A.receiving ),
    .B(\deser_A.bit_idx[1] ),
    .C(\deser_A.bit_idx[0] ),
    .D(\deser_A.bit_idx[2] ),
    .X(_11280_));
 sky130_fd_sc_hd__and4_2 _13126_ (.A(\deser_A.bit_idx[3] ),
    .B(\deser_A.bit_idx[5] ),
    .C(\deser_A.bit_idx[4] ),
    .D(_11280_),
    .X(_11281_));
 sky130_fd_sc_hd__inv_2 _13127_ (.A(_11281_),
    .Y(_11282_));
 sky130_fd_sc_hd__and2_2 _13128_ (.A(\deser_A.bit_idx[6] ),
    .B(_11281_),
    .X(_00002_));
 sky130_fd_sc_hd__and4_2 _13129_ (.A(\deser_B.receiving ),
    .B(\deser_B.bit_idx[1] ),
    .C(\deser_B.bit_idx[0] ),
    .D(\deser_B.bit_idx[2] ),
    .X(_11283_));
 sky130_fd_sc_hd__and4_2 _13130_ (.A(\deser_B.bit_idx[3] ),
    .B(\deser_B.bit_idx[5] ),
    .C(\deser_B.bit_idx[4] ),
    .D(_11283_),
    .X(_11284_));
 sky130_fd_sc_hd__inv_2 _13131_ (.A(_11284_),
    .Y(_11285_));
 sky130_fd_sc_hd__and2_2 _13132_ (.A(\deser_B.bit_idx[6] ),
    .B(_11284_),
    .X(_00001_));
 sky130_fd_sc_hd__or4_2 _13133_ (.A(\systolic_inst.cycle_cnt[23] ),
    .B(\systolic_inst.cycle_cnt[22] ),
    .C(\systolic_inst.cycle_cnt[21] ),
    .D(\systolic_inst.cycle_cnt[20] ),
    .X(_11286_));
 sky130_fd_sc_hd__or4_2 _13134_ (.A(\systolic_inst.cycle_cnt[27] ),
    .B(\systolic_inst.cycle_cnt[26] ),
    .C(\systolic_inst.cycle_cnt[25] ),
    .D(\systolic_inst.cycle_cnt[24] ),
    .X(_11287_));
 sky130_fd_sc_hd__or4_2 _13135_ (.A(\systolic_inst.cycle_cnt[19] ),
    .B(\systolic_inst.cycle_cnt[18] ),
    .C(\systolic_inst.cycle_cnt[17] ),
    .D(\systolic_inst.cycle_cnt[16] ),
    .X(_11288_));
 sky130_fd_sc_hd__o21a_2 _13136_ (.A1(\systolic_inst.cycle_cnt[1] ),
    .A2(\systolic_inst.cycle_cnt[2] ),
    .B1(\systolic_inst.cycle_cnt[3] ),
    .X(_11289_));
 sky130_fd_sc_hd__or3_2 _13137_ (.A(_11286_),
    .B(_11287_),
    .C(_11289_),
    .X(_11290_));
 sky130_fd_sc_hd__or4_2 _13138_ (.A(\systolic_inst.cycle_cnt[15] ),
    .B(\systolic_inst.cycle_cnt[14] ),
    .C(\systolic_inst.cycle_cnt[13] ),
    .D(\systolic_inst.cycle_cnt[12] ),
    .X(_11291_));
 sky130_fd_sc_hd__or4_2 _13139_ (.A(\systolic_inst.cycle_cnt[7] ),
    .B(\systolic_inst.cycle_cnt[6] ),
    .C(\systolic_inst.cycle_cnt[5] ),
    .D(\systolic_inst.cycle_cnt[4] ),
    .X(_11292_));
 sky130_fd_sc_hd__or4_2 _13140_ (.A(\systolic_inst.cycle_cnt[30] ),
    .B(\systolic_inst.cycle_cnt[31] ),
    .C(\systolic_inst.cycle_cnt[29] ),
    .D(\systolic_inst.cycle_cnt[28] ),
    .X(_11293_));
 sky130_fd_sc_hd__or4_2 _13141_ (.A(\systolic_inst.cycle_cnt[11] ),
    .B(\systolic_inst.cycle_cnt[10] ),
    .C(\systolic_inst.cycle_cnt[9] ),
    .D(\systolic_inst.cycle_cnt[8] ),
    .X(_11294_));
 sky130_fd_sc_hd__or3_2 _13142_ (.A(_11291_),
    .B(_11292_),
    .C(_11293_),
    .X(_11295_));
 sky130_fd_sc_hd__or2_2 _13143_ (.A(_11294_),
    .B(_11295_),
    .X(_11296_));
 sky130_fd_sc_hd__o31ai_2 _13144_ (.A1(_11288_),
    .A2(_11290_),
    .A3(_11296_),
    .B1(\systolic_inst.ce_local ),
    .Y(_11297_));
 sky130_fd_sc_hd__inv_2 _13145_ (.A(_11297_),
    .Y(_00000_));
 sky130_fd_sc_hd__and4_2 _13146_ (.A(\ser_C.bit_idx[4] ),
    .B(\ser_C.bit_idx[5] ),
    .C(\ser_C.bit_idx[6] ),
    .D(\ser_C.bit_idx[7] ),
    .X(_11298_));
 sky130_fd_sc_hd__and3_2 _13147_ (.A(\ser_C.bit_idx[0] ),
    .B(\ser_C.bit_idx[3] ),
    .C(_11298_),
    .X(_11299_));
 sky130_fd_sc_hd__and3_2 _13148_ (.A(\ser_C.bit_idx[1] ),
    .B(\ser_C.bit_idx[2] ),
    .C(_11299_),
    .X(_11300_));
 sky130_fd_sc_hd__a21bo_2 _13149_ (.A1(\ser_C.bit_idx[8] ),
    .A2(_11300_),
    .B1_N(C_out_frame_sync),
    .X(_11301_));
 sky130_fd_sc_hd__and2b_2 _13150_ (.A_N(C_out_frame_sync),
    .B(done),
    .X(_11302_));
 sky130_fd_sc_hd__nand2b_2 _13151_ (.A_N(C_out_frame_sync),
    .B(done),
    .Y(_11303_));
 sky130_fd_sc_hd__nand2_2 _13152_ (.A(_11301_),
    .B(_11303_),
    .Y(_00007_));
 sky130_fd_sc_hd__nor2_2 _13153_ (.A(A_in_frame_sync),
    .B(\deser_A.receiving ),
    .Y(_11304_));
 sky130_fd_sc_hd__nor2_2 _13154_ (.A(_00002_),
    .B(_11304_),
    .Y(_00004_));
 sky130_fd_sc_hd__xor2_2 _13155_ (.A(\deser_A.serial_toggle_sync2 ),
    .B(\deser_A.serial_toggle_sync1 ),
    .X(_00003_));
 sky130_fd_sc_hd__nor2_2 _13156_ (.A(B_in_frame_sync),
    .B(\deser_B.receiving ),
    .Y(_11305_));
 sky130_fd_sc_hd__nor2_2 _13157_ (.A(_00001_),
    .B(_11305_),
    .Y(_00006_));
 sky130_fd_sc_hd__xor2_2 _13158_ (.A(\deser_B.serial_toggle_sync2 ),
    .B(\deser_B.serial_toggle_sync1 ),
    .X(_00005_));
 sky130_fd_sc_hd__a31o_2 _13159_ (.A1(B_in_valid),
    .A2(A_in_valid),
    .A3(start),
    .B1(\systolic_inst.ce_local ),
    .X(_11306_));
 sky130_fd_sc_hd__inv_2 _13160_ (.A(_11306_),
    .Y(_11307_));
 sky130_fd_sc_hd__nor2_2 _13161_ (.A(_00000_),
    .B(_11307_),
    .Y(_00009_));
 sky130_fd_sc_hd__mux2_1 _13162_ (.A0(\deser_A.word_buffer[0] ),
    .A1(\deser_A.serial_word[0] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _13163_ (.A0(\deser_A.word_buffer[1] ),
    .A1(\deser_A.serial_word[1] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _13164_ (.A0(\deser_A.word_buffer[2] ),
    .A1(\deser_A.serial_word[2] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _13165_ (.A0(\deser_A.word_buffer[3] ),
    .A1(\deser_A.serial_word[3] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _13166_ (.A0(\deser_A.word_buffer[4] ),
    .A1(\deser_A.serial_word[4] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _13167_ (.A0(\deser_A.word_buffer[5] ),
    .A1(\deser_A.serial_word[5] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _13168_ (.A0(\deser_A.word_buffer[6] ),
    .A1(\deser_A.serial_word[6] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _13169_ (.A0(\deser_A.word_buffer[7] ),
    .A1(\deser_A.serial_word[7] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _13170_ (.A0(\deser_A.word_buffer[8] ),
    .A1(\deser_A.serial_word[8] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _13171_ (.A0(\deser_A.word_buffer[9] ),
    .A1(\deser_A.serial_word[9] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _13172_ (.A0(\deser_A.word_buffer[10] ),
    .A1(\deser_A.serial_word[10] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _13173_ (.A0(\deser_A.word_buffer[11] ),
    .A1(\deser_A.serial_word[11] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _13174_ (.A0(\deser_A.word_buffer[12] ),
    .A1(\deser_A.serial_word[12] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _13175_ (.A0(\deser_A.word_buffer[13] ),
    .A1(\deser_A.serial_word[13] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(\deser_A.word_buffer[14] ),
    .A1(\deser_A.serial_word[14] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _13177_ (.A0(\deser_A.word_buffer[15] ),
    .A1(\deser_A.serial_word[15] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _13178_ (.A0(\deser_A.word_buffer[16] ),
    .A1(\deser_A.serial_word[16] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _13179_ (.A0(\deser_A.word_buffer[17] ),
    .A1(\deser_A.serial_word[17] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _13180_ (.A0(\deser_A.word_buffer[18] ),
    .A1(\deser_A.serial_word[18] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _13181_ (.A0(\deser_A.word_buffer[19] ),
    .A1(\deser_A.serial_word[19] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _13182_ (.A0(\deser_A.word_buffer[20] ),
    .A1(\deser_A.serial_word[20] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _13183_ (.A0(\deser_A.word_buffer[21] ),
    .A1(\deser_A.serial_word[21] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _13184_ (.A0(\deser_A.word_buffer[22] ),
    .A1(\deser_A.serial_word[22] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(\deser_A.word_buffer[23] ),
    .A1(\deser_A.serial_word[23] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _13186_ (.A0(\deser_A.word_buffer[24] ),
    .A1(\deser_A.serial_word[24] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _13187_ (.A0(\deser_A.word_buffer[25] ),
    .A1(\deser_A.serial_word[25] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _13188_ (.A0(\deser_A.word_buffer[26] ),
    .A1(\deser_A.serial_word[26] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _13189_ (.A0(\deser_A.word_buffer[27] ),
    .A1(\deser_A.serial_word[27] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(\deser_A.word_buffer[28] ),
    .A1(\deser_A.serial_word[28] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _13191_ (.A0(\deser_A.word_buffer[29] ),
    .A1(\deser_A.serial_word[29] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _13192_ (.A0(\deser_A.word_buffer[30] ),
    .A1(\deser_A.serial_word[30] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _13193_ (.A0(\deser_A.word_buffer[31] ),
    .A1(\deser_A.serial_word[31] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_1 _13194_ (.A0(\deser_A.word_buffer[32] ),
    .A1(\deser_A.serial_word[32] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _13195_ (.A0(\deser_A.word_buffer[33] ),
    .A1(\deser_A.serial_word[33] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _13196_ (.A0(\deser_A.word_buffer[34] ),
    .A1(\deser_A.serial_word[34] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _13197_ (.A0(\deser_A.word_buffer[35] ),
    .A1(\deser_A.serial_word[35] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _13198_ (.A0(\deser_A.word_buffer[36] ),
    .A1(\deser_A.serial_word[36] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _13199_ (.A0(\deser_A.word_buffer[37] ),
    .A1(\deser_A.serial_word[37] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _13200_ (.A0(\deser_A.word_buffer[38] ),
    .A1(\deser_A.serial_word[38] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _13201_ (.A0(\deser_A.word_buffer[39] ),
    .A1(\deser_A.serial_word[39] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _13202_ (.A0(\deser_A.word_buffer[40] ),
    .A1(\deser_A.serial_word[40] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _13203_ (.A0(\deser_A.word_buffer[41] ),
    .A1(\deser_A.serial_word[41] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _13204_ (.A0(\deser_A.word_buffer[42] ),
    .A1(\deser_A.serial_word[42] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _13205_ (.A0(\deser_A.word_buffer[43] ),
    .A1(\deser_A.serial_word[43] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _13206_ (.A0(\deser_A.word_buffer[44] ),
    .A1(\deser_A.serial_word[44] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _13207_ (.A0(\deser_A.word_buffer[45] ),
    .A1(\deser_A.serial_word[45] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _13208_ (.A0(\deser_A.word_buffer[46] ),
    .A1(\deser_A.serial_word[46] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _13209_ (.A0(\deser_A.word_buffer[47] ),
    .A1(\deser_A.serial_word[47] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _13210_ (.A0(\deser_A.word_buffer[48] ),
    .A1(\deser_A.serial_word[48] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _13211_ (.A0(\deser_A.word_buffer[49] ),
    .A1(\deser_A.serial_word[49] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _13212_ (.A0(\deser_A.word_buffer[50] ),
    .A1(\deser_A.serial_word[50] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _13213_ (.A0(\deser_A.word_buffer[51] ),
    .A1(\deser_A.serial_word[51] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _13214_ (.A0(\deser_A.word_buffer[52] ),
    .A1(\deser_A.serial_word[52] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _13215_ (.A0(\deser_A.word_buffer[53] ),
    .A1(\deser_A.serial_word[53] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _13216_ (.A0(\deser_A.word_buffer[54] ),
    .A1(\deser_A.serial_word[54] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(\deser_A.word_buffer[55] ),
    .A1(\deser_A.serial_word[55] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _13218_ (.A0(\deser_A.word_buffer[56] ),
    .A1(\deser_A.serial_word[56] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(\deser_A.word_buffer[57] ),
    .A1(\deser_A.serial_word[57] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _13220_ (.A0(\deser_A.word_buffer[58] ),
    .A1(\deser_A.serial_word[58] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(\deser_A.word_buffer[59] ),
    .A1(\deser_A.serial_word[59] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _13222_ (.A0(\deser_A.word_buffer[60] ),
    .A1(\deser_A.serial_word[60] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _13223_ (.A0(\deser_A.word_buffer[61] ),
    .A1(\deser_A.serial_word[61] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _13224_ (.A0(\deser_A.word_buffer[62] ),
    .A1(\deser_A.serial_word[62] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _13225_ (.A0(\deser_A.word_buffer[63] ),
    .A1(\deser_A.serial_word[63] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _13226_ (.A0(\deser_A.word_buffer[64] ),
    .A1(\deser_A.serial_word[64] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _13227_ (.A0(\deser_A.word_buffer[65] ),
    .A1(\deser_A.serial_word[65] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _13228_ (.A0(\deser_A.word_buffer[66] ),
    .A1(\deser_A.serial_word[66] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _13229_ (.A0(\deser_A.word_buffer[67] ),
    .A1(\deser_A.serial_word[67] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _13230_ (.A0(\deser_A.word_buffer[68] ),
    .A1(\deser_A.serial_word[68] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _13231_ (.A0(\deser_A.word_buffer[69] ),
    .A1(\deser_A.serial_word[69] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _13232_ (.A0(\deser_A.word_buffer[70] ),
    .A1(\deser_A.serial_word[70] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _13233_ (.A0(\deser_A.word_buffer[71] ),
    .A1(\deser_A.serial_word[71] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _13234_ (.A0(\deser_A.word_buffer[72] ),
    .A1(\deser_A.serial_word[72] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _13235_ (.A0(\deser_A.word_buffer[73] ),
    .A1(\deser_A.serial_word[73] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _13236_ (.A0(\deser_A.word_buffer[74] ),
    .A1(\deser_A.serial_word[74] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _13237_ (.A0(\deser_A.word_buffer[75] ),
    .A1(\deser_A.serial_word[75] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _13238_ (.A0(\deser_A.word_buffer[76] ),
    .A1(\deser_A.serial_word[76] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _13239_ (.A0(\deser_A.word_buffer[77] ),
    .A1(\deser_A.serial_word[77] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _13240_ (.A0(\deser_A.word_buffer[78] ),
    .A1(\deser_A.serial_word[78] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _13241_ (.A0(\deser_A.word_buffer[79] ),
    .A1(\deser_A.serial_word[79] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _13242_ (.A0(\deser_A.word_buffer[80] ),
    .A1(\deser_A.serial_word[80] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _13243_ (.A0(\deser_A.word_buffer[81] ),
    .A1(\deser_A.serial_word[81] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _13244_ (.A0(\deser_A.word_buffer[82] ),
    .A1(\deser_A.serial_word[82] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _13245_ (.A0(\deser_A.word_buffer[83] ),
    .A1(\deser_A.serial_word[83] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _13246_ (.A0(\deser_A.word_buffer[84] ),
    .A1(\deser_A.serial_word[84] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _13247_ (.A0(\deser_A.word_buffer[85] ),
    .A1(\deser_A.serial_word[85] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _13248_ (.A0(\deser_A.word_buffer[86] ),
    .A1(\deser_A.serial_word[86] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _13249_ (.A0(\deser_A.word_buffer[87] ),
    .A1(\deser_A.serial_word[87] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _13250_ (.A0(\deser_A.word_buffer[88] ),
    .A1(\deser_A.serial_word[88] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _13251_ (.A0(\deser_A.word_buffer[89] ),
    .A1(\deser_A.serial_word[89] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _13252_ (.A0(\deser_A.word_buffer[90] ),
    .A1(\deser_A.serial_word[90] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _13253_ (.A0(\deser_A.word_buffer[91] ),
    .A1(\deser_A.serial_word[91] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _13254_ (.A0(\deser_A.word_buffer[92] ),
    .A1(\deser_A.serial_word[92] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _13255_ (.A0(\deser_A.word_buffer[93] ),
    .A1(\deser_A.serial_word[93] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _13256_ (.A0(\deser_A.word_buffer[94] ),
    .A1(\deser_A.serial_word[94] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _13257_ (.A0(\deser_A.word_buffer[95] ),
    .A1(\deser_A.serial_word[95] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _13258_ (.A0(\deser_A.word_buffer[96] ),
    .A1(\deser_A.serial_word[96] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _13259_ (.A0(\deser_A.word_buffer[97] ),
    .A1(\deser_A.serial_word[97] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _13260_ (.A0(\deser_A.word_buffer[98] ),
    .A1(\deser_A.serial_word[98] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _13261_ (.A0(\deser_A.word_buffer[99] ),
    .A1(\deser_A.serial_word[99] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _13262_ (.A0(\deser_A.word_buffer[100] ),
    .A1(\deser_A.serial_word[100] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _13263_ (.A0(\deser_A.word_buffer[101] ),
    .A1(\deser_A.serial_word[101] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _13264_ (.A0(\deser_A.word_buffer[102] ),
    .A1(\deser_A.serial_word[102] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _13265_ (.A0(\deser_A.word_buffer[103] ),
    .A1(\deser_A.serial_word[103] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _13266_ (.A0(\deser_A.word_buffer[104] ),
    .A1(\deser_A.serial_word[104] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _13267_ (.A0(\deser_A.word_buffer[105] ),
    .A1(\deser_A.serial_word[105] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _13268_ (.A0(\deser_A.word_buffer[106] ),
    .A1(\deser_A.serial_word[106] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _13269_ (.A0(\deser_A.word_buffer[107] ),
    .A1(\deser_A.serial_word[107] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _13270_ (.A0(\deser_A.word_buffer[108] ),
    .A1(\deser_A.serial_word[108] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _13271_ (.A0(\deser_A.word_buffer[109] ),
    .A1(\deser_A.serial_word[109] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _13272_ (.A0(\deser_A.word_buffer[110] ),
    .A1(\deser_A.serial_word[110] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _13273_ (.A0(\deser_A.word_buffer[111] ),
    .A1(\deser_A.serial_word[111] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _13274_ (.A0(\deser_A.word_buffer[112] ),
    .A1(\deser_A.serial_word[112] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _13275_ (.A0(\deser_A.word_buffer[113] ),
    .A1(\deser_A.serial_word[113] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _13276_ (.A0(\deser_A.word_buffer[114] ),
    .A1(\deser_A.serial_word[114] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _13277_ (.A0(\deser_A.word_buffer[115] ),
    .A1(\deser_A.serial_word[115] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _13278_ (.A0(\deser_A.word_buffer[116] ),
    .A1(\deser_A.serial_word[116] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _13279_ (.A0(\deser_A.word_buffer[117] ),
    .A1(\deser_A.serial_word[117] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _13280_ (.A0(\deser_A.word_buffer[118] ),
    .A1(\deser_A.serial_word[118] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _13281_ (.A0(\deser_A.word_buffer[119] ),
    .A1(\deser_A.serial_word[119] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _13282_ (.A0(\deser_A.word_buffer[120] ),
    .A1(\deser_A.serial_word[120] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _13283_ (.A0(\deser_A.word_buffer[121] ),
    .A1(\deser_A.serial_word[121] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _13284_ (.A0(\deser_A.word_buffer[122] ),
    .A1(\deser_A.serial_word[122] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _13285_ (.A0(\deser_A.word_buffer[123] ),
    .A1(\deser_A.serial_word[123] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _13286_ (.A0(\deser_A.word_buffer[124] ),
    .A1(\deser_A.serial_word[124] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _13287_ (.A0(\deser_A.word_buffer[125] ),
    .A1(\deser_A.serial_word[125] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _13288_ (.A0(\deser_A.word_buffer[126] ),
    .A1(\deser_A.serial_word[126] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _13289_ (.A0(\deser_A.word_buffer[127] ),
    .A1(\deser_A.serial_word[127] ),
    .S(\deser_A.serial_word_ready ),
    .X(_00137_));
 sky130_fd_sc_hd__xor2_2 _13290_ (.A(\deser_A.serial_toggle ),
    .B(\deser_A.serial_word_ready ),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _13291_ (.A0(\A_in[0] ),
    .A1(\deser_A.word_buffer[0] ),
    .S(_00003_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _13292_ (.A0(\A_in[1] ),
    .A1(\deser_A.word_buffer[1] ),
    .S(_00003_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _13293_ (.A0(\A_in[2] ),
    .A1(\deser_A.word_buffer[2] ),
    .S(_00003_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _13294_ (.A0(\A_in[3] ),
    .A1(\deser_A.word_buffer[3] ),
    .S(_00003_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _13295_ (.A0(\A_in[4] ),
    .A1(\deser_A.word_buffer[4] ),
    .S(_00003_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _13296_ (.A0(\A_in[5] ),
    .A1(\deser_A.word_buffer[5] ),
    .S(_00003_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _13297_ (.A0(\A_in[6] ),
    .A1(\deser_A.word_buffer[6] ),
    .S(_00003_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _13298_ (.A0(\A_in[7] ),
    .A1(\deser_A.word_buffer[7] ),
    .S(_00003_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _13299_ (.A0(\A_in[8] ),
    .A1(\deser_A.word_buffer[8] ),
    .S(_00003_),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _13300_ (.A0(\A_in[9] ),
    .A1(\deser_A.word_buffer[9] ),
    .S(_00003_),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _13301_ (.A0(\A_in[10] ),
    .A1(\deser_A.word_buffer[10] ),
    .S(_00003_),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _13302_ (.A0(\A_in[11] ),
    .A1(\deser_A.word_buffer[11] ),
    .S(_00003_),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _13303_ (.A0(\A_in[12] ),
    .A1(\deser_A.word_buffer[12] ),
    .S(_00003_),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _13304_ (.A0(\A_in[13] ),
    .A1(\deser_A.word_buffer[13] ),
    .S(_00003_),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _13305_ (.A0(\A_in[14] ),
    .A1(\deser_A.word_buffer[14] ),
    .S(_00003_),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _13306_ (.A0(\A_in[15] ),
    .A1(\deser_A.word_buffer[15] ),
    .S(_00003_),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _13307_ (.A0(\A_in[16] ),
    .A1(\deser_A.word_buffer[16] ),
    .S(_00003_),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _13308_ (.A0(\A_in[17] ),
    .A1(\deser_A.word_buffer[17] ),
    .S(_00003_),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _13309_ (.A0(\A_in[18] ),
    .A1(\deser_A.word_buffer[18] ),
    .S(_00003_),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _13310_ (.A0(\A_in[19] ),
    .A1(\deser_A.word_buffer[19] ),
    .S(_00003_),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _13311_ (.A0(\A_in[20] ),
    .A1(\deser_A.word_buffer[20] ),
    .S(_00003_),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _13312_ (.A0(\A_in[21] ),
    .A1(\deser_A.word_buffer[21] ),
    .S(_00003_),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _13313_ (.A0(\A_in[22] ),
    .A1(\deser_A.word_buffer[22] ),
    .S(_00003_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _13314_ (.A0(\A_in[23] ),
    .A1(\deser_A.word_buffer[23] ),
    .S(_00003_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _13315_ (.A0(\A_in[24] ),
    .A1(\deser_A.word_buffer[24] ),
    .S(_00003_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _13316_ (.A0(\A_in[25] ),
    .A1(\deser_A.word_buffer[25] ),
    .S(_00003_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _13317_ (.A0(\A_in[26] ),
    .A1(\deser_A.word_buffer[26] ),
    .S(_00003_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _13318_ (.A0(\A_in[27] ),
    .A1(\deser_A.word_buffer[27] ),
    .S(_00003_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _13319_ (.A0(\A_in[28] ),
    .A1(\deser_A.word_buffer[28] ),
    .S(_00003_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _13320_ (.A0(\A_in[29] ),
    .A1(\deser_A.word_buffer[29] ),
    .S(_00003_),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _13321_ (.A0(\A_in[30] ),
    .A1(\deser_A.word_buffer[30] ),
    .S(_00003_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _13322_ (.A0(\A_in[31] ),
    .A1(\deser_A.word_buffer[31] ),
    .S(_00003_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _13323_ (.A0(\A_in[32] ),
    .A1(\deser_A.word_buffer[32] ),
    .S(_00003_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _13324_ (.A0(\A_in[33] ),
    .A1(\deser_A.word_buffer[33] ),
    .S(_00003_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _13325_ (.A0(\A_in[34] ),
    .A1(\deser_A.word_buffer[34] ),
    .S(_00003_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _13326_ (.A0(\A_in[35] ),
    .A1(\deser_A.word_buffer[35] ),
    .S(_00003_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _13327_ (.A0(\A_in[36] ),
    .A1(\deser_A.word_buffer[36] ),
    .S(_00003_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _13328_ (.A0(\A_in[37] ),
    .A1(\deser_A.word_buffer[37] ),
    .S(_00003_),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _13329_ (.A0(\A_in[38] ),
    .A1(\deser_A.word_buffer[38] ),
    .S(_00003_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _13330_ (.A0(\A_in[39] ),
    .A1(\deser_A.word_buffer[39] ),
    .S(_00003_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _13331_ (.A0(\A_in[40] ),
    .A1(\deser_A.word_buffer[40] ),
    .S(_00003_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _13332_ (.A0(\A_in[41] ),
    .A1(\deser_A.word_buffer[41] ),
    .S(_00003_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _13333_ (.A0(\A_in[42] ),
    .A1(\deser_A.word_buffer[42] ),
    .S(_00003_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _13334_ (.A0(\A_in[43] ),
    .A1(\deser_A.word_buffer[43] ),
    .S(_00003_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _13335_ (.A0(\A_in[44] ),
    .A1(\deser_A.word_buffer[44] ),
    .S(_00003_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _13336_ (.A0(\A_in[45] ),
    .A1(\deser_A.word_buffer[45] ),
    .S(_00003_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _13337_ (.A0(\A_in[46] ),
    .A1(\deser_A.word_buffer[46] ),
    .S(_00003_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _13338_ (.A0(\A_in[47] ),
    .A1(\deser_A.word_buffer[47] ),
    .S(_00003_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _13339_ (.A0(\A_in[48] ),
    .A1(\deser_A.word_buffer[48] ),
    .S(_00003_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _13340_ (.A0(\A_in[49] ),
    .A1(\deser_A.word_buffer[49] ),
    .S(_00003_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _13341_ (.A0(\A_in[50] ),
    .A1(\deser_A.word_buffer[50] ),
    .S(_00003_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _13342_ (.A0(\A_in[51] ),
    .A1(\deser_A.word_buffer[51] ),
    .S(_00003_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _13343_ (.A0(\A_in[52] ),
    .A1(\deser_A.word_buffer[52] ),
    .S(_00003_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _13344_ (.A0(\A_in[53] ),
    .A1(\deser_A.word_buffer[53] ),
    .S(_00003_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _13345_ (.A0(\A_in[54] ),
    .A1(\deser_A.word_buffer[54] ),
    .S(_00003_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _13346_ (.A0(\A_in[55] ),
    .A1(\deser_A.word_buffer[55] ),
    .S(_00003_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _13347_ (.A0(\A_in[56] ),
    .A1(\deser_A.word_buffer[56] ),
    .S(_00003_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _13348_ (.A0(\A_in[57] ),
    .A1(\deser_A.word_buffer[57] ),
    .S(_00003_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _13349_ (.A0(\A_in[58] ),
    .A1(\deser_A.word_buffer[58] ),
    .S(_00003_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _13350_ (.A0(\A_in[59] ),
    .A1(\deser_A.word_buffer[59] ),
    .S(_00003_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _13351_ (.A0(\A_in[60] ),
    .A1(\deser_A.word_buffer[60] ),
    .S(_00003_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _13352_ (.A0(\A_in[61] ),
    .A1(\deser_A.word_buffer[61] ),
    .S(_00003_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _13353_ (.A0(\A_in[62] ),
    .A1(\deser_A.word_buffer[62] ),
    .S(_00003_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _13354_ (.A0(\A_in[63] ),
    .A1(\deser_A.word_buffer[63] ),
    .S(_00003_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _13355_ (.A0(\A_in[64] ),
    .A1(\deser_A.word_buffer[64] ),
    .S(_00003_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _13356_ (.A0(\A_in[65] ),
    .A1(\deser_A.word_buffer[65] ),
    .S(_00003_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _13357_ (.A0(\A_in[66] ),
    .A1(\deser_A.word_buffer[66] ),
    .S(_00003_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _13358_ (.A0(\A_in[67] ),
    .A1(\deser_A.word_buffer[67] ),
    .S(_00003_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _13359_ (.A0(\A_in[68] ),
    .A1(\deser_A.word_buffer[68] ),
    .S(_00003_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _13360_ (.A0(\A_in[69] ),
    .A1(\deser_A.word_buffer[69] ),
    .S(_00003_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _13361_ (.A0(\A_in[70] ),
    .A1(\deser_A.word_buffer[70] ),
    .S(_00003_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _13362_ (.A0(\A_in[71] ),
    .A1(\deser_A.word_buffer[71] ),
    .S(_00003_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _13363_ (.A0(\A_in[72] ),
    .A1(\deser_A.word_buffer[72] ),
    .S(_00003_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _13364_ (.A0(\A_in[73] ),
    .A1(\deser_A.word_buffer[73] ),
    .S(_00003_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _13365_ (.A0(\A_in[74] ),
    .A1(\deser_A.word_buffer[74] ),
    .S(_00003_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _13366_ (.A0(\A_in[75] ),
    .A1(\deser_A.word_buffer[75] ),
    .S(_00003_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _13367_ (.A0(\A_in[76] ),
    .A1(\deser_A.word_buffer[76] ),
    .S(_00003_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _13368_ (.A0(\A_in[77] ),
    .A1(\deser_A.word_buffer[77] ),
    .S(_00003_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _13369_ (.A0(\A_in[78] ),
    .A1(\deser_A.word_buffer[78] ),
    .S(_00003_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _13370_ (.A0(\A_in[79] ),
    .A1(\deser_A.word_buffer[79] ),
    .S(_00003_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _13371_ (.A0(\A_in[80] ),
    .A1(\deser_A.word_buffer[80] ),
    .S(_00003_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _13372_ (.A0(\A_in[81] ),
    .A1(\deser_A.word_buffer[81] ),
    .S(_00003_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _13373_ (.A0(\A_in[82] ),
    .A1(\deser_A.word_buffer[82] ),
    .S(_00003_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _13374_ (.A0(\A_in[83] ),
    .A1(\deser_A.word_buffer[83] ),
    .S(_00003_),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _13375_ (.A0(\A_in[84] ),
    .A1(\deser_A.word_buffer[84] ),
    .S(_00003_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _13376_ (.A0(\A_in[85] ),
    .A1(\deser_A.word_buffer[85] ),
    .S(_00003_),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _13377_ (.A0(\A_in[86] ),
    .A1(\deser_A.word_buffer[86] ),
    .S(_00003_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _13378_ (.A0(\A_in[87] ),
    .A1(\deser_A.word_buffer[87] ),
    .S(_00003_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _13379_ (.A0(\A_in[88] ),
    .A1(\deser_A.word_buffer[88] ),
    .S(_00003_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _13380_ (.A0(\A_in[89] ),
    .A1(\deser_A.word_buffer[89] ),
    .S(_00003_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _13381_ (.A0(\A_in[90] ),
    .A1(\deser_A.word_buffer[90] ),
    .S(_00003_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _13382_ (.A0(\A_in[91] ),
    .A1(\deser_A.word_buffer[91] ),
    .S(_00003_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _13383_ (.A0(\A_in[92] ),
    .A1(\deser_A.word_buffer[92] ),
    .S(_00003_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _13384_ (.A0(\A_in[93] ),
    .A1(\deser_A.word_buffer[93] ),
    .S(_00003_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _13385_ (.A0(\A_in[94] ),
    .A1(\deser_A.word_buffer[94] ),
    .S(_00003_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _13386_ (.A0(\A_in[95] ),
    .A1(\deser_A.word_buffer[95] ),
    .S(_00003_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _13387_ (.A0(\A_in[96] ),
    .A1(\deser_A.word_buffer[96] ),
    .S(_00003_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _13388_ (.A0(\A_in[97] ),
    .A1(\deser_A.word_buffer[97] ),
    .S(_00003_),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _13389_ (.A0(\A_in[98] ),
    .A1(\deser_A.word_buffer[98] ),
    .S(_00003_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _13390_ (.A0(\A_in[99] ),
    .A1(\deser_A.word_buffer[99] ),
    .S(_00003_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _13391_ (.A0(\A_in[100] ),
    .A1(\deser_A.word_buffer[100] ),
    .S(_00003_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _13392_ (.A0(\A_in[101] ),
    .A1(\deser_A.word_buffer[101] ),
    .S(_00003_),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _13393_ (.A0(\A_in[102] ),
    .A1(\deser_A.word_buffer[102] ),
    .S(_00003_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _13394_ (.A0(\A_in[103] ),
    .A1(\deser_A.word_buffer[103] ),
    .S(_00003_),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _13395_ (.A0(\A_in[104] ),
    .A1(\deser_A.word_buffer[104] ),
    .S(_00003_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _13396_ (.A0(\A_in[105] ),
    .A1(\deser_A.word_buffer[105] ),
    .S(_00003_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _13397_ (.A0(\A_in[106] ),
    .A1(\deser_A.word_buffer[106] ),
    .S(_00003_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _13398_ (.A0(\A_in[107] ),
    .A1(\deser_A.word_buffer[107] ),
    .S(_00003_),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _13399_ (.A0(\A_in[108] ),
    .A1(\deser_A.word_buffer[108] ),
    .S(_00003_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _13400_ (.A0(\A_in[109] ),
    .A1(\deser_A.word_buffer[109] ),
    .S(_00003_),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _13401_ (.A0(\A_in[110] ),
    .A1(\deser_A.word_buffer[110] ),
    .S(_00003_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _13402_ (.A0(\A_in[111] ),
    .A1(\deser_A.word_buffer[111] ),
    .S(_00003_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _13403_ (.A0(\A_in[112] ),
    .A1(\deser_A.word_buffer[112] ),
    .S(_00003_),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _13404_ (.A0(\A_in[113] ),
    .A1(\deser_A.word_buffer[113] ),
    .S(_00003_),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _13405_ (.A0(\A_in[114] ),
    .A1(\deser_A.word_buffer[114] ),
    .S(_00003_),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _13406_ (.A0(\A_in[115] ),
    .A1(\deser_A.word_buffer[115] ),
    .S(_00003_),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _13407_ (.A0(\A_in[116] ),
    .A1(\deser_A.word_buffer[116] ),
    .S(_00003_),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _13408_ (.A0(\A_in[117] ),
    .A1(\deser_A.word_buffer[117] ),
    .S(_00003_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _13409_ (.A0(\A_in[118] ),
    .A1(\deser_A.word_buffer[118] ),
    .S(_00003_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _13410_ (.A0(\A_in[119] ),
    .A1(\deser_A.word_buffer[119] ),
    .S(_00003_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _13411_ (.A0(\A_in[120] ),
    .A1(\deser_A.word_buffer[120] ),
    .S(_00003_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _13412_ (.A0(\A_in[121] ),
    .A1(\deser_A.word_buffer[121] ),
    .S(_00003_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _13413_ (.A0(\A_in[122] ),
    .A1(\deser_A.word_buffer[122] ),
    .S(_00003_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _13414_ (.A0(\A_in[123] ),
    .A1(\deser_A.word_buffer[123] ),
    .S(_00003_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _13415_ (.A0(\A_in[124] ),
    .A1(\deser_A.word_buffer[124] ),
    .S(_00003_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _13416_ (.A0(\A_in[125] ),
    .A1(\deser_A.word_buffer[125] ),
    .S(_00003_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _13417_ (.A0(\A_in[126] ),
    .A1(\deser_A.word_buffer[126] ),
    .S(_00003_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _13418_ (.A0(\A_in[127] ),
    .A1(\deser_A.word_buffer[127] ),
    .S(_00003_),
    .X(_00266_));
 sky130_fd_sc_hd__o21a_2 _13419_ (.A1(A_in_frame_sync),
    .A2(\deser_A.receiving ),
    .B1(\deser_A.bit_idx[0] ),
    .X(_11308_));
 sky130_fd_sc_hd__o21ba_2 _13420_ (.A1(\deser_A.receiving ),
    .A2(\deser_A.bit_idx[0] ),
    .B1_N(_11308_),
    .X(_00267_));
 sky130_fd_sc_hd__and2_2 _13421_ (.A(\deser_A.bit_idx[1] ),
    .B(_11308_),
    .X(_11309_));
 sky130_fd_sc_hd__nand2b_2 _13422_ (.A_N(\deser_A.receiving ),
    .B(A_in_frame_sync),
    .Y(_11310_));
 sky130_fd_sc_hd__o21ai_2 _13423_ (.A1(\deser_A.bit_idx[1] ),
    .A2(_11308_),
    .B1(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__nor2_2 _13424_ (.A(_11309_),
    .B(_11311_),
    .Y(_00268_));
 sky130_fd_sc_hd__and3_2 _13425_ (.A(\deser_A.bit_idx[1] ),
    .B(\deser_A.bit_idx[2] ),
    .C(_11308_),
    .X(_11312_));
 sky130_fd_sc_hd__o21ai_2 _13426_ (.A1(\deser_A.bit_idx[2] ),
    .A2(_11309_),
    .B1(_11310_),
    .Y(_11313_));
 sky130_fd_sc_hd__nor2_2 _13427_ (.A(_11312_),
    .B(_11313_),
    .Y(_00269_));
 sky130_fd_sc_hd__o21ai_2 _13428_ (.A1(\deser_A.bit_idx[3] ),
    .A2(_11312_),
    .B1(_11310_),
    .Y(_11314_));
 sky130_fd_sc_hd__a21oi_2 _13429_ (.A1(\deser_A.bit_idx[3] ),
    .A2(_11312_),
    .B1(_11314_),
    .Y(_00270_));
 sky130_fd_sc_hd__a31o_2 _13430_ (.A1(\deser_A.bit_idx[3] ),
    .A2(\deser_A.bit_idx[2] ),
    .A3(_11309_),
    .B1(\deser_A.bit_idx[4] ),
    .X(_11315_));
 sky130_fd_sc_hd__and3_2 _13431_ (.A(\deser_A.bit_idx[3] ),
    .B(\deser_A.bit_idx[4] ),
    .C(_11312_),
    .X(_11316_));
 sky130_fd_sc_hd__inv_2 _13432_ (.A(_11316_),
    .Y(_11317_));
 sky130_fd_sc_hd__and3_2 _13433_ (.A(_11310_),
    .B(_11315_),
    .C(_11317_),
    .X(_00271_));
 sky130_fd_sc_hd__o211a_2 _13434_ (.A1(\deser_A.bit_idx[5] ),
    .A2(_11316_),
    .B1(_11310_),
    .C1(_11282_),
    .X(_00272_));
 sky130_fd_sc_hd__a21o_2 _13435_ (.A1(\deser_A.bit_idx[5] ),
    .A2(_11316_),
    .B1(\deser_A.bit_idx[6] ),
    .X(_11318_));
 sky130_fd_sc_hd__and3b_2 _13436_ (.A_N(_00002_),
    .B(_11310_),
    .C(_11318_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _13437_ (.A0(\deser_A.shift_reg[1] ),
    .A1(\deser_A.shift_reg[2] ),
    .S(\deser_A.receiving ),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _13438_ (.A0(\deser_A.shift_reg[2] ),
    .A1(\deser_A.shift_reg[3] ),
    .S(\deser_A.receiving ),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _13439_ (.A0(\deser_A.shift_reg[3] ),
    .A1(\deser_A.shift_reg[4] ),
    .S(\deser_A.receiving ),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _13440_ (.A0(\deser_A.shift_reg[4] ),
    .A1(\deser_A.shift_reg[5] ),
    .S(\deser_A.receiving ),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _13441_ (.A0(\deser_A.shift_reg[5] ),
    .A1(\deser_A.shift_reg[6] ),
    .S(\deser_A.receiving ),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _13442_ (.A0(\deser_A.shift_reg[6] ),
    .A1(\deser_A.shift_reg[7] ),
    .S(\deser_A.receiving ),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _13443_ (.A0(\deser_A.shift_reg[7] ),
    .A1(\deser_A.shift_reg[8] ),
    .S(\deser_A.receiving ),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _13444_ (.A0(\deser_A.shift_reg[8] ),
    .A1(\deser_A.shift_reg[9] ),
    .S(\deser_A.receiving ),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _13445_ (.A0(\deser_A.shift_reg[9] ),
    .A1(\deser_A.shift_reg[10] ),
    .S(\deser_A.receiving ),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _13446_ (.A0(\deser_A.shift_reg[10] ),
    .A1(\deser_A.shift_reg[11] ),
    .S(\deser_A.receiving ),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _13447_ (.A0(\deser_A.shift_reg[11] ),
    .A1(\deser_A.shift_reg[12] ),
    .S(\deser_A.receiving ),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _13448_ (.A0(\deser_A.shift_reg[12] ),
    .A1(\deser_A.shift_reg[13] ),
    .S(\deser_A.receiving ),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _13449_ (.A0(\deser_A.shift_reg[13] ),
    .A1(\deser_A.shift_reg[14] ),
    .S(\deser_A.receiving ),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _13450_ (.A0(\deser_A.shift_reg[14] ),
    .A1(\deser_A.shift_reg[15] ),
    .S(\deser_A.receiving ),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _13451_ (.A0(\deser_A.shift_reg[15] ),
    .A1(\deser_A.shift_reg[16] ),
    .S(\deser_A.receiving ),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _13452_ (.A0(\deser_A.shift_reg[16] ),
    .A1(\deser_A.shift_reg[17] ),
    .S(\deser_A.receiving ),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _13453_ (.A0(\deser_A.shift_reg[17] ),
    .A1(\deser_A.shift_reg[18] ),
    .S(\deser_A.receiving ),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _13454_ (.A0(\deser_A.shift_reg[18] ),
    .A1(\deser_A.shift_reg[19] ),
    .S(\deser_A.receiving ),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _13455_ (.A0(\deser_A.shift_reg[19] ),
    .A1(\deser_A.shift_reg[20] ),
    .S(\deser_A.receiving ),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _13456_ (.A0(\deser_A.shift_reg[20] ),
    .A1(\deser_A.shift_reg[21] ),
    .S(\deser_A.receiving ),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _13457_ (.A0(\deser_A.shift_reg[21] ),
    .A1(\deser_A.shift_reg[22] ),
    .S(\deser_A.receiving ),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _13458_ (.A0(\deser_A.shift_reg[22] ),
    .A1(\deser_A.shift_reg[23] ),
    .S(\deser_A.receiving ),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _13459_ (.A0(\deser_A.shift_reg[23] ),
    .A1(\deser_A.shift_reg[24] ),
    .S(\deser_A.receiving ),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _13460_ (.A0(\deser_A.shift_reg[24] ),
    .A1(\deser_A.shift_reg[25] ),
    .S(\deser_A.receiving ),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _13461_ (.A0(\deser_A.shift_reg[25] ),
    .A1(\deser_A.shift_reg[26] ),
    .S(\deser_A.receiving ),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _13462_ (.A0(\deser_A.shift_reg[26] ),
    .A1(\deser_A.shift_reg[27] ),
    .S(\deser_A.receiving ),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _13463_ (.A0(\deser_A.shift_reg[27] ),
    .A1(\deser_A.shift_reg[28] ),
    .S(\deser_A.receiving ),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _13464_ (.A0(\deser_A.shift_reg[28] ),
    .A1(\deser_A.shift_reg[29] ),
    .S(\deser_A.receiving ),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _13465_ (.A0(\deser_A.shift_reg[29] ),
    .A1(\deser_A.shift_reg[30] ),
    .S(\deser_A.receiving ),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _13466_ (.A0(\deser_A.shift_reg[30] ),
    .A1(\deser_A.shift_reg[31] ),
    .S(\deser_A.receiving ),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _13467_ (.A0(\deser_A.shift_reg[31] ),
    .A1(\deser_A.shift_reg[32] ),
    .S(\deser_A.receiving ),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _13468_ (.A0(\deser_A.shift_reg[32] ),
    .A1(\deser_A.shift_reg[33] ),
    .S(\deser_A.receiving ),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _13469_ (.A0(\deser_A.shift_reg[33] ),
    .A1(\deser_A.shift_reg[34] ),
    .S(\deser_A.receiving ),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _13470_ (.A0(\deser_A.shift_reg[34] ),
    .A1(\deser_A.shift_reg[35] ),
    .S(\deser_A.receiving ),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _13471_ (.A0(\deser_A.shift_reg[35] ),
    .A1(\deser_A.shift_reg[36] ),
    .S(\deser_A.receiving ),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _13472_ (.A0(\deser_A.shift_reg[36] ),
    .A1(\deser_A.shift_reg[37] ),
    .S(\deser_A.receiving ),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _13473_ (.A0(\deser_A.shift_reg[37] ),
    .A1(\deser_A.shift_reg[38] ),
    .S(\deser_A.receiving ),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _13474_ (.A0(\deser_A.shift_reg[38] ),
    .A1(\deser_A.shift_reg[39] ),
    .S(\deser_A.receiving ),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(\deser_A.shift_reg[39] ),
    .A1(\deser_A.shift_reg[40] ),
    .S(\deser_A.receiving ),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _13476_ (.A0(\deser_A.shift_reg[40] ),
    .A1(\deser_A.shift_reg[41] ),
    .S(\deser_A.receiving ),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _13477_ (.A0(\deser_A.shift_reg[41] ),
    .A1(\deser_A.shift_reg[42] ),
    .S(\deser_A.receiving ),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _13478_ (.A0(\deser_A.shift_reg[42] ),
    .A1(\deser_A.shift_reg[43] ),
    .S(\deser_A.receiving ),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _13479_ (.A0(\deser_A.shift_reg[43] ),
    .A1(\deser_A.shift_reg[44] ),
    .S(\deser_A.receiving ),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _13480_ (.A0(\deser_A.shift_reg[44] ),
    .A1(\deser_A.shift_reg[45] ),
    .S(\deser_A.receiving ),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _13481_ (.A0(\deser_A.shift_reg[45] ),
    .A1(\deser_A.shift_reg[46] ),
    .S(\deser_A.receiving ),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _13482_ (.A0(\deser_A.shift_reg[46] ),
    .A1(\deser_A.shift_reg[47] ),
    .S(\deser_A.receiving ),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _13483_ (.A0(\deser_A.shift_reg[47] ),
    .A1(\deser_A.shift_reg[48] ),
    .S(\deser_A.receiving ),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _13484_ (.A0(\deser_A.shift_reg[48] ),
    .A1(\deser_A.shift_reg[49] ),
    .S(\deser_A.receiving ),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _13485_ (.A0(\deser_A.shift_reg[49] ),
    .A1(\deser_A.shift_reg[50] ),
    .S(\deser_A.receiving ),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _13486_ (.A0(\deser_A.shift_reg[50] ),
    .A1(\deser_A.shift_reg[51] ),
    .S(\deser_A.receiving ),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _13487_ (.A0(\deser_A.shift_reg[51] ),
    .A1(\deser_A.shift_reg[52] ),
    .S(\deser_A.receiving ),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _13488_ (.A0(\deser_A.shift_reg[52] ),
    .A1(\deser_A.shift_reg[53] ),
    .S(\deser_A.receiving ),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _13489_ (.A0(\deser_A.shift_reg[53] ),
    .A1(\deser_A.shift_reg[54] ),
    .S(\deser_A.receiving ),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _13490_ (.A0(\deser_A.shift_reg[54] ),
    .A1(\deser_A.shift_reg[55] ),
    .S(\deser_A.receiving ),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _13491_ (.A0(\deser_A.shift_reg[55] ),
    .A1(\deser_A.shift_reg[56] ),
    .S(\deser_A.receiving ),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _13492_ (.A0(\deser_A.shift_reg[56] ),
    .A1(\deser_A.shift_reg[57] ),
    .S(\deser_A.receiving ),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _13493_ (.A0(\deser_A.shift_reg[57] ),
    .A1(\deser_A.shift_reg[58] ),
    .S(\deser_A.receiving ),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _13494_ (.A0(\deser_A.shift_reg[58] ),
    .A1(\deser_A.shift_reg[59] ),
    .S(\deser_A.receiving ),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _13495_ (.A0(\deser_A.shift_reg[59] ),
    .A1(\deser_A.shift_reg[60] ),
    .S(\deser_A.receiving ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _13496_ (.A0(\deser_A.shift_reg[60] ),
    .A1(\deser_A.shift_reg[61] ),
    .S(\deser_A.receiving ),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _13497_ (.A0(\deser_A.shift_reg[61] ),
    .A1(\deser_A.shift_reg[62] ),
    .S(\deser_A.receiving ),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _13498_ (.A0(\deser_A.shift_reg[62] ),
    .A1(\deser_A.shift_reg[63] ),
    .S(\deser_A.receiving ),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _13499_ (.A0(\deser_A.shift_reg[63] ),
    .A1(\deser_A.shift_reg[64] ),
    .S(\deser_A.receiving ),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _13500_ (.A0(\deser_A.shift_reg[64] ),
    .A1(\deser_A.shift_reg[65] ),
    .S(\deser_A.receiving ),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _13501_ (.A0(\deser_A.shift_reg[65] ),
    .A1(\deser_A.shift_reg[66] ),
    .S(\deser_A.receiving ),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _13502_ (.A0(\deser_A.shift_reg[66] ),
    .A1(\deser_A.shift_reg[67] ),
    .S(\deser_A.receiving ),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _13503_ (.A0(\deser_A.shift_reg[67] ),
    .A1(\deser_A.shift_reg[68] ),
    .S(\deser_A.receiving ),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _13504_ (.A0(\deser_A.shift_reg[68] ),
    .A1(\deser_A.shift_reg[69] ),
    .S(\deser_A.receiving ),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _13505_ (.A0(\deser_A.shift_reg[69] ),
    .A1(\deser_A.shift_reg[70] ),
    .S(\deser_A.receiving ),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _13506_ (.A0(\deser_A.shift_reg[70] ),
    .A1(\deser_A.shift_reg[71] ),
    .S(\deser_A.receiving ),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _13507_ (.A0(\deser_A.shift_reg[71] ),
    .A1(\deser_A.shift_reg[72] ),
    .S(\deser_A.receiving ),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _13508_ (.A0(\deser_A.shift_reg[72] ),
    .A1(\deser_A.shift_reg[73] ),
    .S(\deser_A.receiving ),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _13509_ (.A0(\deser_A.shift_reg[73] ),
    .A1(\deser_A.shift_reg[74] ),
    .S(\deser_A.receiving ),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _13510_ (.A0(\deser_A.shift_reg[74] ),
    .A1(\deser_A.shift_reg[75] ),
    .S(\deser_A.receiving ),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _13511_ (.A0(\deser_A.shift_reg[75] ),
    .A1(\deser_A.shift_reg[76] ),
    .S(\deser_A.receiving ),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _13512_ (.A0(\deser_A.shift_reg[76] ),
    .A1(\deser_A.shift_reg[77] ),
    .S(\deser_A.receiving ),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _13513_ (.A0(\deser_A.shift_reg[77] ),
    .A1(\deser_A.shift_reg[78] ),
    .S(\deser_A.receiving ),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _13514_ (.A0(\deser_A.shift_reg[78] ),
    .A1(\deser_A.shift_reg[79] ),
    .S(\deser_A.receiving ),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _13515_ (.A0(\deser_A.shift_reg[79] ),
    .A1(\deser_A.shift_reg[80] ),
    .S(\deser_A.receiving ),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _13516_ (.A0(\deser_A.shift_reg[80] ),
    .A1(\deser_A.shift_reg[81] ),
    .S(\deser_A.receiving ),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _13517_ (.A0(\deser_A.shift_reg[81] ),
    .A1(\deser_A.shift_reg[82] ),
    .S(\deser_A.receiving ),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _13518_ (.A0(\deser_A.shift_reg[82] ),
    .A1(\deser_A.shift_reg[83] ),
    .S(\deser_A.receiving ),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _13519_ (.A0(\deser_A.shift_reg[83] ),
    .A1(\deser_A.shift_reg[84] ),
    .S(\deser_A.receiving ),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _13520_ (.A0(\deser_A.shift_reg[84] ),
    .A1(\deser_A.shift_reg[85] ),
    .S(\deser_A.receiving ),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _13521_ (.A0(\deser_A.shift_reg[85] ),
    .A1(\deser_A.shift_reg[86] ),
    .S(\deser_A.receiving ),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _13522_ (.A0(\deser_A.shift_reg[86] ),
    .A1(\deser_A.shift_reg[87] ),
    .S(\deser_A.receiving ),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _13523_ (.A0(\deser_A.shift_reg[87] ),
    .A1(\deser_A.shift_reg[88] ),
    .S(\deser_A.receiving ),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(\deser_A.shift_reg[88] ),
    .A1(\deser_A.shift_reg[89] ),
    .S(\deser_A.receiving ),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _13525_ (.A0(\deser_A.shift_reg[89] ),
    .A1(\deser_A.shift_reg[90] ),
    .S(\deser_A.receiving ),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _13526_ (.A0(\deser_A.shift_reg[90] ),
    .A1(\deser_A.shift_reg[91] ),
    .S(\deser_A.receiving ),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _13527_ (.A0(\deser_A.shift_reg[91] ),
    .A1(\deser_A.shift_reg[92] ),
    .S(\deser_A.receiving ),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(\deser_A.shift_reg[92] ),
    .A1(\deser_A.shift_reg[93] ),
    .S(\deser_A.receiving ),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _13529_ (.A0(\deser_A.shift_reg[93] ),
    .A1(\deser_A.shift_reg[94] ),
    .S(\deser_A.receiving ),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _13530_ (.A0(\deser_A.shift_reg[94] ),
    .A1(\deser_A.shift_reg[95] ),
    .S(\deser_A.receiving ),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _13531_ (.A0(\deser_A.shift_reg[95] ),
    .A1(\deser_A.shift_reg[96] ),
    .S(\deser_A.receiving ),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(\deser_A.shift_reg[96] ),
    .A1(\deser_A.shift_reg[97] ),
    .S(\deser_A.receiving ),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _13533_ (.A0(\deser_A.shift_reg[97] ),
    .A1(\deser_A.shift_reg[98] ),
    .S(\deser_A.receiving ),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _13534_ (.A0(\deser_A.shift_reg[98] ),
    .A1(\deser_A.shift_reg[99] ),
    .S(\deser_A.receiving ),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _13535_ (.A0(\deser_A.shift_reg[99] ),
    .A1(\deser_A.shift_reg[100] ),
    .S(\deser_A.receiving ),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _13536_ (.A0(\deser_A.shift_reg[100] ),
    .A1(\deser_A.shift_reg[101] ),
    .S(\deser_A.receiving ),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _13537_ (.A0(\deser_A.shift_reg[101] ),
    .A1(\deser_A.shift_reg[102] ),
    .S(\deser_A.receiving ),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _13538_ (.A0(\deser_A.shift_reg[102] ),
    .A1(\deser_A.shift_reg[103] ),
    .S(\deser_A.receiving ),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _13539_ (.A0(\deser_A.shift_reg[103] ),
    .A1(\deser_A.shift_reg[104] ),
    .S(\deser_A.receiving ),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _13540_ (.A0(\deser_A.shift_reg[104] ),
    .A1(\deser_A.shift_reg[105] ),
    .S(\deser_A.receiving ),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _13541_ (.A0(\deser_A.shift_reg[105] ),
    .A1(\deser_A.shift_reg[106] ),
    .S(\deser_A.receiving ),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _13542_ (.A0(\deser_A.shift_reg[106] ),
    .A1(\deser_A.shift_reg[107] ),
    .S(\deser_A.receiving ),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _13543_ (.A0(\deser_A.shift_reg[107] ),
    .A1(\deser_A.shift_reg[108] ),
    .S(\deser_A.receiving ),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _13544_ (.A0(\deser_A.shift_reg[108] ),
    .A1(\deser_A.shift_reg[109] ),
    .S(\deser_A.receiving ),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _13545_ (.A0(\deser_A.shift_reg[109] ),
    .A1(\deser_A.shift_reg[110] ),
    .S(\deser_A.receiving ),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _13546_ (.A0(\deser_A.shift_reg[110] ),
    .A1(\deser_A.shift_reg[111] ),
    .S(\deser_A.receiving ),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _13547_ (.A0(\deser_A.shift_reg[111] ),
    .A1(\deser_A.shift_reg[112] ),
    .S(\deser_A.receiving ),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _13548_ (.A0(\deser_A.shift_reg[112] ),
    .A1(\deser_A.shift_reg[113] ),
    .S(\deser_A.receiving ),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _13549_ (.A0(\deser_A.shift_reg[113] ),
    .A1(\deser_A.shift_reg[114] ),
    .S(\deser_A.receiving ),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _13550_ (.A0(\deser_A.shift_reg[114] ),
    .A1(\deser_A.shift_reg[115] ),
    .S(\deser_A.receiving ),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _13551_ (.A0(\deser_A.shift_reg[115] ),
    .A1(\deser_A.shift_reg[116] ),
    .S(\deser_A.receiving ),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _13552_ (.A0(\deser_A.shift_reg[116] ),
    .A1(\deser_A.shift_reg[117] ),
    .S(\deser_A.receiving ),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _13553_ (.A0(\deser_A.shift_reg[117] ),
    .A1(\deser_A.shift_reg[118] ),
    .S(\deser_A.receiving ),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _13554_ (.A0(\deser_A.shift_reg[118] ),
    .A1(\deser_A.shift_reg[119] ),
    .S(\deser_A.receiving ),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _13555_ (.A0(\deser_A.shift_reg[119] ),
    .A1(\deser_A.shift_reg[120] ),
    .S(\deser_A.receiving ),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _13556_ (.A0(\deser_A.shift_reg[120] ),
    .A1(\deser_A.shift_reg[121] ),
    .S(\deser_A.receiving ),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _13557_ (.A0(\deser_A.shift_reg[121] ),
    .A1(\deser_A.shift_reg[122] ),
    .S(\deser_A.receiving ),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(\deser_A.shift_reg[122] ),
    .A1(\deser_A.shift_reg[123] ),
    .S(\deser_A.receiving ),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _13559_ (.A0(\deser_A.shift_reg[123] ),
    .A1(\deser_A.shift_reg[124] ),
    .S(\deser_A.receiving ),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _13560_ (.A0(\deser_A.shift_reg[124] ),
    .A1(\deser_A.shift_reg[125] ),
    .S(\deser_A.receiving ),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _13561_ (.A0(\deser_A.shift_reg[125] ),
    .A1(\deser_A.shift_reg[126] ),
    .S(\deser_A.receiving ),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _13562_ (.A0(\deser_A.shift_reg[126] ),
    .A1(\deser_A.shift_reg[127] ),
    .S(\deser_A.receiving ),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _13563_ (.A0(\deser_A.shift_reg[127] ),
    .A1(A_in_serial_data),
    .S(\deser_A.receiving ),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _13564_ (.A0(\deser_B.word_buffer[0] ),
    .A1(\deser_B.serial_word[0] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _13565_ (.A0(\deser_B.word_buffer[1] ),
    .A1(\deser_B.serial_word[1] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _13566_ (.A0(\deser_B.word_buffer[2] ),
    .A1(\deser_B.serial_word[2] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _13567_ (.A0(\deser_B.word_buffer[3] ),
    .A1(\deser_B.serial_word[3] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _13568_ (.A0(\deser_B.word_buffer[4] ),
    .A1(\deser_B.serial_word[4] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _13569_ (.A0(\deser_B.word_buffer[5] ),
    .A1(\deser_B.serial_word[5] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _13570_ (.A0(\deser_B.word_buffer[6] ),
    .A1(\deser_B.serial_word[6] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _13571_ (.A0(\deser_B.word_buffer[7] ),
    .A1(\deser_B.serial_word[7] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _13572_ (.A0(\deser_B.word_buffer[8] ),
    .A1(\deser_B.serial_word[8] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _13573_ (.A0(\deser_B.word_buffer[9] ),
    .A1(\deser_B.serial_word[9] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _13574_ (.A0(\deser_B.word_buffer[10] ),
    .A1(\deser_B.serial_word[10] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _13575_ (.A0(\deser_B.word_buffer[11] ),
    .A1(\deser_B.serial_word[11] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _13576_ (.A0(\deser_B.word_buffer[12] ),
    .A1(\deser_B.serial_word[12] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _13577_ (.A0(\deser_B.word_buffer[13] ),
    .A1(\deser_B.serial_word[13] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _13578_ (.A0(\deser_B.word_buffer[14] ),
    .A1(\deser_B.serial_word[14] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _13579_ (.A0(\deser_B.word_buffer[15] ),
    .A1(\deser_B.serial_word[15] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _13580_ (.A0(\deser_B.word_buffer[16] ),
    .A1(\deser_B.serial_word[16] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _13581_ (.A0(\deser_B.word_buffer[17] ),
    .A1(\deser_B.serial_word[17] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _13582_ (.A0(\deser_B.word_buffer[18] ),
    .A1(\deser_B.serial_word[18] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _13583_ (.A0(\deser_B.word_buffer[19] ),
    .A1(\deser_B.serial_word[19] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _13584_ (.A0(\deser_B.word_buffer[20] ),
    .A1(\deser_B.serial_word[20] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _13585_ (.A0(\deser_B.word_buffer[21] ),
    .A1(\deser_B.serial_word[21] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _13586_ (.A0(\deser_B.word_buffer[22] ),
    .A1(\deser_B.serial_word[22] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _13587_ (.A0(\deser_B.word_buffer[23] ),
    .A1(\deser_B.serial_word[23] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _13588_ (.A0(\deser_B.word_buffer[24] ),
    .A1(\deser_B.serial_word[24] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _13589_ (.A0(\deser_B.word_buffer[25] ),
    .A1(\deser_B.serial_word[25] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _13590_ (.A0(\deser_B.word_buffer[26] ),
    .A1(\deser_B.serial_word[26] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _13591_ (.A0(\deser_B.word_buffer[27] ),
    .A1(\deser_B.serial_word[27] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _13592_ (.A0(\deser_B.word_buffer[28] ),
    .A1(\deser_B.serial_word[28] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _13593_ (.A0(\deser_B.word_buffer[29] ),
    .A1(\deser_B.serial_word[29] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _13594_ (.A0(\deser_B.word_buffer[30] ),
    .A1(\deser_B.serial_word[30] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _13595_ (.A0(\deser_B.word_buffer[31] ),
    .A1(\deser_B.serial_word[31] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _13596_ (.A0(\deser_B.word_buffer[32] ),
    .A1(\deser_B.serial_word[32] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _13597_ (.A0(\deser_B.word_buffer[33] ),
    .A1(\deser_B.serial_word[33] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _13598_ (.A0(\deser_B.word_buffer[34] ),
    .A1(\deser_B.serial_word[34] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _13599_ (.A0(\deser_B.word_buffer[35] ),
    .A1(\deser_B.serial_word[35] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _13600_ (.A0(\deser_B.word_buffer[36] ),
    .A1(\deser_B.serial_word[36] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _13601_ (.A0(\deser_B.word_buffer[37] ),
    .A1(\deser_B.serial_word[37] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _13602_ (.A0(\deser_B.word_buffer[38] ),
    .A1(\deser_B.serial_word[38] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _13603_ (.A0(\deser_B.word_buffer[39] ),
    .A1(\deser_B.serial_word[39] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _13604_ (.A0(\deser_B.word_buffer[40] ),
    .A1(\deser_B.serial_word[40] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _13605_ (.A0(\deser_B.word_buffer[41] ),
    .A1(\deser_B.serial_word[41] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _13606_ (.A0(\deser_B.word_buffer[42] ),
    .A1(\deser_B.serial_word[42] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _13607_ (.A0(\deser_B.word_buffer[43] ),
    .A1(\deser_B.serial_word[43] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _13608_ (.A0(\deser_B.word_buffer[44] ),
    .A1(\deser_B.serial_word[44] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _13609_ (.A0(\deser_B.word_buffer[45] ),
    .A1(\deser_B.serial_word[45] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _13610_ (.A0(\deser_B.word_buffer[46] ),
    .A1(\deser_B.serial_word[46] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _13611_ (.A0(\deser_B.word_buffer[47] ),
    .A1(\deser_B.serial_word[47] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _13612_ (.A0(\deser_B.word_buffer[48] ),
    .A1(\deser_B.serial_word[48] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _13613_ (.A0(\deser_B.word_buffer[49] ),
    .A1(\deser_B.serial_word[49] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _13614_ (.A0(\deser_B.word_buffer[50] ),
    .A1(\deser_B.serial_word[50] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _13615_ (.A0(\deser_B.word_buffer[51] ),
    .A1(\deser_B.serial_word[51] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _13616_ (.A0(\deser_B.word_buffer[52] ),
    .A1(\deser_B.serial_word[52] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _13617_ (.A0(\deser_B.word_buffer[53] ),
    .A1(\deser_B.serial_word[53] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _13618_ (.A0(\deser_B.word_buffer[54] ),
    .A1(\deser_B.serial_word[54] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _13619_ (.A0(\deser_B.word_buffer[55] ),
    .A1(\deser_B.serial_word[55] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _13620_ (.A0(\deser_B.word_buffer[56] ),
    .A1(\deser_B.serial_word[56] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _13621_ (.A0(\deser_B.word_buffer[57] ),
    .A1(\deser_B.serial_word[57] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _13622_ (.A0(\deser_B.word_buffer[58] ),
    .A1(\deser_B.serial_word[58] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _13623_ (.A0(\deser_B.word_buffer[59] ),
    .A1(\deser_B.serial_word[59] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _13624_ (.A0(\deser_B.word_buffer[60] ),
    .A1(\deser_B.serial_word[60] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _13625_ (.A0(\deser_B.word_buffer[61] ),
    .A1(\deser_B.serial_word[61] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _13626_ (.A0(\deser_B.word_buffer[62] ),
    .A1(\deser_B.serial_word[62] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _13627_ (.A0(\deser_B.word_buffer[63] ),
    .A1(\deser_B.serial_word[63] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _13628_ (.A0(\deser_B.word_buffer[64] ),
    .A1(\deser_B.serial_word[64] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _13629_ (.A0(\deser_B.word_buffer[65] ),
    .A1(\deser_B.serial_word[65] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _13630_ (.A0(\deser_B.word_buffer[66] ),
    .A1(\deser_B.serial_word[66] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _13631_ (.A0(\deser_B.word_buffer[67] ),
    .A1(\deser_B.serial_word[67] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _13632_ (.A0(\deser_B.word_buffer[68] ),
    .A1(\deser_B.serial_word[68] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _13633_ (.A0(\deser_B.word_buffer[69] ),
    .A1(\deser_B.serial_word[69] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _13634_ (.A0(\deser_B.word_buffer[70] ),
    .A1(\deser_B.serial_word[70] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _13635_ (.A0(\deser_B.word_buffer[71] ),
    .A1(\deser_B.serial_word[71] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _13636_ (.A0(\deser_B.word_buffer[72] ),
    .A1(\deser_B.serial_word[72] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _13637_ (.A0(\deser_B.word_buffer[73] ),
    .A1(\deser_B.serial_word[73] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _13638_ (.A0(\deser_B.word_buffer[74] ),
    .A1(\deser_B.serial_word[74] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _13639_ (.A0(\deser_B.word_buffer[75] ),
    .A1(\deser_B.serial_word[75] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _13640_ (.A0(\deser_B.word_buffer[76] ),
    .A1(\deser_B.serial_word[76] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _13641_ (.A0(\deser_B.word_buffer[77] ),
    .A1(\deser_B.serial_word[77] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _13642_ (.A0(\deser_B.word_buffer[78] ),
    .A1(\deser_B.serial_word[78] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _13643_ (.A0(\deser_B.word_buffer[79] ),
    .A1(\deser_B.serial_word[79] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _13644_ (.A0(\deser_B.word_buffer[80] ),
    .A1(\deser_B.serial_word[80] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _13645_ (.A0(\deser_B.word_buffer[81] ),
    .A1(\deser_B.serial_word[81] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _13646_ (.A0(\deser_B.word_buffer[82] ),
    .A1(\deser_B.serial_word[82] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _13647_ (.A0(\deser_B.word_buffer[83] ),
    .A1(\deser_B.serial_word[83] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _13648_ (.A0(\deser_B.word_buffer[84] ),
    .A1(\deser_B.serial_word[84] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _13649_ (.A0(\deser_B.word_buffer[85] ),
    .A1(\deser_B.serial_word[85] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _13650_ (.A0(\deser_B.word_buffer[86] ),
    .A1(\deser_B.serial_word[86] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _13651_ (.A0(\deser_B.word_buffer[87] ),
    .A1(\deser_B.serial_word[87] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _13652_ (.A0(\deser_B.word_buffer[88] ),
    .A1(\deser_B.serial_word[88] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _13653_ (.A0(\deser_B.word_buffer[89] ),
    .A1(\deser_B.serial_word[89] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _13654_ (.A0(\deser_B.word_buffer[90] ),
    .A1(\deser_B.serial_word[90] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _13655_ (.A0(\deser_B.word_buffer[91] ),
    .A1(\deser_B.serial_word[91] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _13656_ (.A0(\deser_B.word_buffer[92] ),
    .A1(\deser_B.serial_word[92] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _13657_ (.A0(\deser_B.word_buffer[93] ),
    .A1(\deser_B.serial_word[93] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _13658_ (.A0(\deser_B.word_buffer[94] ),
    .A1(\deser_B.serial_word[94] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _13659_ (.A0(\deser_B.word_buffer[95] ),
    .A1(\deser_B.serial_word[95] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _13660_ (.A0(\deser_B.word_buffer[96] ),
    .A1(\deser_B.serial_word[96] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _13661_ (.A0(\deser_B.word_buffer[97] ),
    .A1(\deser_B.serial_word[97] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _13662_ (.A0(\deser_B.word_buffer[98] ),
    .A1(\deser_B.serial_word[98] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _13663_ (.A0(\deser_B.word_buffer[99] ),
    .A1(\deser_B.serial_word[99] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _13664_ (.A0(\deser_B.word_buffer[100] ),
    .A1(\deser_B.serial_word[100] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _13665_ (.A0(\deser_B.word_buffer[101] ),
    .A1(\deser_B.serial_word[101] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _13666_ (.A0(\deser_B.word_buffer[102] ),
    .A1(\deser_B.serial_word[102] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _13667_ (.A0(\deser_B.word_buffer[103] ),
    .A1(\deser_B.serial_word[103] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _13668_ (.A0(\deser_B.word_buffer[104] ),
    .A1(\deser_B.serial_word[104] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _13669_ (.A0(\deser_B.word_buffer[105] ),
    .A1(\deser_B.serial_word[105] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _13670_ (.A0(\deser_B.word_buffer[106] ),
    .A1(\deser_B.serial_word[106] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _13671_ (.A0(\deser_B.word_buffer[107] ),
    .A1(\deser_B.serial_word[107] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _13672_ (.A0(\deser_B.word_buffer[108] ),
    .A1(\deser_B.serial_word[108] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _13673_ (.A0(\deser_B.word_buffer[109] ),
    .A1(\deser_B.serial_word[109] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _13674_ (.A0(\deser_B.word_buffer[110] ),
    .A1(\deser_B.serial_word[110] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _13675_ (.A0(\deser_B.word_buffer[111] ),
    .A1(\deser_B.serial_word[111] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _13676_ (.A0(\deser_B.word_buffer[112] ),
    .A1(\deser_B.serial_word[112] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _13677_ (.A0(\deser_B.word_buffer[113] ),
    .A1(\deser_B.serial_word[113] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _13678_ (.A0(\deser_B.word_buffer[114] ),
    .A1(\deser_B.serial_word[114] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _13679_ (.A0(\deser_B.word_buffer[115] ),
    .A1(\deser_B.serial_word[115] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _13680_ (.A0(\deser_B.word_buffer[116] ),
    .A1(\deser_B.serial_word[116] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _13681_ (.A0(\deser_B.word_buffer[117] ),
    .A1(\deser_B.serial_word[117] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _13682_ (.A0(\deser_B.word_buffer[118] ),
    .A1(\deser_B.serial_word[118] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _13683_ (.A0(\deser_B.word_buffer[119] ),
    .A1(\deser_B.serial_word[119] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _13684_ (.A0(\deser_B.word_buffer[120] ),
    .A1(\deser_B.serial_word[120] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _13685_ (.A0(\deser_B.word_buffer[121] ),
    .A1(\deser_B.serial_word[121] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _13686_ (.A0(\deser_B.word_buffer[122] ),
    .A1(\deser_B.serial_word[122] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _13687_ (.A0(\deser_B.word_buffer[123] ),
    .A1(\deser_B.serial_word[123] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _13688_ (.A0(\deser_B.word_buffer[124] ),
    .A1(\deser_B.serial_word[124] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _13689_ (.A0(\deser_B.word_buffer[125] ),
    .A1(\deser_B.serial_word[125] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _13690_ (.A0(\deser_B.word_buffer[126] ),
    .A1(\deser_B.serial_word[126] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _13691_ (.A0(\deser_B.word_buffer[127] ),
    .A1(\deser_B.serial_word[127] ),
    .S(\deser_B.serial_word_ready ),
    .X(_00528_));
 sky130_fd_sc_hd__xor2_2 _13692_ (.A(\deser_B.serial_toggle ),
    .B(\deser_B.serial_word_ready ),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _13693_ (.A0(\B_in[0] ),
    .A1(\deser_B.word_buffer[0] ),
    .S(_00005_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _13694_ (.A0(\B_in[1] ),
    .A1(\deser_B.word_buffer[1] ),
    .S(_00005_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _13695_ (.A0(\B_in[2] ),
    .A1(\deser_B.word_buffer[2] ),
    .S(_00005_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _13696_ (.A0(\B_in[3] ),
    .A1(\deser_B.word_buffer[3] ),
    .S(_00005_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _13697_ (.A0(\B_in[4] ),
    .A1(\deser_B.word_buffer[4] ),
    .S(_00005_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _13698_ (.A0(\B_in[5] ),
    .A1(\deser_B.word_buffer[5] ),
    .S(_00005_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _13699_ (.A0(\B_in[6] ),
    .A1(\deser_B.word_buffer[6] ),
    .S(_00005_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _13700_ (.A0(\B_in[7] ),
    .A1(\deser_B.word_buffer[7] ),
    .S(_00005_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _13701_ (.A0(\B_in[8] ),
    .A1(\deser_B.word_buffer[8] ),
    .S(_00005_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _13702_ (.A0(\B_in[9] ),
    .A1(\deser_B.word_buffer[9] ),
    .S(_00005_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _13703_ (.A0(\B_in[10] ),
    .A1(\deser_B.word_buffer[10] ),
    .S(_00005_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _13704_ (.A0(\B_in[11] ),
    .A1(\deser_B.word_buffer[11] ),
    .S(_00005_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _13705_ (.A0(\B_in[12] ),
    .A1(\deser_B.word_buffer[12] ),
    .S(_00005_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _13706_ (.A0(\B_in[13] ),
    .A1(\deser_B.word_buffer[13] ),
    .S(_00005_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _13707_ (.A0(\B_in[14] ),
    .A1(\deser_B.word_buffer[14] ),
    .S(_00005_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _13708_ (.A0(\B_in[15] ),
    .A1(\deser_B.word_buffer[15] ),
    .S(_00005_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _13709_ (.A0(\B_in[16] ),
    .A1(\deser_B.word_buffer[16] ),
    .S(_00005_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _13710_ (.A0(\B_in[17] ),
    .A1(\deser_B.word_buffer[17] ),
    .S(_00005_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _13711_ (.A0(\B_in[18] ),
    .A1(\deser_B.word_buffer[18] ),
    .S(_00005_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _13712_ (.A0(\B_in[19] ),
    .A1(\deser_B.word_buffer[19] ),
    .S(_00005_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _13713_ (.A0(\B_in[20] ),
    .A1(\deser_B.word_buffer[20] ),
    .S(_00005_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _13714_ (.A0(\B_in[21] ),
    .A1(\deser_B.word_buffer[21] ),
    .S(_00005_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _13715_ (.A0(\B_in[22] ),
    .A1(\deser_B.word_buffer[22] ),
    .S(_00005_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _13716_ (.A0(\B_in[23] ),
    .A1(\deser_B.word_buffer[23] ),
    .S(_00005_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _13717_ (.A0(\B_in[24] ),
    .A1(\deser_B.word_buffer[24] ),
    .S(_00005_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _13718_ (.A0(\B_in[25] ),
    .A1(\deser_B.word_buffer[25] ),
    .S(_00005_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _13719_ (.A0(\B_in[26] ),
    .A1(\deser_B.word_buffer[26] ),
    .S(_00005_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _13720_ (.A0(\B_in[27] ),
    .A1(\deser_B.word_buffer[27] ),
    .S(_00005_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _13721_ (.A0(\B_in[28] ),
    .A1(\deser_B.word_buffer[28] ),
    .S(_00005_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _13722_ (.A0(\B_in[29] ),
    .A1(\deser_B.word_buffer[29] ),
    .S(_00005_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _13723_ (.A0(\B_in[30] ),
    .A1(\deser_B.word_buffer[30] ),
    .S(_00005_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _13724_ (.A0(\B_in[31] ),
    .A1(\deser_B.word_buffer[31] ),
    .S(_00005_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _13725_ (.A0(\B_in[32] ),
    .A1(\deser_B.word_buffer[32] ),
    .S(_00005_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _13726_ (.A0(\B_in[33] ),
    .A1(\deser_B.word_buffer[33] ),
    .S(_00005_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _13727_ (.A0(\B_in[34] ),
    .A1(\deser_B.word_buffer[34] ),
    .S(_00005_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _13728_ (.A0(\B_in[35] ),
    .A1(\deser_B.word_buffer[35] ),
    .S(_00005_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _13729_ (.A0(\B_in[36] ),
    .A1(\deser_B.word_buffer[36] ),
    .S(_00005_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _13730_ (.A0(\B_in[37] ),
    .A1(\deser_B.word_buffer[37] ),
    .S(_00005_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _13731_ (.A0(\B_in[38] ),
    .A1(\deser_B.word_buffer[38] ),
    .S(_00005_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _13732_ (.A0(\B_in[39] ),
    .A1(\deser_B.word_buffer[39] ),
    .S(_00005_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _13733_ (.A0(\B_in[40] ),
    .A1(\deser_B.word_buffer[40] ),
    .S(_00005_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _13734_ (.A0(\B_in[41] ),
    .A1(\deser_B.word_buffer[41] ),
    .S(_00005_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _13735_ (.A0(\B_in[42] ),
    .A1(\deser_B.word_buffer[42] ),
    .S(_00005_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _13736_ (.A0(\B_in[43] ),
    .A1(\deser_B.word_buffer[43] ),
    .S(_00005_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _13737_ (.A0(\B_in[44] ),
    .A1(\deser_B.word_buffer[44] ),
    .S(_00005_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _13738_ (.A0(\B_in[45] ),
    .A1(\deser_B.word_buffer[45] ),
    .S(_00005_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _13739_ (.A0(\B_in[46] ),
    .A1(\deser_B.word_buffer[46] ),
    .S(_00005_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _13740_ (.A0(\B_in[47] ),
    .A1(\deser_B.word_buffer[47] ),
    .S(_00005_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _13741_ (.A0(\B_in[48] ),
    .A1(\deser_B.word_buffer[48] ),
    .S(_00005_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _13742_ (.A0(\B_in[49] ),
    .A1(\deser_B.word_buffer[49] ),
    .S(_00005_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _13743_ (.A0(\B_in[50] ),
    .A1(\deser_B.word_buffer[50] ),
    .S(_00005_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _13744_ (.A0(\B_in[51] ),
    .A1(\deser_B.word_buffer[51] ),
    .S(_00005_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _13745_ (.A0(\B_in[52] ),
    .A1(\deser_B.word_buffer[52] ),
    .S(_00005_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _13746_ (.A0(\B_in[53] ),
    .A1(\deser_B.word_buffer[53] ),
    .S(_00005_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _13747_ (.A0(\B_in[54] ),
    .A1(\deser_B.word_buffer[54] ),
    .S(_00005_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _13748_ (.A0(\B_in[55] ),
    .A1(\deser_B.word_buffer[55] ),
    .S(_00005_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _13749_ (.A0(\B_in[56] ),
    .A1(\deser_B.word_buffer[56] ),
    .S(_00005_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _13750_ (.A0(\B_in[57] ),
    .A1(\deser_B.word_buffer[57] ),
    .S(_00005_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _13751_ (.A0(\B_in[58] ),
    .A1(\deser_B.word_buffer[58] ),
    .S(_00005_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _13752_ (.A0(\B_in[59] ),
    .A1(\deser_B.word_buffer[59] ),
    .S(_00005_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _13753_ (.A0(\B_in[60] ),
    .A1(\deser_B.word_buffer[60] ),
    .S(_00005_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _13754_ (.A0(\B_in[61] ),
    .A1(\deser_B.word_buffer[61] ),
    .S(_00005_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _13755_ (.A0(\B_in[62] ),
    .A1(\deser_B.word_buffer[62] ),
    .S(_00005_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _13756_ (.A0(\B_in[63] ),
    .A1(\deser_B.word_buffer[63] ),
    .S(_00005_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _13757_ (.A0(\B_in[64] ),
    .A1(\deser_B.word_buffer[64] ),
    .S(_00005_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _13758_ (.A0(\B_in[65] ),
    .A1(\deser_B.word_buffer[65] ),
    .S(_00005_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _13759_ (.A0(\B_in[66] ),
    .A1(\deser_B.word_buffer[66] ),
    .S(_00005_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _13760_ (.A0(\B_in[67] ),
    .A1(\deser_B.word_buffer[67] ),
    .S(_00005_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _13761_ (.A0(\B_in[68] ),
    .A1(\deser_B.word_buffer[68] ),
    .S(_00005_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _13762_ (.A0(\B_in[69] ),
    .A1(\deser_B.word_buffer[69] ),
    .S(_00005_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _13763_ (.A0(\B_in[70] ),
    .A1(\deser_B.word_buffer[70] ),
    .S(_00005_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _13764_ (.A0(\B_in[71] ),
    .A1(\deser_B.word_buffer[71] ),
    .S(_00005_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _13765_ (.A0(\B_in[72] ),
    .A1(\deser_B.word_buffer[72] ),
    .S(_00005_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _13766_ (.A0(\B_in[73] ),
    .A1(\deser_B.word_buffer[73] ),
    .S(_00005_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _13767_ (.A0(\B_in[74] ),
    .A1(\deser_B.word_buffer[74] ),
    .S(_00005_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _13768_ (.A0(\B_in[75] ),
    .A1(\deser_B.word_buffer[75] ),
    .S(_00005_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _13769_ (.A0(\B_in[76] ),
    .A1(\deser_B.word_buffer[76] ),
    .S(_00005_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _13770_ (.A0(\B_in[77] ),
    .A1(\deser_B.word_buffer[77] ),
    .S(_00005_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _13771_ (.A0(\B_in[78] ),
    .A1(\deser_B.word_buffer[78] ),
    .S(_00005_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _13772_ (.A0(\B_in[79] ),
    .A1(\deser_B.word_buffer[79] ),
    .S(_00005_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _13773_ (.A0(\B_in[80] ),
    .A1(\deser_B.word_buffer[80] ),
    .S(_00005_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _13774_ (.A0(\B_in[81] ),
    .A1(\deser_B.word_buffer[81] ),
    .S(_00005_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _13775_ (.A0(\B_in[82] ),
    .A1(\deser_B.word_buffer[82] ),
    .S(_00005_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _13776_ (.A0(\B_in[83] ),
    .A1(\deser_B.word_buffer[83] ),
    .S(_00005_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _13777_ (.A0(\B_in[84] ),
    .A1(\deser_B.word_buffer[84] ),
    .S(_00005_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _13778_ (.A0(\B_in[85] ),
    .A1(\deser_B.word_buffer[85] ),
    .S(_00005_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _13779_ (.A0(\B_in[86] ),
    .A1(\deser_B.word_buffer[86] ),
    .S(_00005_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _13780_ (.A0(\B_in[87] ),
    .A1(\deser_B.word_buffer[87] ),
    .S(_00005_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _13781_ (.A0(\B_in[88] ),
    .A1(\deser_B.word_buffer[88] ),
    .S(_00005_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _13782_ (.A0(\B_in[89] ),
    .A1(\deser_B.word_buffer[89] ),
    .S(_00005_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _13783_ (.A0(\B_in[90] ),
    .A1(\deser_B.word_buffer[90] ),
    .S(_00005_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _13784_ (.A0(\B_in[91] ),
    .A1(\deser_B.word_buffer[91] ),
    .S(_00005_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _13785_ (.A0(\B_in[92] ),
    .A1(\deser_B.word_buffer[92] ),
    .S(_00005_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _13786_ (.A0(\B_in[93] ),
    .A1(\deser_B.word_buffer[93] ),
    .S(_00005_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _13787_ (.A0(\B_in[94] ),
    .A1(\deser_B.word_buffer[94] ),
    .S(_00005_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _13788_ (.A0(\B_in[95] ),
    .A1(\deser_B.word_buffer[95] ),
    .S(_00005_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _13789_ (.A0(\B_in[96] ),
    .A1(\deser_B.word_buffer[96] ),
    .S(_00005_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _13790_ (.A0(\B_in[97] ),
    .A1(\deser_B.word_buffer[97] ),
    .S(_00005_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _13791_ (.A0(\B_in[98] ),
    .A1(\deser_B.word_buffer[98] ),
    .S(_00005_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _13792_ (.A0(\B_in[99] ),
    .A1(\deser_B.word_buffer[99] ),
    .S(_00005_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _13793_ (.A0(\B_in[100] ),
    .A1(\deser_B.word_buffer[100] ),
    .S(_00005_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _13794_ (.A0(\B_in[101] ),
    .A1(\deser_B.word_buffer[101] ),
    .S(_00005_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _13795_ (.A0(\B_in[102] ),
    .A1(\deser_B.word_buffer[102] ),
    .S(_00005_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _13796_ (.A0(\B_in[103] ),
    .A1(\deser_B.word_buffer[103] ),
    .S(_00005_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _13797_ (.A0(\B_in[104] ),
    .A1(\deser_B.word_buffer[104] ),
    .S(_00005_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _13798_ (.A0(\B_in[105] ),
    .A1(\deser_B.word_buffer[105] ),
    .S(_00005_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _13799_ (.A0(\B_in[106] ),
    .A1(\deser_B.word_buffer[106] ),
    .S(_00005_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _13800_ (.A0(\B_in[107] ),
    .A1(\deser_B.word_buffer[107] ),
    .S(_00005_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _13801_ (.A0(\B_in[108] ),
    .A1(\deser_B.word_buffer[108] ),
    .S(_00005_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _13802_ (.A0(\B_in[109] ),
    .A1(\deser_B.word_buffer[109] ),
    .S(_00005_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _13803_ (.A0(\B_in[110] ),
    .A1(\deser_B.word_buffer[110] ),
    .S(_00005_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _13804_ (.A0(\B_in[111] ),
    .A1(\deser_B.word_buffer[111] ),
    .S(_00005_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _13805_ (.A0(\B_in[112] ),
    .A1(\deser_B.word_buffer[112] ),
    .S(_00005_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _13806_ (.A0(\B_in[113] ),
    .A1(\deser_B.word_buffer[113] ),
    .S(_00005_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _13807_ (.A0(\B_in[114] ),
    .A1(\deser_B.word_buffer[114] ),
    .S(_00005_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _13808_ (.A0(\B_in[115] ),
    .A1(\deser_B.word_buffer[115] ),
    .S(_00005_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _13809_ (.A0(\B_in[116] ),
    .A1(\deser_B.word_buffer[116] ),
    .S(_00005_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _13810_ (.A0(\B_in[117] ),
    .A1(\deser_B.word_buffer[117] ),
    .S(_00005_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _13811_ (.A0(\B_in[118] ),
    .A1(\deser_B.word_buffer[118] ),
    .S(_00005_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _13812_ (.A0(\B_in[119] ),
    .A1(\deser_B.word_buffer[119] ),
    .S(_00005_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _13813_ (.A0(\B_in[120] ),
    .A1(\deser_B.word_buffer[120] ),
    .S(_00005_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _13814_ (.A0(\B_in[121] ),
    .A1(\deser_B.word_buffer[121] ),
    .S(_00005_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _13815_ (.A0(\B_in[122] ),
    .A1(\deser_B.word_buffer[122] ),
    .S(_00005_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _13816_ (.A0(\B_in[123] ),
    .A1(\deser_B.word_buffer[123] ),
    .S(_00005_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _13817_ (.A0(\B_in[124] ),
    .A1(\deser_B.word_buffer[124] ),
    .S(_00005_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _13818_ (.A0(\B_in[125] ),
    .A1(\deser_B.word_buffer[125] ),
    .S(_00005_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _13819_ (.A0(\B_in[126] ),
    .A1(\deser_B.word_buffer[126] ),
    .S(_00005_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _13820_ (.A0(\B_in[127] ),
    .A1(\deser_B.word_buffer[127] ),
    .S(_00005_),
    .X(_00657_));
 sky130_fd_sc_hd__o21a_2 _13821_ (.A1(B_in_frame_sync),
    .A2(\deser_B.receiving ),
    .B1(\deser_B.bit_idx[0] ),
    .X(_11319_));
 sky130_fd_sc_hd__o21ba_2 _13822_ (.A1(\deser_B.receiving ),
    .A2(\deser_B.bit_idx[0] ),
    .B1_N(_11319_),
    .X(_00658_));
 sky130_fd_sc_hd__and2_2 _13823_ (.A(\deser_B.bit_idx[1] ),
    .B(_11319_),
    .X(_11320_));
 sky130_fd_sc_hd__nand2b_2 _13824_ (.A_N(\deser_B.receiving ),
    .B(B_in_frame_sync),
    .Y(_11321_));
 sky130_fd_sc_hd__o21ai_2 _13825_ (.A1(\deser_B.bit_idx[1] ),
    .A2(_11319_),
    .B1(_11321_),
    .Y(_11322_));
 sky130_fd_sc_hd__nor2_2 _13826_ (.A(_11320_),
    .B(_11322_),
    .Y(_00659_));
 sky130_fd_sc_hd__and3_2 _13827_ (.A(\deser_B.bit_idx[1] ),
    .B(\deser_B.bit_idx[2] ),
    .C(_11319_),
    .X(_11323_));
 sky130_fd_sc_hd__o21ai_2 _13828_ (.A1(\deser_B.bit_idx[2] ),
    .A2(_11320_),
    .B1(_11321_),
    .Y(_11324_));
 sky130_fd_sc_hd__nor2_2 _13829_ (.A(_11323_),
    .B(_11324_),
    .Y(_00660_));
 sky130_fd_sc_hd__o21ai_2 _13830_ (.A1(\deser_B.bit_idx[3] ),
    .A2(_11323_),
    .B1(_11321_),
    .Y(_11325_));
 sky130_fd_sc_hd__a21oi_2 _13831_ (.A1(\deser_B.bit_idx[3] ),
    .A2(_11323_),
    .B1(_11325_),
    .Y(_00661_));
 sky130_fd_sc_hd__a31o_2 _13832_ (.A1(\deser_B.bit_idx[3] ),
    .A2(\deser_B.bit_idx[2] ),
    .A3(_11320_),
    .B1(\deser_B.bit_idx[4] ),
    .X(_11326_));
 sky130_fd_sc_hd__and3_2 _13833_ (.A(\deser_B.bit_idx[3] ),
    .B(\deser_B.bit_idx[4] ),
    .C(_11323_),
    .X(_11327_));
 sky130_fd_sc_hd__inv_2 _13834_ (.A(_11327_),
    .Y(_11328_));
 sky130_fd_sc_hd__and3_2 _13835_ (.A(_11321_),
    .B(_11326_),
    .C(_11328_),
    .X(_00662_));
 sky130_fd_sc_hd__o211a_2 _13836_ (.A1(\deser_B.bit_idx[5] ),
    .A2(_11327_),
    .B1(_11321_),
    .C1(_11285_),
    .X(_00663_));
 sky130_fd_sc_hd__a21o_2 _13837_ (.A1(\deser_B.bit_idx[5] ),
    .A2(_11327_),
    .B1(\deser_B.bit_idx[6] ),
    .X(_11329_));
 sky130_fd_sc_hd__and3b_2 _13838_ (.A_N(_00001_),
    .B(_11321_),
    .C(_11329_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _13839_ (.A0(\deser_A.serial_word[0] ),
    .A1(\deser_A.shift_reg[0] ),
    .S(_00002_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _13840_ (.A0(\deser_A.serial_word[1] ),
    .A1(\deser_A.shift_reg[1] ),
    .S(_00002_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _13841_ (.A0(\deser_A.serial_word[2] ),
    .A1(\deser_A.shift_reg[2] ),
    .S(_00002_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _13842_ (.A0(\deser_A.serial_word[3] ),
    .A1(\deser_A.shift_reg[3] ),
    .S(_00002_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _13843_ (.A0(\deser_A.serial_word[4] ),
    .A1(\deser_A.shift_reg[4] ),
    .S(_00002_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _13844_ (.A0(\deser_A.serial_word[5] ),
    .A1(\deser_A.shift_reg[5] ),
    .S(_00002_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _13845_ (.A0(\deser_A.serial_word[6] ),
    .A1(\deser_A.shift_reg[6] ),
    .S(_00002_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _13846_ (.A0(\deser_A.serial_word[7] ),
    .A1(\deser_A.shift_reg[7] ),
    .S(_00002_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _13847_ (.A0(\deser_A.serial_word[8] ),
    .A1(\deser_A.shift_reg[8] ),
    .S(_00002_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _13848_ (.A0(\deser_A.serial_word[9] ),
    .A1(\deser_A.shift_reg[9] ),
    .S(_00002_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _13849_ (.A0(\deser_A.serial_word[10] ),
    .A1(\deser_A.shift_reg[10] ),
    .S(_00002_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _13850_ (.A0(\deser_A.serial_word[11] ),
    .A1(\deser_A.shift_reg[11] ),
    .S(_00002_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _13851_ (.A0(\deser_A.serial_word[12] ),
    .A1(\deser_A.shift_reg[12] ),
    .S(_00002_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _13852_ (.A0(\deser_A.serial_word[13] ),
    .A1(\deser_A.shift_reg[13] ),
    .S(_00002_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _13853_ (.A0(\deser_A.serial_word[14] ),
    .A1(\deser_A.shift_reg[14] ),
    .S(_00002_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _13854_ (.A0(\deser_A.serial_word[15] ),
    .A1(\deser_A.shift_reg[15] ),
    .S(_00002_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _13855_ (.A0(\deser_A.serial_word[16] ),
    .A1(\deser_A.shift_reg[16] ),
    .S(_00002_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _13856_ (.A0(\deser_A.serial_word[17] ),
    .A1(\deser_A.shift_reg[17] ),
    .S(_00002_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _13857_ (.A0(\deser_A.serial_word[18] ),
    .A1(\deser_A.shift_reg[18] ),
    .S(_00002_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _13858_ (.A0(\deser_A.serial_word[19] ),
    .A1(\deser_A.shift_reg[19] ),
    .S(_00002_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _13859_ (.A0(\deser_A.serial_word[20] ),
    .A1(\deser_A.shift_reg[20] ),
    .S(_00002_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _13860_ (.A0(\deser_A.serial_word[21] ),
    .A1(\deser_A.shift_reg[21] ),
    .S(_00002_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _13861_ (.A0(\deser_A.serial_word[22] ),
    .A1(\deser_A.shift_reg[22] ),
    .S(_00002_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _13862_ (.A0(\deser_A.serial_word[23] ),
    .A1(\deser_A.shift_reg[23] ),
    .S(_00002_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _13863_ (.A0(\deser_A.serial_word[24] ),
    .A1(\deser_A.shift_reg[24] ),
    .S(_00002_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _13864_ (.A0(\deser_A.serial_word[25] ),
    .A1(\deser_A.shift_reg[25] ),
    .S(_00002_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _13865_ (.A0(\deser_A.serial_word[26] ),
    .A1(\deser_A.shift_reg[26] ),
    .S(_00002_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _13866_ (.A0(\deser_A.serial_word[27] ),
    .A1(\deser_A.shift_reg[27] ),
    .S(_00002_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _13867_ (.A0(\deser_A.serial_word[28] ),
    .A1(\deser_A.shift_reg[28] ),
    .S(_00002_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _13868_ (.A0(\deser_A.serial_word[29] ),
    .A1(\deser_A.shift_reg[29] ),
    .S(_00002_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _13869_ (.A0(\deser_A.serial_word[30] ),
    .A1(\deser_A.shift_reg[30] ),
    .S(_00002_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _13870_ (.A0(\deser_A.serial_word[31] ),
    .A1(\deser_A.shift_reg[31] ),
    .S(_00002_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _13871_ (.A0(\deser_A.serial_word[32] ),
    .A1(\deser_A.shift_reg[32] ),
    .S(_00002_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _13872_ (.A0(\deser_A.serial_word[33] ),
    .A1(\deser_A.shift_reg[33] ),
    .S(_00002_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _13873_ (.A0(\deser_A.serial_word[34] ),
    .A1(\deser_A.shift_reg[34] ),
    .S(_00002_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _13874_ (.A0(\deser_A.serial_word[35] ),
    .A1(\deser_A.shift_reg[35] ),
    .S(_00002_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _13875_ (.A0(\deser_A.serial_word[36] ),
    .A1(\deser_A.shift_reg[36] ),
    .S(_00002_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _13876_ (.A0(\deser_A.serial_word[37] ),
    .A1(\deser_A.shift_reg[37] ),
    .S(_00002_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _13877_ (.A0(\deser_A.serial_word[38] ),
    .A1(\deser_A.shift_reg[38] ),
    .S(_00002_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _13878_ (.A0(\deser_A.serial_word[39] ),
    .A1(\deser_A.shift_reg[39] ),
    .S(_00002_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _13879_ (.A0(\deser_A.serial_word[40] ),
    .A1(\deser_A.shift_reg[40] ),
    .S(_00002_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _13880_ (.A0(\deser_A.serial_word[41] ),
    .A1(\deser_A.shift_reg[41] ),
    .S(_00002_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _13881_ (.A0(\deser_A.serial_word[42] ),
    .A1(\deser_A.shift_reg[42] ),
    .S(_00002_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _13882_ (.A0(\deser_A.serial_word[43] ),
    .A1(\deser_A.shift_reg[43] ),
    .S(_00002_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _13883_ (.A0(\deser_A.serial_word[44] ),
    .A1(\deser_A.shift_reg[44] ),
    .S(_00002_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _13884_ (.A0(\deser_A.serial_word[45] ),
    .A1(\deser_A.shift_reg[45] ),
    .S(_00002_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _13885_ (.A0(\deser_A.serial_word[46] ),
    .A1(\deser_A.shift_reg[46] ),
    .S(_00002_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _13886_ (.A0(\deser_A.serial_word[47] ),
    .A1(\deser_A.shift_reg[47] ),
    .S(_00002_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _13887_ (.A0(\deser_A.serial_word[48] ),
    .A1(\deser_A.shift_reg[48] ),
    .S(_00002_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _13888_ (.A0(\deser_A.serial_word[49] ),
    .A1(\deser_A.shift_reg[49] ),
    .S(_00002_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _13889_ (.A0(\deser_A.serial_word[50] ),
    .A1(\deser_A.shift_reg[50] ),
    .S(_00002_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _13890_ (.A0(\deser_A.serial_word[51] ),
    .A1(\deser_A.shift_reg[51] ),
    .S(_00002_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _13891_ (.A0(\deser_A.serial_word[52] ),
    .A1(\deser_A.shift_reg[52] ),
    .S(_00002_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _13892_ (.A0(\deser_A.serial_word[53] ),
    .A1(\deser_A.shift_reg[53] ),
    .S(_00002_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _13893_ (.A0(\deser_A.serial_word[54] ),
    .A1(\deser_A.shift_reg[54] ),
    .S(_00002_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _13894_ (.A0(\deser_A.serial_word[55] ),
    .A1(\deser_A.shift_reg[55] ),
    .S(_00002_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _13895_ (.A0(\deser_A.serial_word[56] ),
    .A1(\deser_A.shift_reg[56] ),
    .S(_00002_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _13896_ (.A0(\deser_A.serial_word[57] ),
    .A1(\deser_A.shift_reg[57] ),
    .S(_00002_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _13897_ (.A0(\deser_A.serial_word[58] ),
    .A1(\deser_A.shift_reg[58] ),
    .S(_00002_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _13898_ (.A0(\deser_A.serial_word[59] ),
    .A1(\deser_A.shift_reg[59] ),
    .S(_00002_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _13899_ (.A0(\deser_A.serial_word[60] ),
    .A1(\deser_A.shift_reg[60] ),
    .S(_00002_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _13900_ (.A0(\deser_A.serial_word[61] ),
    .A1(\deser_A.shift_reg[61] ),
    .S(_00002_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _13901_ (.A0(\deser_A.serial_word[62] ),
    .A1(\deser_A.shift_reg[62] ),
    .S(_00002_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _13902_ (.A0(\deser_A.serial_word[63] ),
    .A1(\deser_A.shift_reg[63] ),
    .S(_00002_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _13903_ (.A0(\deser_A.serial_word[64] ),
    .A1(\deser_A.shift_reg[64] ),
    .S(_00002_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _13904_ (.A0(\deser_A.serial_word[65] ),
    .A1(\deser_A.shift_reg[65] ),
    .S(_00002_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _13905_ (.A0(\deser_A.serial_word[66] ),
    .A1(\deser_A.shift_reg[66] ),
    .S(_00002_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _13906_ (.A0(\deser_A.serial_word[67] ),
    .A1(\deser_A.shift_reg[67] ),
    .S(_00002_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _13907_ (.A0(\deser_A.serial_word[68] ),
    .A1(\deser_A.shift_reg[68] ),
    .S(_00002_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _13908_ (.A0(\deser_A.serial_word[69] ),
    .A1(\deser_A.shift_reg[69] ),
    .S(_00002_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _13909_ (.A0(\deser_A.serial_word[70] ),
    .A1(\deser_A.shift_reg[70] ),
    .S(_00002_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _13910_ (.A0(\deser_A.serial_word[71] ),
    .A1(\deser_A.shift_reg[71] ),
    .S(_00002_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _13911_ (.A0(\deser_A.serial_word[72] ),
    .A1(\deser_A.shift_reg[72] ),
    .S(_00002_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _13912_ (.A0(\deser_A.serial_word[73] ),
    .A1(\deser_A.shift_reg[73] ),
    .S(_00002_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _13913_ (.A0(\deser_A.serial_word[74] ),
    .A1(\deser_A.shift_reg[74] ),
    .S(_00002_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _13914_ (.A0(\deser_A.serial_word[75] ),
    .A1(\deser_A.shift_reg[75] ),
    .S(_00002_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _13915_ (.A0(\deser_A.serial_word[76] ),
    .A1(\deser_A.shift_reg[76] ),
    .S(_00002_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _13916_ (.A0(\deser_A.serial_word[77] ),
    .A1(\deser_A.shift_reg[77] ),
    .S(_00002_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _13917_ (.A0(\deser_A.serial_word[78] ),
    .A1(\deser_A.shift_reg[78] ),
    .S(_00002_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _13918_ (.A0(\deser_A.serial_word[79] ),
    .A1(\deser_A.shift_reg[79] ),
    .S(_00002_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _13919_ (.A0(\deser_A.serial_word[80] ),
    .A1(\deser_A.shift_reg[80] ),
    .S(_00002_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _13920_ (.A0(\deser_A.serial_word[81] ),
    .A1(\deser_A.shift_reg[81] ),
    .S(_00002_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _13921_ (.A0(\deser_A.serial_word[82] ),
    .A1(\deser_A.shift_reg[82] ),
    .S(_00002_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _13922_ (.A0(\deser_A.serial_word[83] ),
    .A1(\deser_A.shift_reg[83] ),
    .S(_00002_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _13923_ (.A0(\deser_A.serial_word[84] ),
    .A1(\deser_A.shift_reg[84] ),
    .S(_00002_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _13924_ (.A0(\deser_A.serial_word[85] ),
    .A1(\deser_A.shift_reg[85] ),
    .S(_00002_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _13925_ (.A0(\deser_A.serial_word[86] ),
    .A1(\deser_A.shift_reg[86] ),
    .S(_00002_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _13926_ (.A0(\deser_A.serial_word[87] ),
    .A1(\deser_A.shift_reg[87] ),
    .S(_00002_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _13927_ (.A0(\deser_A.serial_word[88] ),
    .A1(\deser_A.shift_reg[88] ),
    .S(_00002_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _13928_ (.A0(\deser_A.serial_word[89] ),
    .A1(\deser_A.shift_reg[89] ),
    .S(_00002_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _13929_ (.A0(\deser_A.serial_word[90] ),
    .A1(\deser_A.shift_reg[90] ),
    .S(_00002_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _13930_ (.A0(\deser_A.serial_word[91] ),
    .A1(\deser_A.shift_reg[91] ),
    .S(_00002_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _13931_ (.A0(\deser_A.serial_word[92] ),
    .A1(\deser_A.shift_reg[92] ),
    .S(_00002_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _13932_ (.A0(\deser_A.serial_word[93] ),
    .A1(\deser_A.shift_reg[93] ),
    .S(_00002_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _13933_ (.A0(\deser_A.serial_word[94] ),
    .A1(\deser_A.shift_reg[94] ),
    .S(_00002_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _13934_ (.A0(\deser_A.serial_word[95] ),
    .A1(\deser_A.shift_reg[95] ),
    .S(_00002_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _13935_ (.A0(\deser_A.serial_word[96] ),
    .A1(\deser_A.shift_reg[96] ),
    .S(_00002_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _13936_ (.A0(\deser_A.serial_word[97] ),
    .A1(\deser_A.shift_reg[97] ),
    .S(_00002_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _13937_ (.A0(\deser_A.serial_word[98] ),
    .A1(\deser_A.shift_reg[98] ),
    .S(_00002_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _13938_ (.A0(\deser_A.serial_word[99] ),
    .A1(\deser_A.shift_reg[99] ),
    .S(_00002_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _13939_ (.A0(\deser_A.serial_word[100] ),
    .A1(\deser_A.shift_reg[100] ),
    .S(_00002_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _13940_ (.A0(\deser_A.serial_word[101] ),
    .A1(\deser_A.shift_reg[101] ),
    .S(_00002_),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _13941_ (.A0(\deser_A.serial_word[102] ),
    .A1(\deser_A.shift_reg[102] ),
    .S(_00002_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _13942_ (.A0(\deser_A.serial_word[103] ),
    .A1(\deser_A.shift_reg[103] ),
    .S(_00002_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _13943_ (.A0(\deser_A.serial_word[104] ),
    .A1(\deser_A.shift_reg[104] ),
    .S(_00002_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _13944_ (.A0(\deser_A.serial_word[105] ),
    .A1(\deser_A.shift_reg[105] ),
    .S(_00002_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _13945_ (.A0(\deser_A.serial_word[106] ),
    .A1(\deser_A.shift_reg[106] ),
    .S(_00002_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _13946_ (.A0(\deser_A.serial_word[107] ),
    .A1(\deser_A.shift_reg[107] ),
    .S(_00002_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _13947_ (.A0(\deser_A.serial_word[108] ),
    .A1(\deser_A.shift_reg[108] ),
    .S(_00002_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _13948_ (.A0(\deser_A.serial_word[109] ),
    .A1(\deser_A.shift_reg[109] ),
    .S(_00002_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _13949_ (.A0(\deser_A.serial_word[110] ),
    .A1(\deser_A.shift_reg[110] ),
    .S(_00002_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _13950_ (.A0(\deser_A.serial_word[111] ),
    .A1(\deser_A.shift_reg[111] ),
    .S(_00002_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _13951_ (.A0(\deser_A.serial_word[112] ),
    .A1(\deser_A.shift_reg[112] ),
    .S(_00002_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _13952_ (.A0(\deser_A.serial_word[113] ),
    .A1(\deser_A.shift_reg[113] ),
    .S(_00002_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _13953_ (.A0(\deser_A.serial_word[114] ),
    .A1(\deser_A.shift_reg[114] ),
    .S(_00002_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _13954_ (.A0(\deser_A.serial_word[115] ),
    .A1(\deser_A.shift_reg[115] ),
    .S(_00002_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _13955_ (.A0(\deser_A.serial_word[116] ),
    .A1(\deser_A.shift_reg[116] ),
    .S(_00002_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _13956_ (.A0(\deser_A.serial_word[117] ),
    .A1(\deser_A.shift_reg[117] ),
    .S(_00002_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _13957_ (.A0(\deser_A.serial_word[118] ),
    .A1(\deser_A.shift_reg[118] ),
    .S(_00002_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _13958_ (.A0(\deser_A.serial_word[119] ),
    .A1(\deser_A.shift_reg[119] ),
    .S(_00002_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _13959_ (.A0(\deser_A.serial_word[120] ),
    .A1(\deser_A.shift_reg[120] ),
    .S(_00002_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _13960_ (.A0(\deser_A.serial_word[121] ),
    .A1(\deser_A.shift_reg[121] ),
    .S(_00002_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _13961_ (.A0(\deser_A.serial_word[122] ),
    .A1(\deser_A.shift_reg[122] ),
    .S(_00002_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _13962_ (.A0(\deser_A.serial_word[123] ),
    .A1(\deser_A.shift_reg[123] ),
    .S(_00002_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _13963_ (.A0(\deser_A.serial_word[124] ),
    .A1(\deser_A.shift_reg[124] ),
    .S(_00002_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _13964_ (.A0(\deser_A.serial_word[125] ),
    .A1(\deser_A.shift_reg[125] ),
    .S(_00002_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _13965_ (.A0(\deser_A.serial_word[126] ),
    .A1(\deser_A.shift_reg[126] ),
    .S(_00002_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _13966_ (.A0(\deser_A.serial_word[127] ),
    .A1(\deser_A.shift_reg[127] ),
    .S(_00002_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _13967_ (.A0(\deser_B.shift_reg[1] ),
    .A1(\deser_B.shift_reg[2] ),
    .S(\deser_B.receiving ),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _13968_ (.A0(\deser_B.shift_reg[2] ),
    .A1(\deser_B.shift_reg[3] ),
    .S(\deser_B.receiving ),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _13969_ (.A0(\deser_B.shift_reg[3] ),
    .A1(\deser_B.shift_reg[4] ),
    .S(\deser_B.receiving ),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _13970_ (.A0(\deser_B.shift_reg[4] ),
    .A1(\deser_B.shift_reg[5] ),
    .S(\deser_B.receiving ),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _13971_ (.A0(\deser_B.shift_reg[5] ),
    .A1(\deser_B.shift_reg[6] ),
    .S(\deser_B.receiving ),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _13972_ (.A0(\deser_B.shift_reg[6] ),
    .A1(\deser_B.shift_reg[7] ),
    .S(\deser_B.receiving ),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _13973_ (.A0(\deser_B.shift_reg[7] ),
    .A1(\deser_B.shift_reg[8] ),
    .S(\deser_B.receiving ),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _13974_ (.A0(\deser_B.shift_reg[8] ),
    .A1(\deser_B.shift_reg[9] ),
    .S(\deser_B.receiving ),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _13975_ (.A0(\deser_B.shift_reg[9] ),
    .A1(\deser_B.shift_reg[10] ),
    .S(\deser_B.receiving ),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _13976_ (.A0(\deser_B.shift_reg[10] ),
    .A1(\deser_B.shift_reg[11] ),
    .S(\deser_B.receiving ),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _13977_ (.A0(\deser_B.shift_reg[11] ),
    .A1(\deser_B.shift_reg[12] ),
    .S(\deser_B.receiving ),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _13978_ (.A0(\deser_B.shift_reg[12] ),
    .A1(\deser_B.shift_reg[13] ),
    .S(\deser_B.receiving ),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _13979_ (.A0(\deser_B.shift_reg[13] ),
    .A1(\deser_B.shift_reg[14] ),
    .S(\deser_B.receiving ),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _13980_ (.A0(\deser_B.shift_reg[14] ),
    .A1(\deser_B.shift_reg[15] ),
    .S(\deser_B.receiving ),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _13981_ (.A0(\deser_B.shift_reg[15] ),
    .A1(\deser_B.shift_reg[16] ),
    .S(\deser_B.receiving ),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _13982_ (.A0(\deser_B.shift_reg[16] ),
    .A1(\deser_B.shift_reg[17] ),
    .S(\deser_B.receiving ),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _13983_ (.A0(\deser_B.shift_reg[17] ),
    .A1(\deser_B.shift_reg[18] ),
    .S(\deser_B.receiving ),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _13984_ (.A0(\deser_B.shift_reg[18] ),
    .A1(\deser_B.shift_reg[19] ),
    .S(\deser_B.receiving ),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _13985_ (.A0(\deser_B.shift_reg[19] ),
    .A1(\deser_B.shift_reg[20] ),
    .S(\deser_B.receiving ),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _13986_ (.A0(\deser_B.shift_reg[20] ),
    .A1(\deser_B.shift_reg[21] ),
    .S(\deser_B.receiving ),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _13987_ (.A0(\deser_B.shift_reg[21] ),
    .A1(\deser_B.shift_reg[22] ),
    .S(\deser_B.receiving ),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _13988_ (.A0(\deser_B.shift_reg[22] ),
    .A1(\deser_B.shift_reg[23] ),
    .S(\deser_B.receiving ),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _13989_ (.A0(\deser_B.shift_reg[23] ),
    .A1(\deser_B.shift_reg[24] ),
    .S(\deser_B.receiving ),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _13990_ (.A0(\deser_B.shift_reg[24] ),
    .A1(\deser_B.shift_reg[25] ),
    .S(\deser_B.receiving ),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _13991_ (.A0(\deser_B.shift_reg[25] ),
    .A1(\deser_B.shift_reg[26] ),
    .S(\deser_B.receiving ),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _13992_ (.A0(\deser_B.shift_reg[26] ),
    .A1(\deser_B.shift_reg[27] ),
    .S(\deser_B.receiving ),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _13993_ (.A0(\deser_B.shift_reg[27] ),
    .A1(\deser_B.shift_reg[28] ),
    .S(\deser_B.receiving ),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _13994_ (.A0(\deser_B.shift_reg[28] ),
    .A1(\deser_B.shift_reg[29] ),
    .S(\deser_B.receiving ),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _13995_ (.A0(\deser_B.shift_reg[29] ),
    .A1(\deser_B.shift_reg[30] ),
    .S(\deser_B.receiving ),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _13996_ (.A0(\deser_B.shift_reg[30] ),
    .A1(\deser_B.shift_reg[31] ),
    .S(\deser_B.receiving ),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _13997_ (.A0(\deser_B.shift_reg[31] ),
    .A1(\deser_B.shift_reg[32] ),
    .S(\deser_B.receiving ),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _13998_ (.A0(\deser_B.shift_reg[32] ),
    .A1(\deser_B.shift_reg[33] ),
    .S(\deser_B.receiving ),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _13999_ (.A0(\deser_B.shift_reg[33] ),
    .A1(\deser_B.shift_reg[34] ),
    .S(\deser_B.receiving ),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _14000_ (.A0(\deser_B.shift_reg[34] ),
    .A1(\deser_B.shift_reg[35] ),
    .S(\deser_B.receiving ),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _14001_ (.A0(\deser_B.shift_reg[35] ),
    .A1(\deser_B.shift_reg[36] ),
    .S(\deser_B.receiving ),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _14002_ (.A0(\deser_B.shift_reg[36] ),
    .A1(\deser_B.shift_reg[37] ),
    .S(\deser_B.receiving ),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _14003_ (.A0(\deser_B.shift_reg[37] ),
    .A1(\deser_B.shift_reg[38] ),
    .S(\deser_B.receiving ),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _14004_ (.A0(\deser_B.shift_reg[38] ),
    .A1(\deser_B.shift_reg[39] ),
    .S(\deser_B.receiving ),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _14005_ (.A0(\deser_B.shift_reg[39] ),
    .A1(\deser_B.shift_reg[40] ),
    .S(\deser_B.receiving ),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _14006_ (.A0(\deser_B.shift_reg[40] ),
    .A1(\deser_B.shift_reg[41] ),
    .S(\deser_B.receiving ),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _14007_ (.A0(\deser_B.shift_reg[41] ),
    .A1(\deser_B.shift_reg[42] ),
    .S(\deser_B.receiving ),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _14008_ (.A0(\deser_B.shift_reg[42] ),
    .A1(\deser_B.shift_reg[43] ),
    .S(\deser_B.receiving ),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _14009_ (.A0(\deser_B.shift_reg[43] ),
    .A1(\deser_B.shift_reg[44] ),
    .S(\deser_B.receiving ),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _14010_ (.A0(\deser_B.shift_reg[44] ),
    .A1(\deser_B.shift_reg[45] ),
    .S(\deser_B.receiving ),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _14011_ (.A0(\deser_B.shift_reg[45] ),
    .A1(\deser_B.shift_reg[46] ),
    .S(\deser_B.receiving ),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _14012_ (.A0(\deser_B.shift_reg[46] ),
    .A1(\deser_B.shift_reg[47] ),
    .S(\deser_B.receiving ),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _14013_ (.A0(\deser_B.shift_reg[47] ),
    .A1(\deser_B.shift_reg[48] ),
    .S(\deser_B.receiving ),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _14014_ (.A0(\deser_B.shift_reg[48] ),
    .A1(\deser_B.shift_reg[49] ),
    .S(\deser_B.receiving ),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _14015_ (.A0(\deser_B.shift_reg[49] ),
    .A1(\deser_B.shift_reg[50] ),
    .S(\deser_B.receiving ),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _14016_ (.A0(\deser_B.shift_reg[50] ),
    .A1(\deser_B.shift_reg[51] ),
    .S(\deser_B.receiving ),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _14017_ (.A0(\deser_B.shift_reg[51] ),
    .A1(\deser_B.shift_reg[52] ),
    .S(\deser_B.receiving ),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _14018_ (.A0(\deser_B.shift_reg[52] ),
    .A1(\deser_B.shift_reg[53] ),
    .S(\deser_B.receiving ),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _14019_ (.A0(\deser_B.shift_reg[53] ),
    .A1(\deser_B.shift_reg[54] ),
    .S(\deser_B.receiving ),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _14020_ (.A0(\deser_B.shift_reg[54] ),
    .A1(\deser_B.shift_reg[55] ),
    .S(\deser_B.receiving ),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _14021_ (.A0(\deser_B.shift_reg[55] ),
    .A1(\deser_B.shift_reg[56] ),
    .S(\deser_B.receiving ),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _14022_ (.A0(\deser_B.shift_reg[56] ),
    .A1(\deser_B.shift_reg[57] ),
    .S(\deser_B.receiving ),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _14023_ (.A0(\deser_B.shift_reg[57] ),
    .A1(\deser_B.shift_reg[58] ),
    .S(\deser_B.receiving ),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _14024_ (.A0(\deser_B.shift_reg[58] ),
    .A1(\deser_B.shift_reg[59] ),
    .S(\deser_B.receiving ),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _14025_ (.A0(\deser_B.shift_reg[59] ),
    .A1(\deser_B.shift_reg[60] ),
    .S(\deser_B.receiving ),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _14026_ (.A0(\deser_B.shift_reg[60] ),
    .A1(\deser_B.shift_reg[61] ),
    .S(\deser_B.receiving ),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _14027_ (.A0(\deser_B.shift_reg[61] ),
    .A1(\deser_B.shift_reg[62] ),
    .S(\deser_B.receiving ),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _14028_ (.A0(\deser_B.shift_reg[62] ),
    .A1(\deser_B.shift_reg[63] ),
    .S(\deser_B.receiving ),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _14029_ (.A0(\deser_B.shift_reg[63] ),
    .A1(\deser_B.shift_reg[64] ),
    .S(\deser_B.receiving ),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _14030_ (.A0(\deser_B.shift_reg[64] ),
    .A1(\deser_B.shift_reg[65] ),
    .S(\deser_B.receiving ),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _14031_ (.A0(\deser_B.shift_reg[65] ),
    .A1(\deser_B.shift_reg[66] ),
    .S(\deser_B.receiving ),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _14032_ (.A0(\deser_B.shift_reg[66] ),
    .A1(\deser_B.shift_reg[67] ),
    .S(\deser_B.receiving ),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _14033_ (.A0(\deser_B.shift_reg[67] ),
    .A1(\deser_B.shift_reg[68] ),
    .S(\deser_B.receiving ),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _14034_ (.A0(\deser_B.shift_reg[68] ),
    .A1(\deser_B.shift_reg[69] ),
    .S(\deser_B.receiving ),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _14035_ (.A0(\deser_B.shift_reg[69] ),
    .A1(\deser_B.shift_reg[70] ),
    .S(\deser_B.receiving ),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _14036_ (.A0(\deser_B.shift_reg[70] ),
    .A1(\deser_B.shift_reg[71] ),
    .S(\deser_B.receiving ),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _14037_ (.A0(\deser_B.shift_reg[71] ),
    .A1(\deser_B.shift_reg[72] ),
    .S(\deser_B.receiving ),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _14038_ (.A0(\deser_B.shift_reg[72] ),
    .A1(\deser_B.shift_reg[73] ),
    .S(\deser_B.receiving ),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _14039_ (.A0(\deser_B.shift_reg[73] ),
    .A1(\deser_B.shift_reg[74] ),
    .S(\deser_B.receiving ),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _14040_ (.A0(\deser_B.shift_reg[74] ),
    .A1(\deser_B.shift_reg[75] ),
    .S(\deser_B.receiving ),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _14041_ (.A0(\deser_B.shift_reg[75] ),
    .A1(\deser_B.shift_reg[76] ),
    .S(\deser_B.receiving ),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _14042_ (.A0(\deser_B.shift_reg[76] ),
    .A1(\deser_B.shift_reg[77] ),
    .S(\deser_B.receiving ),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _14043_ (.A0(\deser_B.shift_reg[77] ),
    .A1(\deser_B.shift_reg[78] ),
    .S(\deser_B.receiving ),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _14044_ (.A0(\deser_B.shift_reg[78] ),
    .A1(\deser_B.shift_reg[79] ),
    .S(\deser_B.receiving ),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _14045_ (.A0(\deser_B.shift_reg[79] ),
    .A1(\deser_B.shift_reg[80] ),
    .S(\deser_B.receiving ),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _14046_ (.A0(\deser_B.shift_reg[80] ),
    .A1(\deser_B.shift_reg[81] ),
    .S(\deser_B.receiving ),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _14047_ (.A0(\deser_B.shift_reg[81] ),
    .A1(\deser_B.shift_reg[82] ),
    .S(\deser_B.receiving ),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _14048_ (.A0(\deser_B.shift_reg[82] ),
    .A1(\deser_B.shift_reg[83] ),
    .S(\deser_B.receiving ),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _14049_ (.A0(\deser_B.shift_reg[83] ),
    .A1(\deser_B.shift_reg[84] ),
    .S(\deser_B.receiving ),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _14050_ (.A0(\deser_B.shift_reg[84] ),
    .A1(\deser_B.shift_reg[85] ),
    .S(\deser_B.receiving ),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _14051_ (.A0(\deser_B.shift_reg[85] ),
    .A1(\deser_B.shift_reg[86] ),
    .S(\deser_B.receiving ),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _14052_ (.A0(\deser_B.shift_reg[86] ),
    .A1(\deser_B.shift_reg[87] ),
    .S(\deser_B.receiving ),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _14053_ (.A0(\deser_B.shift_reg[87] ),
    .A1(\deser_B.shift_reg[88] ),
    .S(\deser_B.receiving ),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _14054_ (.A0(\deser_B.shift_reg[88] ),
    .A1(\deser_B.shift_reg[89] ),
    .S(\deser_B.receiving ),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _14055_ (.A0(\deser_B.shift_reg[89] ),
    .A1(\deser_B.shift_reg[90] ),
    .S(\deser_B.receiving ),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _14056_ (.A0(\deser_B.shift_reg[90] ),
    .A1(\deser_B.shift_reg[91] ),
    .S(\deser_B.receiving ),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _14057_ (.A0(\deser_B.shift_reg[91] ),
    .A1(\deser_B.shift_reg[92] ),
    .S(\deser_B.receiving ),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _14058_ (.A0(\deser_B.shift_reg[92] ),
    .A1(\deser_B.shift_reg[93] ),
    .S(\deser_B.receiving ),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _14059_ (.A0(\deser_B.shift_reg[93] ),
    .A1(\deser_B.shift_reg[94] ),
    .S(\deser_B.receiving ),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _14060_ (.A0(\deser_B.shift_reg[94] ),
    .A1(\deser_B.shift_reg[95] ),
    .S(\deser_B.receiving ),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _14061_ (.A0(\deser_B.shift_reg[95] ),
    .A1(\deser_B.shift_reg[96] ),
    .S(\deser_B.receiving ),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _14062_ (.A0(\deser_B.shift_reg[96] ),
    .A1(\deser_B.shift_reg[97] ),
    .S(\deser_B.receiving ),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _14063_ (.A0(\deser_B.shift_reg[97] ),
    .A1(\deser_B.shift_reg[98] ),
    .S(\deser_B.receiving ),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _14064_ (.A0(\deser_B.shift_reg[98] ),
    .A1(\deser_B.shift_reg[99] ),
    .S(\deser_B.receiving ),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _14065_ (.A0(\deser_B.shift_reg[99] ),
    .A1(\deser_B.shift_reg[100] ),
    .S(\deser_B.receiving ),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _14066_ (.A0(\deser_B.shift_reg[100] ),
    .A1(\deser_B.shift_reg[101] ),
    .S(\deser_B.receiving ),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _14067_ (.A0(\deser_B.shift_reg[101] ),
    .A1(\deser_B.shift_reg[102] ),
    .S(\deser_B.receiving ),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _14068_ (.A0(\deser_B.shift_reg[102] ),
    .A1(\deser_B.shift_reg[103] ),
    .S(\deser_B.receiving ),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _14069_ (.A0(\deser_B.shift_reg[103] ),
    .A1(\deser_B.shift_reg[104] ),
    .S(\deser_B.receiving ),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _14070_ (.A0(\deser_B.shift_reg[104] ),
    .A1(\deser_B.shift_reg[105] ),
    .S(\deser_B.receiving ),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _14071_ (.A0(\deser_B.shift_reg[105] ),
    .A1(\deser_B.shift_reg[106] ),
    .S(\deser_B.receiving ),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _14072_ (.A0(\deser_B.shift_reg[106] ),
    .A1(\deser_B.shift_reg[107] ),
    .S(\deser_B.receiving ),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _14073_ (.A0(\deser_B.shift_reg[107] ),
    .A1(\deser_B.shift_reg[108] ),
    .S(\deser_B.receiving ),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _14074_ (.A0(\deser_B.shift_reg[108] ),
    .A1(\deser_B.shift_reg[109] ),
    .S(\deser_B.receiving ),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _14075_ (.A0(\deser_B.shift_reg[109] ),
    .A1(\deser_B.shift_reg[110] ),
    .S(\deser_B.receiving ),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _14076_ (.A0(\deser_B.shift_reg[110] ),
    .A1(\deser_B.shift_reg[111] ),
    .S(\deser_B.receiving ),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _14077_ (.A0(\deser_B.shift_reg[111] ),
    .A1(\deser_B.shift_reg[112] ),
    .S(\deser_B.receiving ),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _14078_ (.A0(\deser_B.shift_reg[112] ),
    .A1(\deser_B.shift_reg[113] ),
    .S(\deser_B.receiving ),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _14079_ (.A0(\deser_B.shift_reg[113] ),
    .A1(\deser_B.shift_reg[114] ),
    .S(\deser_B.receiving ),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _14080_ (.A0(\deser_B.shift_reg[114] ),
    .A1(\deser_B.shift_reg[115] ),
    .S(\deser_B.receiving ),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _14081_ (.A0(\deser_B.shift_reg[115] ),
    .A1(\deser_B.shift_reg[116] ),
    .S(\deser_B.receiving ),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _14082_ (.A0(\deser_B.shift_reg[116] ),
    .A1(\deser_B.shift_reg[117] ),
    .S(\deser_B.receiving ),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _14083_ (.A0(\deser_B.shift_reg[117] ),
    .A1(\deser_B.shift_reg[118] ),
    .S(\deser_B.receiving ),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _14084_ (.A0(\deser_B.shift_reg[118] ),
    .A1(\deser_B.shift_reg[119] ),
    .S(\deser_B.receiving ),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _14085_ (.A0(\deser_B.shift_reg[119] ),
    .A1(\deser_B.shift_reg[120] ),
    .S(\deser_B.receiving ),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _14086_ (.A0(\deser_B.shift_reg[120] ),
    .A1(\deser_B.shift_reg[121] ),
    .S(\deser_B.receiving ),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _14087_ (.A0(\deser_B.shift_reg[121] ),
    .A1(\deser_B.shift_reg[122] ),
    .S(\deser_B.receiving ),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _14088_ (.A0(\deser_B.shift_reg[122] ),
    .A1(\deser_B.shift_reg[123] ),
    .S(\deser_B.receiving ),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _14089_ (.A0(\deser_B.shift_reg[123] ),
    .A1(\deser_B.shift_reg[124] ),
    .S(\deser_B.receiving ),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _14090_ (.A0(\deser_B.shift_reg[124] ),
    .A1(\deser_B.shift_reg[125] ),
    .S(\deser_B.receiving ),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _14091_ (.A0(\deser_B.shift_reg[125] ),
    .A1(\deser_B.shift_reg[126] ),
    .S(\deser_B.receiving ),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _14092_ (.A0(\deser_B.shift_reg[126] ),
    .A1(\deser_B.shift_reg[127] ),
    .S(\deser_B.receiving ),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _14093_ (.A0(\deser_B.shift_reg[127] ),
    .A1(B_in_serial_data),
    .S(\deser_B.receiving ),
    .X(_00919_));
 sky130_fd_sc_hd__and3b_2 _14094_ (.A_N(\deser_A.receiving ),
    .B(A_in_serial_data),
    .C(A_in_frame_sync),
    .X(_11330_));
 sky130_fd_sc_hd__a221o_2 _14095_ (.A1(\deser_A.receiving ),
    .A2(\deser_A.shift_reg[1] ),
    .B1(\deser_A.shift_reg[0] ),
    .B2(_11304_),
    .C1(_11330_),
    .X(_00920_));
 sky130_fd_sc_hd__and3b_2 _14096_ (.A_N(\deser_B.receiving ),
    .B(B_in_serial_data),
    .C(B_in_frame_sync),
    .X(_11331_));
 sky130_fd_sc_hd__a221o_2 _14097_ (.A1(\deser_B.receiving ),
    .A2(\deser_B.shift_reg[1] ),
    .B1(\deser_B.shift_reg[0] ),
    .B2(_11305_),
    .C1(_11331_),
    .X(_00921_));
 sky130_fd_sc_hd__nand2_2 _14098_ (.A(rst_n),
    .B(_11306_),
    .Y(_11332_));
 sky130_fd_sc_hd__and2_2 _14099_ (.A(rst_n),
    .B(_00008_),
    .X(_11333_));
 sky130_fd_sc_hd__a22o_2 _14100_ (.A1(\systolic_inst.A_shift[12][0] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[56] ),
    .X(_00922_));
 sky130_fd_sc_hd__a22o_2 _14101_ (.A1(\systolic_inst.A_shift[12][1] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[57] ),
    .X(_00923_));
 sky130_fd_sc_hd__a22o_2 _14102_ (.A1(\systolic_inst.A_shift[12][2] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[58] ),
    .X(_00924_));
 sky130_fd_sc_hd__a22o_2 _14103_ (.A1(\systolic_inst.A_shift[12][3] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[59] ),
    .X(_00925_));
 sky130_fd_sc_hd__a22o_2 _14104_ (.A1(\systolic_inst.A_shift[12][4] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[60] ),
    .X(_00926_));
 sky130_fd_sc_hd__a22o_2 _14105_ (.A1(\systolic_inst.A_shift[12][5] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[61] ),
    .X(_00927_));
 sky130_fd_sc_hd__a22o_2 _14106_ (.A1(\systolic_inst.A_shift[12][6] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[62] ),
    .X(_00928_));
 sky130_fd_sc_hd__a22o_2 _14107_ (.A1(\systolic_inst.A_shift[12][7] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[63] ),
    .X(_00929_));
 sky130_fd_sc_hd__a22o_2 _14108_ (.A1(\systolic_inst.B_shift[12][0] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[96] ),
    .X(_00930_));
 sky130_fd_sc_hd__a22o_2 _14109_ (.A1(\systolic_inst.B_shift[12][1] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[97] ),
    .X(_00931_));
 sky130_fd_sc_hd__a22o_2 _14110_ (.A1(\systolic_inst.B_shift[12][2] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[98] ),
    .X(_00932_));
 sky130_fd_sc_hd__a22o_2 _14111_ (.A1(\systolic_inst.B_shift[12][3] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[99] ),
    .X(_00933_));
 sky130_fd_sc_hd__a22o_2 _14112_ (.A1(\systolic_inst.B_shift[12][4] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[100] ),
    .X(_00934_));
 sky130_fd_sc_hd__a22o_2 _14113_ (.A1(\systolic_inst.B_shift[12][5] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[101] ),
    .X(_00935_));
 sky130_fd_sc_hd__a22o_2 _14114_ (.A1(\systolic_inst.B_shift[12][6] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[102] ),
    .X(_00936_));
 sky130_fd_sc_hd__a22o_2 _14115_ (.A1(\systolic_inst.B_shift[12][7] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[103] ),
    .X(_00937_));
 sky130_fd_sc_hd__a22o_2 _14116_ (.A1(\systolic_inst.A_shift[21][0] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[88] ),
    .X(_00938_));
 sky130_fd_sc_hd__a22o_2 _14117_ (.A1(\systolic_inst.A_shift[21][1] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[89] ),
    .X(_00939_));
 sky130_fd_sc_hd__a22o_2 _14118_ (.A1(\systolic_inst.A_shift[21][2] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[90] ),
    .X(_00940_));
 sky130_fd_sc_hd__a22o_2 _14119_ (.A1(\systolic_inst.A_shift[21][3] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[91] ),
    .X(_00941_));
 sky130_fd_sc_hd__a22o_2 _14120_ (.A1(\systolic_inst.A_shift[21][4] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[92] ),
    .X(_00942_));
 sky130_fd_sc_hd__a22o_2 _14121_ (.A1(\systolic_inst.A_shift[21][5] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[93] ),
    .X(_00943_));
 sky130_fd_sc_hd__a22o_2 _14122_ (.A1(\systolic_inst.A_shift[21][6] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[94] ),
    .X(_00944_));
 sky130_fd_sc_hd__a22o_2 _14123_ (.A1(\systolic_inst.A_shift[21][7] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[95] ),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _14124_ (.A0(\systolic_inst.A_outs[15][0] ),
    .A1(\systolic_inst.A_outs[14][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _14125_ (.A0(\systolic_inst.A_outs[15][1] ),
    .A1(\systolic_inst.A_outs[14][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _14126_ (.A0(\systolic_inst.A_outs[15][2] ),
    .A1(\systolic_inst.A_outs[14][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _14127_ (.A0(\systolic_inst.A_outs[15][3] ),
    .A1(\systolic_inst.A_outs[14][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _14128_ (.A0(\systolic_inst.A_outs[15][4] ),
    .A1(\systolic_inst.A_outs[14][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _14129_ (.A0(\systolic_inst.A_outs[15][5] ),
    .A1(\systolic_inst.A_outs[14][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _14130_ (.A0(\systolic_inst.A_outs[15][6] ),
    .A1(\systolic_inst.A_outs[14][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _14131_ (.A0(\systolic_inst.A_outs[15][7] ),
    .A1(\systolic_inst.A_outs[14][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _14132_ (.A0(\systolic_inst.B_outs[14][0] ),
    .A1(\systolic_inst.B_outs[10][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _14133_ (.A0(\systolic_inst.B_outs[14][1] ),
    .A1(\systolic_inst.B_outs[10][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _14134_ (.A0(\systolic_inst.B_outs[14][2] ),
    .A1(\systolic_inst.B_outs[10][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _14135_ (.A0(\systolic_inst.B_outs[14][3] ),
    .A1(\systolic_inst.B_outs[10][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _14136_ (.A0(\systolic_inst.B_outs[14][4] ),
    .A1(\systolic_inst.B_outs[10][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _14137_ (.A0(\systolic_inst.B_outs[14][5] ),
    .A1(\systolic_inst.B_outs[10][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _14138_ (.A0(\systolic_inst.B_outs[14][6] ),
    .A1(\systolic_inst.B_outs[10][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _14139_ (.A0(\systolic_inst.B_outs[14][7] ),
    .A1(\systolic_inst.B_outs[10][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_00961_));
 sky130_fd_sc_hd__and3_2 _14140_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[15][0] ),
    .C(\systolic_inst.A_outs[15][0] ),
    .X(_11334_));
 sky130_fd_sc_hd__a21o_2 _14141_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[0] ),
    .B1(_11334_),
    .X(_00962_));
 sky130_fd_sc_hd__a22o_2 _14142_ (.A1(\systolic_inst.B_outs[15][0] ),
    .A2(\systolic_inst.A_outs[15][1] ),
    .B1(\systolic_inst.B_outs[15][1] ),
    .B2(\systolic_inst.A_outs[15][0] ),
    .X(_11335_));
 sky130_fd_sc_hd__and4_2 _14143_ (.A(\systolic_inst.B_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][0] ),
    .C(\systolic_inst.A_outs[15][1] ),
    .D(\systolic_inst.B_outs[15][1] ),
    .X(_11336_));
 sky130_fd_sc_hd__nor2_2 _14144_ (.A(_11258_),
    .B(_11336_),
    .Y(_11337_));
 sky130_fd_sc_hd__a22o_2 _14145_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[1] ),
    .B1(_11335_),
    .B2(_11337_),
    .X(_00963_));
 sky130_fd_sc_hd__and2_2 _14146_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[2] ),
    .X(_11338_));
 sky130_fd_sc_hd__a22o_2 _14147_ (.A1(\systolic_inst.A_outs[15][1] ),
    .A2(\systolic_inst.B_outs[15][1] ),
    .B1(\systolic_inst.B_outs[15][2] ),
    .B2(\systolic_inst.A_outs[15][0] ),
    .X(_11339_));
 sky130_fd_sc_hd__nand4_2 _14148_ (.A(\systolic_inst.A_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][1] ),
    .C(\systolic_inst.B_outs[15][1] ),
    .D(\systolic_inst.B_outs[15][2] ),
    .Y(_11340_));
 sky130_fd_sc_hd__and4_2 _14149_ (.A(\systolic_inst.B_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][2] ),
    .C(_11339_),
    .D(_11340_),
    .X(_11341_));
 sky130_fd_sc_hd__a22oi_2 _14150_ (.A1(\systolic_inst.B_outs[15][0] ),
    .A2(\systolic_inst.A_outs[15][2] ),
    .B1(_11339_),
    .B2(_11340_),
    .Y(_11342_));
 sky130_fd_sc_hd__nor2_2 _14151_ (.A(_11341_),
    .B(_11342_),
    .Y(_11343_));
 sky130_fd_sc_hd__or2_2 _14152_ (.A(_11336_),
    .B(_11343_),
    .X(_11344_));
 sky130_fd_sc_hd__nand2_2 _14153_ (.A(_11336_),
    .B(_11343_),
    .Y(_11345_));
 sky130_fd_sc_hd__a31o_2 _14154_ (.A1(\systolic_inst.ce_local ),
    .A2(_11344_),
    .A3(_11345_),
    .B1(_11338_),
    .X(_00964_));
 sky130_fd_sc_hd__a22o_2 _14155_ (.A1(\systolic_inst.B_outs[15][1] ),
    .A2(\systolic_inst.A_outs[15][2] ),
    .B1(\systolic_inst.B_outs[15][2] ),
    .B2(\systolic_inst.A_outs[15][1] ),
    .X(_11346_));
 sky130_fd_sc_hd__nand4_2 _14156_ (.A(\systolic_inst.A_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][1] ),
    .C(\systolic_inst.A_outs[15][2] ),
    .D(\systolic_inst.B_outs[15][2] ),
    .Y(_11347_));
 sky130_fd_sc_hd__nand2_2 _14157_ (.A(_11346_),
    .B(_11347_),
    .Y(_11348_));
 sky130_fd_sc_hd__xnor2_2 _14158_ (.A(_11340_),
    .B(_11348_),
    .Y(_11349_));
 sky130_fd_sc_hd__a22oi_2 _14159_ (.A1(\systolic_inst.A_outs[15][0] ),
    .A2(\systolic_inst.B_outs[15][3] ),
    .B1(\systolic_inst.A_outs[15][3] ),
    .B2(\systolic_inst.B_outs[15][0] ),
    .Y(_11350_));
 sky130_fd_sc_hd__and4_2 _14160_ (.A(\systolic_inst.B_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][0] ),
    .C(\systolic_inst.B_outs[15][3] ),
    .D(\systolic_inst.A_outs[15][3] ),
    .X(_11351_));
 sky130_fd_sc_hd__or2_2 _14161_ (.A(_11350_),
    .B(_11351_),
    .X(_11352_));
 sky130_fd_sc_hd__xor2_2 _14162_ (.A(_11349_),
    .B(_11352_),
    .X(_11353_));
 sky130_fd_sc_hd__nand2_2 _14163_ (.A(_11341_),
    .B(_11353_),
    .Y(_11354_));
 sky130_fd_sc_hd__xnor2_2 _14164_ (.A(_11341_),
    .B(_11353_),
    .Y(_11355_));
 sky130_fd_sc_hd__or2_2 _14165_ (.A(_11345_),
    .B(_11355_),
    .X(_11356_));
 sky130_fd_sc_hd__nand2_2 _14166_ (.A(_11345_),
    .B(_11355_),
    .Y(_11357_));
 sky130_fd_sc_hd__and2_2 _14167_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[3] ),
    .X(_11358_));
 sky130_fd_sc_hd__a31o_2 _14168_ (.A1(\systolic_inst.ce_local ),
    .A2(_11356_),
    .A3(_11357_),
    .B1(_11358_),
    .X(_00965_));
 sky130_fd_sc_hd__a22oi_2 _14169_ (.A1(\systolic_inst.A_outs[15][2] ),
    .A2(\systolic_inst.B_outs[15][2] ),
    .B1(\systolic_inst.A_outs[15][3] ),
    .B2(\systolic_inst.B_outs[15][1] ),
    .Y(_11359_));
 sky130_fd_sc_hd__and4_2 _14170_ (.A(\systolic_inst.B_outs[15][1] ),
    .B(\systolic_inst.A_outs[15][2] ),
    .C(\systolic_inst.B_outs[15][2] ),
    .D(\systolic_inst.A_outs[15][3] ),
    .X(_11360_));
 sky130_fd_sc_hd__nor2_2 _14171_ (.A(_11359_),
    .B(_11360_),
    .Y(_11361_));
 sky130_fd_sc_hd__xnor2_2 _14172_ (.A(_11351_),
    .B(_11361_),
    .Y(_11362_));
 sky130_fd_sc_hd__nor2_2 _14173_ (.A(_11347_),
    .B(_11362_),
    .Y(_11363_));
 sky130_fd_sc_hd__xnor2_2 _14174_ (.A(_11347_),
    .B(_11362_),
    .Y(_11364_));
 sky130_fd_sc_hd__and2_2 _14175_ (.A(\systolic_inst.B_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][4] ),
    .X(_11365_));
 sky130_fd_sc_hd__nand4_2 _14176_ (.A(\systolic_inst.A_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][1] ),
    .C(\systolic_inst.B_outs[15][3] ),
    .D(\systolic_inst.B_outs[15][4] ),
    .Y(_11366_));
 sky130_fd_sc_hd__a22o_2 _14177_ (.A1(\systolic_inst.A_outs[15][1] ),
    .A2(\systolic_inst.B_outs[15][3] ),
    .B1(\systolic_inst.B_outs[15][4] ),
    .B2(\systolic_inst.A_outs[15][0] ),
    .X(_11367_));
 sky130_fd_sc_hd__nand2_2 _14178_ (.A(_11366_),
    .B(_11367_),
    .Y(_11368_));
 sky130_fd_sc_hd__xnor2_2 _14179_ (.A(_11365_),
    .B(_11368_),
    .Y(_11369_));
 sky130_fd_sc_hd__and2b_2 _14180_ (.A_N(_11364_),
    .B(_11369_),
    .X(_11370_));
 sky130_fd_sc_hd__xnor2_2 _14181_ (.A(_11364_),
    .B(_11369_),
    .Y(_11371_));
 sky130_fd_sc_hd__o22ai_2 _14182_ (.A1(_11340_),
    .A2(_11348_),
    .B1(_11349_),
    .B2(_11352_),
    .Y(_11372_));
 sky130_fd_sc_hd__nand2_2 _14183_ (.A(_11371_),
    .B(_11372_),
    .Y(_11373_));
 sky130_fd_sc_hd__xnor2_2 _14184_ (.A(_11371_),
    .B(_11372_),
    .Y(_11374_));
 sky130_fd_sc_hd__a21o_2 _14185_ (.A1(_11354_),
    .A2(_11356_),
    .B1(_11374_),
    .X(_11375_));
 sky130_fd_sc_hd__a31o_2 _14186_ (.A1(_11354_),
    .A2(_11356_),
    .A3(_11374_),
    .B1(_11258_),
    .X(_11376_));
 sky130_fd_sc_hd__and2b_2 _14187_ (.A_N(_11376_),
    .B(_11375_),
    .X(_11377_));
 sky130_fd_sc_hd__a21o_2 _14188_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[4] ),
    .B1(_11377_),
    .X(_00966_));
 sky130_fd_sc_hd__a21o_2 _14189_ (.A1(_11351_),
    .A2(_11361_),
    .B1(_11363_),
    .X(_11378_));
 sky130_fd_sc_hd__a21bo_2 _14190_ (.A1(_11365_),
    .A2(_11367_),
    .B1_N(_11366_),
    .X(_11379_));
 sky130_fd_sc_hd__a22oi_2 _14191_ (.A1(\systolic_inst.B_outs[15][2] ),
    .A2(\systolic_inst.A_outs[15][3] ),
    .B1(\systolic_inst.A_outs[15][4] ),
    .B2(\systolic_inst.B_outs[15][1] ),
    .Y(_11380_));
 sky130_fd_sc_hd__and4_2 _14192_ (.A(\systolic_inst.B_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][2] ),
    .C(\systolic_inst.A_outs[15][3] ),
    .D(\systolic_inst.A_outs[15][4] ),
    .X(_11381_));
 sky130_fd_sc_hd__or2_2 _14193_ (.A(_11380_),
    .B(_11381_),
    .X(_11382_));
 sky130_fd_sc_hd__nand2b_2 _14194_ (.A_N(_11382_),
    .B(_11379_),
    .Y(_11383_));
 sky130_fd_sc_hd__xnor2_2 _14195_ (.A(_11379_),
    .B(_11382_),
    .Y(_11384_));
 sky130_fd_sc_hd__xnor2_2 _14196_ (.A(_11360_),
    .B(_11384_),
    .Y(_11385_));
 sky130_fd_sc_hd__and2_2 _14197_ (.A(\systolic_inst.A_outs[15][0] ),
    .B(\systolic_inst.B_outs[15][5] ),
    .X(_11386_));
 sky130_fd_sc_hd__nand2_2 _14198_ (.A(\systolic_inst.B_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][5] ),
    .Y(_11387_));
 sky130_fd_sc_hd__and4_2 _14199_ (.A(\systolic_inst.A_outs[15][1] ),
    .B(\systolic_inst.A_outs[15][2] ),
    .C(\systolic_inst.B_outs[15][3] ),
    .D(\systolic_inst.B_outs[15][4] ),
    .X(_11388_));
 sky130_fd_sc_hd__a22oi_2 _14200_ (.A1(\systolic_inst.A_outs[15][2] ),
    .A2(\systolic_inst.B_outs[15][3] ),
    .B1(\systolic_inst.B_outs[15][4] ),
    .B2(\systolic_inst.A_outs[15][1] ),
    .Y(_11389_));
 sky130_fd_sc_hd__or3_2 _14201_ (.A(_11387_),
    .B(_11388_),
    .C(_11389_),
    .X(_11390_));
 sky130_fd_sc_hd__o21ai_2 _14202_ (.A1(_11388_),
    .A2(_11389_),
    .B1(_11387_),
    .Y(_11391_));
 sky130_fd_sc_hd__and3_2 _14203_ (.A(_11386_),
    .B(_11390_),
    .C(_11391_),
    .X(_11392_));
 sky130_fd_sc_hd__a21oi_2 _14204_ (.A1(_11390_),
    .A2(_11391_),
    .B1(_11386_),
    .Y(_11393_));
 sky130_fd_sc_hd__or2_2 _14205_ (.A(_11392_),
    .B(_11393_),
    .X(_11394_));
 sky130_fd_sc_hd__nor2_2 _14206_ (.A(_11385_),
    .B(_11394_),
    .Y(_11395_));
 sky130_fd_sc_hd__xor2_2 _14207_ (.A(_11385_),
    .B(_11394_),
    .X(_11396_));
 sky130_fd_sc_hd__nand2_2 _14208_ (.A(_11370_),
    .B(_11396_),
    .Y(_11397_));
 sky130_fd_sc_hd__xor2_2 _14209_ (.A(_11370_),
    .B(_11396_),
    .X(_11398_));
 sky130_fd_sc_hd__nand2_2 _14210_ (.A(_11378_),
    .B(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__xnor2_2 _14211_ (.A(_11378_),
    .B(_11398_),
    .Y(_11400_));
 sky130_fd_sc_hd__a21oi_2 _14212_ (.A1(_11373_),
    .A2(_11375_),
    .B1(_11400_),
    .Y(_11401_));
 sky130_fd_sc_hd__a31o_2 _14213_ (.A1(_11373_),
    .A2(_11375_),
    .A3(_11400_),
    .B1(_11258_),
    .X(_11402_));
 sky130_fd_sc_hd__a2bb2o_2 _14214_ (.A1_N(_11402_),
    .A2_N(_11401_),
    .B1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[5] ),
    .B2(_11258_),
    .X(_00967_));
 sky130_fd_sc_hd__a21bo_2 _14215_ (.A1(_11360_),
    .A2(_11384_),
    .B1_N(_11383_),
    .X(_11403_));
 sky130_fd_sc_hd__o21bai_2 _14216_ (.A1(_11387_),
    .A2(_11389_),
    .B1_N(_11388_),
    .Y(_11404_));
 sky130_fd_sc_hd__a22oi_2 _14217_ (.A1(\systolic_inst.B_outs[15][2] ),
    .A2(\systolic_inst.A_outs[15][4] ),
    .B1(\systolic_inst.A_outs[15][5] ),
    .B2(\systolic_inst.B_outs[15][1] ),
    .Y(_11405_));
 sky130_fd_sc_hd__and4_2 _14218_ (.A(\systolic_inst.B_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][2] ),
    .C(\systolic_inst.A_outs[15][4] ),
    .D(\systolic_inst.A_outs[15][5] ),
    .X(_11406_));
 sky130_fd_sc_hd__or2_2 _14219_ (.A(_11405_),
    .B(_11406_),
    .X(_11407_));
 sky130_fd_sc_hd__and2b_2 _14220_ (.A_N(_11407_),
    .B(_11404_),
    .X(_11408_));
 sky130_fd_sc_hd__xnor2_2 _14221_ (.A(_11404_),
    .B(_11407_),
    .Y(_11409_));
 sky130_fd_sc_hd__xor2_2 _14222_ (.A(_11381_),
    .B(_11409_),
    .X(_11410_));
 sky130_fd_sc_hd__nand4_2 _14223_ (.A(\systolic_inst.A_outs[15][2] ),
    .B(\systolic_inst.B_outs[15][3] ),
    .C(\systolic_inst.A_outs[15][3] ),
    .D(\systolic_inst.B_outs[15][4] ),
    .Y(_11411_));
 sky130_fd_sc_hd__a22o_2 _14224_ (.A1(\systolic_inst.B_outs[15][3] ),
    .A2(\systolic_inst.A_outs[15][3] ),
    .B1(\systolic_inst.B_outs[15][4] ),
    .B2(\systolic_inst.A_outs[15][2] ),
    .X(_11412_));
 sky130_fd_sc_hd__nand4_2 _14225_ (.A(\systolic_inst.B_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][6] ),
    .C(_11411_),
    .D(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__a22o_2 _14226_ (.A1(\systolic_inst.B_outs[15][0] ),
    .A2(\systolic_inst.A_outs[15][6] ),
    .B1(_11411_),
    .B2(_11412_),
    .X(_11414_));
 sky130_fd_sc_hd__a22oi_2 _14227_ (.A1(\systolic_inst.A_outs[15][1] ),
    .A2(\systolic_inst.B_outs[15][5] ),
    .B1(\systolic_inst.B_outs[15][6] ),
    .B2(\systolic_inst.A_outs[15][0] ),
    .Y(_11415_));
 sky130_fd_sc_hd__nand2_2 _14228_ (.A(\systolic_inst.A_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][6] ),
    .Y(_11416_));
 sky130_fd_sc_hd__and4_2 _14229_ (.A(\systolic_inst.A_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][1] ),
    .C(\systolic_inst.B_outs[15][5] ),
    .D(\systolic_inst.B_outs[15][6] ),
    .X(_11417_));
 sky130_fd_sc_hd__nor2_2 _14230_ (.A(_11415_),
    .B(_11417_),
    .Y(_11418_));
 sky130_fd_sc_hd__nand3_2 _14231_ (.A(_11413_),
    .B(_11414_),
    .C(_11418_),
    .Y(_11419_));
 sky130_fd_sc_hd__a21o_2 _14232_ (.A1(_11413_),
    .A2(_11414_),
    .B1(_11418_),
    .X(_11420_));
 sky130_fd_sc_hd__and3_2 _14233_ (.A(_11392_),
    .B(_11419_),
    .C(_11420_),
    .X(_11421_));
 sky130_fd_sc_hd__a21oi_2 _14234_ (.A1(_11419_),
    .A2(_11420_),
    .B1(_11392_),
    .Y(_11422_));
 sky130_fd_sc_hd__or3b_2 _14235_ (.A(_11421_),
    .B(_11422_),
    .C_N(_11410_),
    .X(_11423_));
 sky130_fd_sc_hd__o21bai_2 _14236_ (.A1(_11421_),
    .A2(_11422_),
    .B1_N(_11410_),
    .Y(_11424_));
 sky130_fd_sc_hd__nand3_2 _14237_ (.A(_11395_),
    .B(_11423_),
    .C(_11424_),
    .Y(_11425_));
 sky130_fd_sc_hd__inv_2 _14238_ (.A(_11425_),
    .Y(_11426_));
 sky130_fd_sc_hd__a21o_2 _14239_ (.A1(_11423_),
    .A2(_11424_),
    .B1(_11395_),
    .X(_11427_));
 sky130_fd_sc_hd__and3_2 _14240_ (.A(_11403_),
    .B(_11425_),
    .C(_11427_),
    .X(_11428_));
 sky130_fd_sc_hd__a21oi_2 _14241_ (.A1(_11425_),
    .A2(_11427_),
    .B1(_11403_),
    .Y(_11429_));
 sky130_fd_sc_hd__a211oi_2 _14242_ (.A1(_11397_),
    .A2(_11399_),
    .B1(_11428_),
    .C1(_11429_),
    .Y(_11430_));
 sky130_fd_sc_hd__o211ai_2 _14243_ (.A1(_11428_),
    .A2(_11429_),
    .B1(_11397_),
    .C1(_11399_),
    .Y(_11431_));
 sky130_fd_sc_hd__and2b_2 _14244_ (.A_N(_11430_),
    .B(_11431_),
    .X(_11432_));
 sky130_fd_sc_hd__xor2_2 _14245_ (.A(_11401_),
    .B(_11432_),
    .X(_11433_));
 sky130_fd_sc_hd__mux2_1 _14246_ (.A0(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[6] ),
    .A1(_11433_),
    .S(\systolic_inst.ce_local ),
    .X(_00968_));
 sky130_fd_sc_hd__a21o_2 _14247_ (.A1(_11401_),
    .A2(_11431_),
    .B1(_11430_),
    .X(_11434_));
 sky130_fd_sc_hd__nor2_2 _14248_ (.A(_11426_),
    .B(_11428_),
    .Y(_11435_));
 sky130_fd_sc_hd__a21o_2 _14249_ (.A1(_11381_),
    .A2(_11409_),
    .B1(_11408_),
    .X(_11436_));
 sky130_fd_sc_hd__nand2_2 _14250_ (.A(_11411_),
    .B(_11413_),
    .Y(_11437_));
 sky130_fd_sc_hd__a22o_2 _14251_ (.A1(\systolic_inst.B_outs[15][2] ),
    .A2(\systolic_inst.A_outs[15][5] ),
    .B1(\systolic_inst.A_outs[15][6] ),
    .B2(\systolic_inst.B_outs[15][1] ),
    .X(_11438_));
 sky130_fd_sc_hd__and4_2 _14252_ (.A(\systolic_inst.B_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][2] ),
    .C(\systolic_inst.A_outs[15][5] ),
    .D(\systolic_inst.A_outs[15][6] ),
    .X(_11439_));
 sky130_fd_sc_hd__inv_2 _14253_ (.A(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__and3_2 _14254_ (.A(\systolic_inst.B_outs[15][7] ),
    .B(_11438_),
    .C(_11440_),
    .X(_11441_));
 sky130_fd_sc_hd__a21oi_2 _14255_ (.A1(_11438_),
    .A2(_11440_),
    .B1(\systolic_inst.B_outs[15][7] ),
    .Y(_11442_));
 sky130_fd_sc_hd__or2_2 _14256_ (.A(_11441_),
    .B(_11442_),
    .X(_11443_));
 sky130_fd_sc_hd__and2b_2 _14257_ (.A_N(_11443_),
    .B(_11437_),
    .X(_11444_));
 sky130_fd_sc_hd__xnor2_2 _14258_ (.A(_11437_),
    .B(_11443_),
    .Y(_11445_));
 sky130_fd_sc_hd__xnor2_2 _14259_ (.A(_11406_),
    .B(_11445_),
    .Y(_11446_));
 sky130_fd_sc_hd__nand2_2 _14260_ (.A(\systolic_inst.B_outs[15][0] ),
    .B(\systolic_inst.A_outs[15][7] ),
    .Y(_11447_));
 sky130_fd_sc_hd__and4_2 _14261_ (.A(\systolic_inst.B_outs[15][3] ),
    .B(\systolic_inst.A_outs[15][3] ),
    .C(\systolic_inst.B_outs[15][4] ),
    .D(\systolic_inst.A_outs[15][4] ),
    .X(_11448_));
 sky130_fd_sc_hd__a22oi_2 _14262_ (.A1(\systolic_inst.A_outs[15][3] ),
    .A2(\systolic_inst.B_outs[15][4] ),
    .B1(\systolic_inst.A_outs[15][4] ),
    .B2(\systolic_inst.B_outs[15][3] ),
    .Y(_11449_));
 sky130_fd_sc_hd__or2_2 _14263_ (.A(_11448_),
    .B(_11449_),
    .X(_11450_));
 sky130_fd_sc_hd__xor2_2 _14264_ (.A(_11447_),
    .B(_11450_),
    .X(_11451_));
 sky130_fd_sc_hd__nand2_2 _14265_ (.A(\systolic_inst.A_outs[15][2] ),
    .B(\systolic_inst.B_outs[15][5] ),
    .Y(_11452_));
 sky130_fd_sc_hd__and2b_2 _14266_ (.A_N(\systolic_inst.A_outs[15][0] ),
    .B(\systolic_inst.B_outs[15][7] ),
    .X(_11453_));
 sky130_fd_sc_hd__and3_2 _14267_ (.A(\systolic_inst.A_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][6] ),
    .C(_11453_),
    .X(_11454_));
 sky130_fd_sc_hd__xnor2_2 _14268_ (.A(_11416_),
    .B(_11453_),
    .Y(_11455_));
 sky130_fd_sc_hd__xnor2_2 _14269_ (.A(_11452_),
    .B(_11455_),
    .Y(_11456_));
 sky130_fd_sc_hd__nand2_2 _14270_ (.A(_11417_),
    .B(_11456_),
    .Y(_11457_));
 sky130_fd_sc_hd__or2_2 _14271_ (.A(_11417_),
    .B(_11456_),
    .X(_11458_));
 sky130_fd_sc_hd__xor2_2 _14272_ (.A(_11417_),
    .B(_11456_),
    .X(_11459_));
 sky130_fd_sc_hd__xnor2_2 _14273_ (.A(_11451_),
    .B(_11459_),
    .Y(_11460_));
 sky130_fd_sc_hd__or2_2 _14274_ (.A(_11419_),
    .B(_11460_),
    .X(_11461_));
 sky130_fd_sc_hd__and2_2 _14275_ (.A(_11419_),
    .B(_11460_),
    .X(_11462_));
 sky130_fd_sc_hd__xor2_2 _14276_ (.A(_11419_),
    .B(_11460_),
    .X(_11463_));
 sky130_fd_sc_hd__xnor2_2 _14277_ (.A(_11446_),
    .B(_11463_),
    .Y(_11464_));
 sky130_fd_sc_hd__and2b_2 _14278_ (.A_N(_11421_),
    .B(_11423_),
    .X(_11465_));
 sky130_fd_sc_hd__and2b_2 _14279_ (.A_N(_11465_),
    .B(_11464_),
    .X(_11466_));
 sky130_fd_sc_hd__xnor2_2 _14280_ (.A(_11464_),
    .B(_11465_),
    .Y(_11467_));
 sky130_fd_sc_hd__xnor2_2 _14281_ (.A(_11436_),
    .B(_11467_),
    .Y(_11468_));
 sky130_fd_sc_hd__and2_2 _14282_ (.A(_11435_),
    .B(_11468_),
    .X(_11469_));
 sky130_fd_sc_hd__nor2_2 _14283_ (.A(_11435_),
    .B(_11468_),
    .Y(_11470_));
 sky130_fd_sc_hd__nor2_2 _14284_ (.A(_11469_),
    .B(_11470_),
    .Y(_11471_));
 sky130_fd_sc_hd__a21boi_2 _14285_ (.A1(_11435_),
    .A2(_11468_),
    .B1_N(_11434_),
    .Y(_11472_));
 sky130_fd_sc_hd__o21ba_2 _14286_ (.A1(_11434_),
    .A2(_11471_),
    .B1_N(_11472_),
    .X(_11473_));
 sky130_fd_sc_hd__mux2_1 _14287_ (.A0(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[7] ),
    .A1(_11473_),
    .S(\systolic_inst.ce_local ),
    .X(_00969_));
 sky130_fd_sc_hd__a21o_2 _14288_ (.A1(_11406_),
    .A2(_11445_),
    .B1(_11444_),
    .X(_11474_));
 sky130_fd_sc_hd__or2_2 _14289_ (.A(_11439_),
    .B(_11441_),
    .X(_11475_));
 sky130_fd_sc_hd__o21bai_2 _14290_ (.A1(_11447_),
    .A2(_11449_),
    .B1_N(_11448_),
    .Y(_11476_));
 sky130_fd_sc_hd__a22o_2 _14291_ (.A1(\systolic_inst.B_outs[15][2] ),
    .A2(\systolic_inst.A_outs[15][6] ),
    .B1(\systolic_inst.A_outs[15][7] ),
    .B2(\systolic_inst.B_outs[15][1] ),
    .X(_11477_));
 sky130_fd_sc_hd__and4_2 _14292_ (.A(\systolic_inst.B_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][2] ),
    .C(\systolic_inst.A_outs[15][6] ),
    .D(\systolic_inst.A_outs[15][7] ),
    .X(_11478_));
 sky130_fd_sc_hd__nand4_2 _14293_ (.A(\systolic_inst.B_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][2] ),
    .C(\systolic_inst.A_outs[15][6] ),
    .D(\systolic_inst.A_outs[15][7] ),
    .Y(_11479_));
 sky130_fd_sc_hd__nand2_2 _14294_ (.A(_11477_),
    .B(_11479_),
    .Y(_11480_));
 sky130_fd_sc_hd__xnor2_2 _14295_ (.A(_11476_),
    .B(_11480_),
    .Y(_11481_));
 sky130_fd_sc_hd__xnor2_2 _14296_ (.A(_11475_),
    .B(_11481_),
    .Y(_11482_));
 sky130_fd_sc_hd__and4_2 _14297_ (.A(\systolic_inst.B_outs[15][3] ),
    .B(\systolic_inst.B_outs[15][4] ),
    .C(\systolic_inst.A_outs[15][4] ),
    .D(\systolic_inst.A_outs[15][5] ),
    .X(_11483_));
 sky130_fd_sc_hd__a22oi_2 _14298_ (.A1(\systolic_inst.B_outs[15][4] ),
    .A2(\systolic_inst.A_outs[15][4] ),
    .B1(\systolic_inst.A_outs[15][5] ),
    .B2(\systolic_inst.B_outs[15][3] ),
    .Y(_11484_));
 sky130_fd_sc_hd__nor2_2 _14299_ (.A(_11483_),
    .B(_11484_),
    .Y(_11485_));
 sky130_fd_sc_hd__xnor2_2 _14300_ (.A(_11447_),
    .B(_11485_),
    .Y(_11486_));
 sky130_fd_sc_hd__nand2_2 _14301_ (.A(\systolic_inst.A_outs[15][3] ),
    .B(\systolic_inst.B_outs[15][5] ),
    .Y(_11487_));
 sky130_fd_sc_hd__and2b_2 _14302_ (.A_N(\systolic_inst.A_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][7] ),
    .X(_11488_));
 sky130_fd_sc_hd__nand2_2 _14303_ (.A(\systolic_inst.A_outs[15][2] ),
    .B(\systolic_inst.B_outs[15][6] ),
    .Y(_11489_));
 sky130_fd_sc_hd__and3_2 _14304_ (.A(\systolic_inst.A_outs[15][2] ),
    .B(\systolic_inst.B_outs[15][6] ),
    .C(_11488_),
    .X(_11490_));
 sky130_fd_sc_hd__xnor2_2 _14305_ (.A(_11488_),
    .B(_11489_),
    .Y(_11491_));
 sky130_fd_sc_hd__xnor2_2 _14306_ (.A(_11487_),
    .B(_11491_),
    .Y(_11492_));
 sky130_fd_sc_hd__a31o_2 _14307_ (.A1(\systolic_inst.A_outs[15][2] ),
    .A2(\systolic_inst.B_outs[15][5] ),
    .A3(_11455_),
    .B1(_11454_),
    .X(_11493_));
 sky130_fd_sc_hd__and2_2 _14308_ (.A(_11492_),
    .B(_11493_),
    .X(_11494_));
 sky130_fd_sc_hd__xor2_2 _14309_ (.A(_11492_),
    .B(_11493_),
    .X(_11495_));
 sky130_fd_sc_hd__xnor2_2 _14310_ (.A(_11486_),
    .B(_11495_),
    .Y(_11496_));
 sky130_fd_sc_hd__a21boi_2 _14311_ (.A1(_11451_),
    .A2(_11458_),
    .B1_N(_11457_),
    .Y(_11497_));
 sky130_fd_sc_hd__nor2_2 _14312_ (.A(_11496_),
    .B(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__xnor2_2 _14313_ (.A(_11496_),
    .B(_11497_),
    .Y(_11499_));
 sky130_fd_sc_hd__nor2_2 _14314_ (.A(_11482_),
    .B(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__xor2_2 _14315_ (.A(_11482_),
    .B(_11499_),
    .X(_11501_));
 sky130_fd_sc_hd__o21a_2 _14316_ (.A1(_11446_),
    .A2(_11462_),
    .B1(_11461_),
    .X(_11502_));
 sky130_fd_sc_hd__nand2b_2 _14317_ (.A_N(_11502_),
    .B(_11501_),
    .Y(_11503_));
 sky130_fd_sc_hd__xnor2_2 _14318_ (.A(_11501_),
    .B(_11502_),
    .Y(_11504_));
 sky130_fd_sc_hd__nand2_2 _14319_ (.A(_11474_),
    .B(_11504_),
    .Y(_11505_));
 sky130_fd_sc_hd__xnor2_2 _14320_ (.A(_11474_),
    .B(_11504_),
    .Y(_11506_));
 sky130_fd_sc_hd__a21oi_2 _14321_ (.A1(_11436_),
    .A2(_11467_),
    .B1(_11466_),
    .Y(_11507_));
 sky130_fd_sc_hd__or2_2 _14322_ (.A(_11506_),
    .B(_11507_),
    .X(_11508_));
 sky130_fd_sc_hd__xor2_2 _14323_ (.A(_11506_),
    .B(_11507_),
    .X(_11509_));
 sky130_fd_sc_hd__o21ai_2 _14324_ (.A1(_11470_),
    .A2(_11472_),
    .B1(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__or3_2 _14325_ (.A(_11470_),
    .B(_11472_),
    .C(_11509_),
    .X(_11511_));
 sky130_fd_sc_hd__and3_2 _14326_ (.A(\systolic_inst.ce_local ),
    .B(_11510_),
    .C(_11511_),
    .X(_11512_));
 sky130_fd_sc_hd__a21o_2 _14327_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[8] ),
    .B1(_11512_),
    .X(_00970_));
 sky130_fd_sc_hd__nand2_2 _14328_ (.A(_11503_),
    .B(_11505_),
    .Y(_11513_));
 sky130_fd_sc_hd__a32o_2 _14329_ (.A1(_11476_),
    .A2(_11477_),
    .A3(_11479_),
    .B1(_11481_),
    .B2(_11475_),
    .X(_11514_));
 sky130_fd_sc_hd__a31o_2 _14330_ (.A1(\systolic_inst.B_outs[15][0] ),
    .A2(\systolic_inst.A_outs[15][7] ),
    .A3(_11485_),
    .B1(_11483_),
    .X(_11515_));
 sky130_fd_sc_hd__nand2_2 _14331_ (.A(\systolic_inst.B_outs[15][1] ),
    .B(\systolic_inst.B_outs[15][2] ),
    .Y(_11516_));
 sky130_fd_sc_hd__o21a_2 _14332_ (.A1(\systolic_inst.B_outs[15][1] ),
    .A2(\systolic_inst.B_outs[15][2] ),
    .B1(\systolic_inst.A_outs[15][7] ),
    .X(_11517_));
 sky130_fd_sc_hd__o21ai_2 _14333_ (.A1(\systolic_inst.B_outs[15][1] ),
    .A2(\systolic_inst.B_outs[15][2] ),
    .B1(\systolic_inst.A_outs[15][7] ),
    .Y(_11518_));
 sky130_fd_sc_hd__nand2_2 _14334_ (.A(_11516_),
    .B(_11517_),
    .Y(_11519_));
 sky130_fd_sc_hd__xnor2_2 _14335_ (.A(_11515_),
    .B(_11519_),
    .Y(_11520_));
 sky130_fd_sc_hd__and2_2 _14336_ (.A(_11478_),
    .B(_11520_),
    .X(_11521_));
 sky130_fd_sc_hd__nor2_2 _14337_ (.A(_11478_),
    .B(_11520_),
    .Y(_11522_));
 sky130_fd_sc_hd__or2_2 _14338_ (.A(_11521_),
    .B(_11522_),
    .X(_11523_));
 sky130_fd_sc_hd__a22oi_2 _14339_ (.A1(\systolic_inst.B_outs[15][4] ),
    .A2(\systolic_inst.A_outs[15][5] ),
    .B1(\systolic_inst.A_outs[15][6] ),
    .B2(\systolic_inst.B_outs[15][3] ),
    .Y(_11524_));
 sky130_fd_sc_hd__and4_2 _14340_ (.A(\systolic_inst.B_outs[15][3] ),
    .B(\systolic_inst.B_outs[15][4] ),
    .C(\systolic_inst.A_outs[15][5] ),
    .D(\systolic_inst.A_outs[15][6] ),
    .X(_11525_));
 sky130_fd_sc_hd__nor2_2 _14341_ (.A(_11524_),
    .B(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__xnor2_2 _14342_ (.A(_11447_),
    .B(_11526_),
    .Y(_11527_));
 sky130_fd_sc_hd__nand2_2 _14343_ (.A(\systolic_inst.A_outs[15][4] ),
    .B(\systolic_inst.B_outs[15][5] ),
    .Y(_11528_));
 sky130_fd_sc_hd__and2b_2 _14344_ (.A_N(\systolic_inst.A_outs[15][2] ),
    .B(\systolic_inst.B_outs[15][7] ),
    .X(_11529_));
 sky130_fd_sc_hd__nand2_2 _14345_ (.A(\systolic_inst.A_outs[15][3] ),
    .B(\systolic_inst.B_outs[15][6] ),
    .Y(_11530_));
 sky130_fd_sc_hd__and3_2 _14346_ (.A(\systolic_inst.A_outs[15][3] ),
    .B(\systolic_inst.B_outs[15][6] ),
    .C(_11529_),
    .X(_11531_));
 sky130_fd_sc_hd__xnor2_2 _14347_ (.A(_11529_),
    .B(_11530_),
    .Y(_11532_));
 sky130_fd_sc_hd__xnor2_2 _14348_ (.A(_11528_),
    .B(_11532_),
    .Y(_11533_));
 sky130_fd_sc_hd__a31o_2 _14349_ (.A1(\systolic_inst.A_outs[15][3] ),
    .A2(\systolic_inst.B_outs[15][5] ),
    .A3(_11491_),
    .B1(_11490_),
    .X(_11534_));
 sky130_fd_sc_hd__and2_2 _14350_ (.A(_11533_),
    .B(_11534_),
    .X(_11535_));
 sky130_fd_sc_hd__xor2_2 _14351_ (.A(_11533_),
    .B(_11534_),
    .X(_11536_));
 sky130_fd_sc_hd__xnor2_2 _14352_ (.A(_11527_),
    .B(_11536_),
    .Y(_11537_));
 sky130_fd_sc_hd__a21oi_2 _14353_ (.A1(_11486_),
    .A2(_11495_),
    .B1(_11494_),
    .Y(_11538_));
 sky130_fd_sc_hd__xnor2_2 _14354_ (.A(_11537_),
    .B(_11538_),
    .Y(_11539_));
 sky130_fd_sc_hd__xor2_2 _14355_ (.A(_11523_),
    .B(_11539_),
    .X(_11540_));
 sky130_fd_sc_hd__o21ai_2 _14356_ (.A1(_11498_),
    .A2(_11500_),
    .B1(_11540_),
    .Y(_11541_));
 sky130_fd_sc_hd__or3_2 _14357_ (.A(_11498_),
    .B(_11500_),
    .C(_11540_),
    .X(_11542_));
 sky130_fd_sc_hd__and2_2 _14358_ (.A(_11541_),
    .B(_11542_),
    .X(_11543_));
 sky130_fd_sc_hd__nand2_2 _14359_ (.A(_11514_),
    .B(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__xnor2_2 _14360_ (.A(_11514_),
    .B(_11543_),
    .Y(_11545_));
 sky130_fd_sc_hd__and2b_2 _14361_ (.A_N(_11545_),
    .B(_11513_),
    .X(_11546_));
 sky130_fd_sc_hd__nand2b_2 _14362_ (.A_N(_11545_),
    .B(_11513_),
    .Y(_11547_));
 sky130_fd_sc_hd__and3_2 _14363_ (.A(_11503_),
    .B(_11505_),
    .C(_11545_),
    .X(_11548_));
 sky130_fd_sc_hd__or2_2 _14364_ (.A(_11546_),
    .B(_11548_),
    .X(_11549_));
 sky130_fd_sc_hd__nand2_2 _14365_ (.A(_11508_),
    .B(_11510_),
    .Y(_11550_));
 sky130_fd_sc_hd__xnor2_2 _14366_ (.A(_11549_),
    .B(_11550_),
    .Y(_11551_));
 sky130_fd_sc_hd__mux2_1 _14367_ (.A0(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[9] ),
    .A1(_11551_),
    .S(\systolic_inst.ce_local ),
    .X(_00971_));
 sky130_fd_sc_hd__a31o_2 _14368_ (.A1(_11515_),
    .A2(_11516_),
    .A3(_11517_),
    .B1(_11521_),
    .X(_11552_));
 sky130_fd_sc_hd__o21ba_2 _14369_ (.A1(_11447_),
    .A2(_11524_),
    .B1_N(_11525_),
    .X(_11553_));
 sky130_fd_sc_hd__nor2_2 _14370_ (.A(_11518_),
    .B(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__and2_2 _14371_ (.A(_11518_),
    .B(_11553_),
    .X(_11555_));
 sky130_fd_sc_hd__or2_2 _14372_ (.A(_11554_),
    .B(_11555_),
    .X(_11556_));
 sky130_fd_sc_hd__a22o_2 _14373_ (.A1(\systolic_inst.B_outs[15][4] ),
    .A2(\systolic_inst.A_outs[15][6] ),
    .B1(\systolic_inst.A_outs[15][7] ),
    .B2(\systolic_inst.B_outs[15][3] ),
    .X(_11557_));
 sky130_fd_sc_hd__and3_2 _14374_ (.A(\systolic_inst.B_outs[15][3] ),
    .B(\systolic_inst.B_outs[15][4] ),
    .C(\systolic_inst.A_outs[15][7] ),
    .X(_11558_));
 sky130_fd_sc_hd__a21bo_2 _14375_ (.A1(\systolic_inst.A_outs[15][6] ),
    .A2(_11558_),
    .B1_N(_11557_),
    .X(_11559_));
 sky130_fd_sc_hd__xor2_2 _14376_ (.A(_11447_),
    .B(_11559_),
    .X(_11560_));
 sky130_fd_sc_hd__nand2_2 _14377_ (.A(\systolic_inst.B_outs[15][5] ),
    .B(\systolic_inst.A_outs[15][5] ),
    .Y(_11561_));
 sky130_fd_sc_hd__and4b_2 _14378_ (.A_N(\systolic_inst.A_outs[15][3] ),
    .B(\systolic_inst.A_outs[15][4] ),
    .C(\systolic_inst.B_outs[15][6] ),
    .D(\systolic_inst.B_outs[15][7] ),
    .X(_11562_));
 sky130_fd_sc_hd__o2bb2a_2 _14379_ (.A1_N(\systolic_inst.A_outs[15][4] ),
    .A2_N(\systolic_inst.B_outs[15][6] ),
    .B1(_11273_),
    .B2(\systolic_inst.A_outs[15][3] ),
    .X(_11563_));
 sky130_fd_sc_hd__nor2_2 _14380_ (.A(_11562_),
    .B(_11563_),
    .Y(_11564_));
 sky130_fd_sc_hd__xnor2_2 _14381_ (.A(_11561_),
    .B(_11564_),
    .Y(_11565_));
 sky130_fd_sc_hd__a31oi_2 _14382_ (.A1(\systolic_inst.A_outs[15][4] ),
    .A2(\systolic_inst.B_outs[15][5] ),
    .A3(_11532_),
    .B1(_11531_),
    .Y(_11566_));
 sky130_fd_sc_hd__nand2b_2 _14383_ (.A_N(_11566_),
    .B(_11565_),
    .Y(_11567_));
 sky130_fd_sc_hd__xnor2_2 _14384_ (.A(_11565_),
    .B(_11566_),
    .Y(_11568_));
 sky130_fd_sc_hd__xnor2_2 _14385_ (.A(_11560_),
    .B(_11568_),
    .Y(_11569_));
 sky130_fd_sc_hd__a21o_2 _14386_ (.A1(_11527_),
    .A2(_11536_),
    .B1(_11535_),
    .X(_11570_));
 sky130_fd_sc_hd__and2b_2 _14387_ (.A_N(_11569_),
    .B(_11570_),
    .X(_11571_));
 sky130_fd_sc_hd__xor2_2 _14388_ (.A(_11569_),
    .B(_11570_),
    .X(_11572_));
 sky130_fd_sc_hd__xor2_2 _14389_ (.A(_11556_),
    .B(_11572_),
    .X(_11573_));
 sky130_fd_sc_hd__o32a_2 _14390_ (.A1(_11521_),
    .A2(_11522_),
    .A3(_11539_),
    .B1(_11538_),
    .B2(_11537_),
    .X(_11574_));
 sky130_fd_sc_hd__nand2b_2 _14391_ (.A_N(_11574_),
    .B(_11573_),
    .Y(_11575_));
 sky130_fd_sc_hd__nand2b_2 _14392_ (.A_N(_11573_),
    .B(_11574_),
    .Y(_11576_));
 sky130_fd_sc_hd__nand2_2 _14393_ (.A(_11575_),
    .B(_11576_),
    .Y(_11577_));
 sky130_fd_sc_hd__nand2b_2 _14394_ (.A_N(_11577_),
    .B(_11552_),
    .Y(_11578_));
 sky130_fd_sc_hd__xor2_2 _14395_ (.A(_11552_),
    .B(_11577_),
    .X(_11579_));
 sky130_fd_sc_hd__a21oi_2 _14396_ (.A1(_11541_),
    .A2(_11544_),
    .B1(_11579_),
    .Y(_11580_));
 sky130_fd_sc_hd__and3_2 _14397_ (.A(_11541_),
    .B(_11544_),
    .C(_11579_),
    .X(_11581_));
 sky130_fd_sc_hd__a31o_2 _14398_ (.A1(_11508_),
    .A2(_11510_),
    .A3(_11547_),
    .B1(_11548_),
    .X(_11582_));
 sky130_fd_sc_hd__o21a_2 _14399_ (.A1(_11580_),
    .A2(_11581_),
    .B1(_11582_),
    .X(_11583_));
 sky130_fd_sc_hd__nor3_2 _14400_ (.A(_11580_),
    .B(_11581_),
    .C(_11582_),
    .Y(_11584_));
 sky130_fd_sc_hd__nor2_2 _14401_ (.A(_11583_),
    .B(_11584_),
    .Y(_11585_));
 sky130_fd_sc_hd__mux2_1 _14402_ (.A0(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[10] ),
    .A1(_11585_),
    .S(\systolic_inst.ce_local ),
    .X(_00972_));
 sky130_fd_sc_hd__or2_2 _14403_ (.A(_11580_),
    .B(_11584_),
    .X(_11586_));
 sky130_fd_sc_hd__o2bb2a_2 _14404_ (.A1_N(\systolic_inst.A_outs[15][6] ),
    .A2_N(_11558_),
    .B1(_11559_),
    .B2(_11447_),
    .X(_11587_));
 sky130_fd_sc_hd__nor2_2 _14405_ (.A(_11518_),
    .B(_11587_),
    .Y(_11588_));
 sky130_fd_sc_hd__and2_2 _14406_ (.A(_11518_),
    .B(_11587_),
    .X(_11589_));
 sky130_fd_sc_hd__or2_2 _14407_ (.A(_11588_),
    .B(_11589_),
    .X(_11590_));
 sky130_fd_sc_hd__or2_2 _14408_ (.A(\systolic_inst.B_outs[15][3] ),
    .B(\systolic_inst.B_outs[15][4] ),
    .X(_11591_));
 sky130_fd_sc_hd__and3b_2 _14409_ (.A_N(_11558_),
    .B(_11591_),
    .C(\systolic_inst.A_outs[15][7] ),
    .X(_11592_));
 sky130_fd_sc_hd__xnor2_2 _14410_ (.A(_11447_),
    .B(_11592_),
    .Y(_11593_));
 sky130_fd_sc_hd__nand2_2 _14411_ (.A(\systolic_inst.B_outs[15][5] ),
    .B(\systolic_inst.A_outs[15][6] ),
    .Y(_11594_));
 sky130_fd_sc_hd__and4b_2 _14412_ (.A_N(\systolic_inst.A_outs[15][4] ),
    .B(\systolic_inst.A_outs[15][5] ),
    .C(\systolic_inst.B_outs[15][6] ),
    .D(\systolic_inst.B_outs[15][7] ),
    .X(_11595_));
 sky130_fd_sc_hd__o2bb2a_2 _14413_ (.A1_N(\systolic_inst.A_outs[15][5] ),
    .A2_N(\systolic_inst.B_outs[15][6] ),
    .B1(_11273_),
    .B2(\systolic_inst.A_outs[15][4] ),
    .X(_11596_));
 sky130_fd_sc_hd__or2_2 _14414_ (.A(_11595_),
    .B(_11596_),
    .X(_11597_));
 sky130_fd_sc_hd__xor2_2 _14415_ (.A(_11594_),
    .B(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__o21ba_2 _14416_ (.A1(_11561_),
    .A2(_11563_),
    .B1_N(_11562_),
    .X(_11599_));
 sky130_fd_sc_hd__nand2b_2 _14417_ (.A_N(_11599_),
    .B(_11598_),
    .Y(_11600_));
 sky130_fd_sc_hd__xnor2_2 _14418_ (.A(_11598_),
    .B(_11599_),
    .Y(_11601_));
 sky130_fd_sc_hd__nand2_2 _14419_ (.A(_11593_),
    .B(_11601_),
    .Y(_11602_));
 sky130_fd_sc_hd__or2_2 _14420_ (.A(_11593_),
    .B(_11601_),
    .X(_11603_));
 sky130_fd_sc_hd__nand2_2 _14421_ (.A(_11602_),
    .B(_11603_),
    .Y(_11604_));
 sky130_fd_sc_hd__a21bo_2 _14422_ (.A1(_11560_),
    .A2(_11568_),
    .B1_N(_11567_),
    .X(_11605_));
 sky130_fd_sc_hd__nand2b_2 _14423_ (.A_N(_11604_),
    .B(_11605_),
    .Y(_11606_));
 sky130_fd_sc_hd__xor2_2 _14424_ (.A(_11604_),
    .B(_11605_),
    .X(_11607_));
 sky130_fd_sc_hd__xor2_2 _14425_ (.A(_11590_),
    .B(_11607_),
    .X(_11608_));
 sky130_fd_sc_hd__o21ba_2 _14426_ (.A1(_11556_),
    .A2(_11572_),
    .B1_N(_11571_),
    .X(_11609_));
 sky130_fd_sc_hd__and2b_2 _14427_ (.A_N(_11609_),
    .B(_11608_),
    .X(_11610_));
 sky130_fd_sc_hd__xnor2_2 _14428_ (.A(_11608_),
    .B(_11609_),
    .Y(_11611_));
 sky130_fd_sc_hd__xnor2_2 _14429_ (.A(_11554_),
    .B(_11611_),
    .Y(_11612_));
 sky130_fd_sc_hd__a21oi_2 _14430_ (.A1(_11575_),
    .A2(_11578_),
    .B1(_11612_),
    .Y(_11613_));
 sky130_fd_sc_hd__and3_2 _14431_ (.A(_11575_),
    .B(_11578_),
    .C(_11612_),
    .X(_11614_));
 sky130_fd_sc_hd__inv_2 _14432_ (.A(_11614_),
    .Y(_11615_));
 sky130_fd_sc_hd__or2_2 _14433_ (.A(_11613_),
    .B(_11614_),
    .X(_11616_));
 sky130_fd_sc_hd__xnor2_2 _14434_ (.A(_11586_),
    .B(_11616_),
    .Y(_11617_));
 sky130_fd_sc_hd__mux2_1 _14435_ (.A0(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[11] ),
    .A1(_11617_),
    .S(\systolic_inst.ce_local ),
    .X(_00973_));
 sky130_fd_sc_hd__a31o_2 _14436_ (.A1(\systolic_inst.B_outs[15][0] ),
    .A2(\systolic_inst.A_outs[15][7] ),
    .A3(_11591_),
    .B1(_11558_),
    .X(_11618_));
 sky130_fd_sc_hd__or2_2 _14437_ (.A(_11517_),
    .B(_11618_),
    .X(_11619_));
 sky130_fd_sc_hd__and2_2 _14438_ (.A(_11517_),
    .B(_11618_),
    .X(_11620_));
 sky130_fd_sc_hd__inv_2 _14439_ (.A(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__nand2_2 _14440_ (.A(_11619_),
    .B(_11621_),
    .Y(_11622_));
 sky130_fd_sc_hd__o2bb2a_2 _14441_ (.A1_N(\systolic_inst.B_outs[15][6] ),
    .A2_N(\systolic_inst.A_outs[15][6] ),
    .B1(_11273_),
    .B2(\systolic_inst.A_outs[15][5] ),
    .X(_11623_));
 sky130_fd_sc_hd__and4b_2 _14442_ (.A_N(\systolic_inst.A_outs[15][5] ),
    .B(\systolic_inst.B_outs[15][6] ),
    .C(\systolic_inst.A_outs[15][6] ),
    .D(\systolic_inst.B_outs[15][7] ),
    .X(_11624_));
 sky130_fd_sc_hd__nor2_2 _14443_ (.A(_11623_),
    .B(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__nand2_2 _14444_ (.A(\systolic_inst.B_outs[15][5] ),
    .B(\systolic_inst.A_outs[15][7] ),
    .Y(_11626_));
 sky130_fd_sc_hd__xnor2_2 _14445_ (.A(_11625_),
    .B(_11626_),
    .Y(_11627_));
 sky130_fd_sc_hd__o21ba_2 _14446_ (.A1(_11594_),
    .A2(_11596_),
    .B1_N(_11595_),
    .X(_11628_));
 sky130_fd_sc_hd__nand2b_2 _14447_ (.A_N(_11628_),
    .B(_11627_),
    .Y(_11629_));
 sky130_fd_sc_hd__xnor2_2 _14448_ (.A(_11627_),
    .B(_11628_),
    .Y(_11630_));
 sky130_fd_sc_hd__xnor2_2 _14449_ (.A(_11593_),
    .B(_11630_),
    .Y(_11631_));
 sky130_fd_sc_hd__a21o_2 _14450_ (.A1(_11600_),
    .A2(_11602_),
    .B1(_11631_),
    .X(_11632_));
 sky130_fd_sc_hd__nand3_2 _14451_ (.A(_11600_),
    .B(_11602_),
    .C(_11631_),
    .Y(_11633_));
 sky130_fd_sc_hd__nand2_2 _14452_ (.A(_11632_),
    .B(_11633_),
    .Y(_11634_));
 sky130_fd_sc_hd__xor2_2 _14453_ (.A(_11622_),
    .B(_11634_),
    .X(_11635_));
 sky130_fd_sc_hd__o21a_2 _14454_ (.A1(_11590_),
    .A2(_11607_),
    .B1(_11606_),
    .X(_11636_));
 sky130_fd_sc_hd__nand2b_2 _14455_ (.A_N(_11636_),
    .B(_11635_),
    .Y(_11637_));
 sky130_fd_sc_hd__xnor2_2 _14456_ (.A(_11635_),
    .B(_11636_),
    .Y(_11638_));
 sky130_fd_sc_hd__nand2_2 _14457_ (.A(_11588_),
    .B(_11638_),
    .Y(_11639_));
 sky130_fd_sc_hd__or2_2 _14458_ (.A(_11588_),
    .B(_11638_),
    .X(_11640_));
 sky130_fd_sc_hd__nand2_2 _14459_ (.A(_11639_),
    .B(_11640_),
    .Y(_11641_));
 sky130_fd_sc_hd__a21oi_2 _14460_ (.A1(_11554_),
    .A2(_11611_),
    .B1(_11610_),
    .Y(_11642_));
 sky130_fd_sc_hd__nor2_2 _14461_ (.A(_11641_),
    .B(_11642_),
    .Y(_11643_));
 sky130_fd_sc_hd__and2_2 _14462_ (.A(_11641_),
    .B(_11642_),
    .X(_11644_));
 sky130_fd_sc_hd__nor2_2 _14463_ (.A(_11643_),
    .B(_11644_),
    .Y(_11645_));
 sky130_fd_sc_hd__o31a_2 _14464_ (.A1(_11580_),
    .A2(_11584_),
    .A3(_11613_),
    .B1(_11615_),
    .X(_11646_));
 sky130_fd_sc_hd__and2_2 _14465_ (.A(_11645_),
    .B(_11646_),
    .X(_11647_));
 sky130_fd_sc_hd__nor2_2 _14466_ (.A(_11645_),
    .B(_11646_),
    .Y(_11648_));
 sky130_fd_sc_hd__nor2_2 _14467_ (.A(_11647_),
    .B(_11648_),
    .Y(_11649_));
 sky130_fd_sc_hd__mux2_1 _14468_ (.A0(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[12] ),
    .A1(_11649_),
    .S(\systolic_inst.ce_local ),
    .X(_00974_));
 sky130_fd_sc_hd__nand2_2 _14469_ (.A(\systolic_inst.B_outs[15][6] ),
    .B(\systolic_inst.A_outs[15][7] ),
    .Y(_11650_));
 sky130_fd_sc_hd__or2_2 _14470_ (.A(\systolic_inst.A_outs[15][6] ),
    .B(_11273_),
    .X(_11651_));
 sky130_fd_sc_hd__and2_2 _14471_ (.A(_11650_),
    .B(_11651_),
    .X(_11652_));
 sky130_fd_sc_hd__nor2_2 _14472_ (.A(_11650_),
    .B(_11651_),
    .Y(_11653_));
 sky130_fd_sc_hd__nor2_2 _14473_ (.A(_11652_),
    .B(_11653_),
    .Y(_11654_));
 sky130_fd_sc_hd__xnor2_2 _14474_ (.A(_11626_),
    .B(_11654_),
    .Y(_11655_));
 sky130_fd_sc_hd__o21ba_2 _14475_ (.A1(_11623_),
    .A2(_11626_),
    .B1_N(_11624_),
    .X(_11656_));
 sky130_fd_sc_hd__nand2b_2 _14476_ (.A_N(_11656_),
    .B(_11655_),
    .Y(_11657_));
 sky130_fd_sc_hd__xnor2_2 _14477_ (.A(_11655_),
    .B(_11656_),
    .Y(_11658_));
 sky130_fd_sc_hd__nand2_2 _14478_ (.A(_11593_),
    .B(_11658_),
    .Y(_11659_));
 sky130_fd_sc_hd__or2_2 _14479_ (.A(_11593_),
    .B(_11658_),
    .X(_11660_));
 sky130_fd_sc_hd__nand2_2 _14480_ (.A(_11659_),
    .B(_11660_),
    .Y(_11661_));
 sky130_fd_sc_hd__a21bo_2 _14481_ (.A1(_11593_),
    .A2(_11630_),
    .B1_N(_11629_),
    .X(_11662_));
 sky130_fd_sc_hd__and2b_2 _14482_ (.A_N(_11661_),
    .B(_11662_),
    .X(_11663_));
 sky130_fd_sc_hd__xor2_2 _14483_ (.A(_11661_),
    .B(_11662_),
    .X(_11664_));
 sky130_fd_sc_hd__xor2_2 _14484_ (.A(_11622_),
    .B(_11664_),
    .X(_11665_));
 sky130_fd_sc_hd__o21a_2 _14485_ (.A1(_11622_),
    .A2(_11634_),
    .B1(_11632_),
    .X(_11666_));
 sky130_fd_sc_hd__and2b_2 _14486_ (.A_N(_11666_),
    .B(_11665_),
    .X(_11667_));
 sky130_fd_sc_hd__and2b_2 _14487_ (.A_N(_11665_),
    .B(_11666_),
    .X(_11668_));
 sky130_fd_sc_hd__nor2_2 _14488_ (.A(_11667_),
    .B(_11668_),
    .Y(_11669_));
 sky130_fd_sc_hd__xnor2_2 _14489_ (.A(_11620_),
    .B(_11669_),
    .Y(_11670_));
 sky130_fd_sc_hd__nand3_2 _14490_ (.A(_11637_),
    .B(_11639_),
    .C(_11670_),
    .Y(_11671_));
 sky130_fd_sc_hd__a21o_2 _14491_ (.A1(_11637_),
    .A2(_11639_),
    .B1(_11670_),
    .X(_11672_));
 sky130_fd_sc_hd__and2_2 _14492_ (.A(_11671_),
    .B(_11672_),
    .X(_11673_));
 sky130_fd_sc_hd__nor2_2 _14493_ (.A(_11643_),
    .B(_11647_),
    .Y(_11674_));
 sky130_fd_sc_hd__xnor2_2 _14494_ (.A(_11673_),
    .B(_11674_),
    .Y(_11675_));
 sky130_fd_sc_hd__mux2_1 _14495_ (.A0(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[13] ),
    .A1(_11675_),
    .S(\systolic_inst.ce_local ),
    .X(_00975_));
 sky130_fd_sc_hd__a31o_2 _14496_ (.A1(\systolic_inst.B_outs[15][5] ),
    .A2(\systolic_inst.A_outs[15][7] ),
    .A3(_11654_),
    .B1(_11653_),
    .X(_11676_));
 sky130_fd_sc_hd__nand3_2 _14497_ (.A(\systolic_inst.B_outs[15][5] ),
    .B(\systolic_inst.B_outs[15][6] ),
    .C(\systolic_inst.A_outs[15][7] ),
    .Y(_11677_));
 sky130_fd_sc_hd__o211a_2 _14498_ (.A1(_11273_),
    .A2(\systolic_inst.A_outs[15][7] ),
    .B1(_11626_),
    .C1(_11650_),
    .X(_11678_));
 sky130_fd_sc_hd__a21oi_2 _14499_ (.A1(_11676_),
    .A2(_11677_),
    .B1(_11678_),
    .Y(_11679_));
 sky130_fd_sc_hd__or2_2 _14500_ (.A(_11593_),
    .B(_11679_),
    .X(_11680_));
 sky130_fd_sc_hd__nand2_2 _14501_ (.A(_11593_),
    .B(_11679_),
    .Y(_11681_));
 sky130_fd_sc_hd__nand2_2 _14502_ (.A(_11680_),
    .B(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__a21oi_2 _14503_ (.A1(_11657_),
    .A2(_11659_),
    .B1(_11682_),
    .Y(_11683_));
 sky130_fd_sc_hd__and3_2 _14504_ (.A(_11657_),
    .B(_11659_),
    .C(_11682_),
    .X(_11684_));
 sky130_fd_sc_hd__nor2_2 _14505_ (.A(_11683_),
    .B(_11684_),
    .Y(_11685_));
 sky130_fd_sc_hd__xnor2_2 _14506_ (.A(_11622_),
    .B(_11685_),
    .Y(_11686_));
 sky130_fd_sc_hd__o21ba_2 _14507_ (.A1(_11622_),
    .A2(_11664_),
    .B1_N(_11663_),
    .X(_11687_));
 sky130_fd_sc_hd__and2b_2 _14508_ (.A_N(_11687_),
    .B(_11686_),
    .X(_11688_));
 sky130_fd_sc_hd__xnor2_2 _14509_ (.A(_11686_),
    .B(_11687_),
    .Y(_11689_));
 sky130_fd_sc_hd__xnor2_2 _14510_ (.A(_11620_),
    .B(_11689_),
    .Y(_11690_));
 sky130_fd_sc_hd__a21oi_2 _14511_ (.A1(_11620_),
    .A2(_11669_),
    .B1(_11667_),
    .Y(_11691_));
 sky130_fd_sc_hd__nor2_2 _14512_ (.A(_11690_),
    .B(_11691_),
    .Y(_11692_));
 sky130_fd_sc_hd__or2_2 _14513_ (.A(_11690_),
    .B(_11691_),
    .X(_11693_));
 sky130_fd_sc_hd__and2_2 _14514_ (.A(_11690_),
    .B(_11691_),
    .X(_11694_));
 sky130_fd_sc_hd__nor2_2 _14515_ (.A(_11692_),
    .B(_11694_),
    .Y(_11695_));
 sky130_fd_sc_hd__a21bo_2 _14516_ (.A1(_11643_),
    .A2(_11671_),
    .B1_N(_11672_),
    .X(_11696_));
 sky130_fd_sc_hd__a21oi_2 _14517_ (.A1(_11647_),
    .A2(_11673_),
    .B1(_11696_),
    .Y(_11697_));
 sky130_fd_sc_hd__xnor2_2 _14518_ (.A(_11695_),
    .B(_11697_),
    .Y(_11698_));
 sky130_fd_sc_hd__mux2_1 _14519_ (.A0(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[14] ),
    .A1(_11698_),
    .S(\systolic_inst.ce_local ),
    .X(_00976_));
 sky130_fd_sc_hd__a21o_2 _14520_ (.A1(_11620_),
    .A2(_11689_),
    .B1(_11688_),
    .X(_11699_));
 sky130_fd_sc_hd__o21ba_2 _14521_ (.A1(_11622_),
    .A2(_11684_),
    .B1_N(_11683_),
    .X(_11700_));
 sky130_fd_sc_hd__xnor2_2 _14522_ (.A(_11619_),
    .B(_11680_),
    .Y(_11701_));
 sky130_fd_sc_hd__xnor2_2 _14523_ (.A(_11700_),
    .B(_11701_),
    .Y(_11702_));
 sky130_fd_sc_hd__xnor2_2 _14524_ (.A(_11699_),
    .B(_11702_),
    .Y(_11703_));
 sky130_fd_sc_hd__o211a_2 _14525_ (.A1(_11694_),
    .A2(_11697_),
    .B1(\systolic_inst.ce_local ),
    .C1(_11693_),
    .X(_11704_));
 sky130_fd_sc_hd__a22o_2 _14526_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B1(_11703_),
    .B2(_11704_),
    .X(_00977_));
 sky130_fd_sc_hd__a21o_2 _14527_ (.A1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[15][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_11705_));
 sky130_fd_sc_hd__a21oi_2 _14528_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[15][0] ),
    .Y(_11706_));
 sky130_fd_sc_hd__a21oi_2 _14529_ (.A1(\systolic_inst.ce_local ),
    .A2(_11705_),
    .B1(_11706_),
    .Y(_00978_));
 sky130_fd_sc_hd__and2_2 _14530_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[15][1] ),
    .X(_11707_));
 sky130_fd_sc_hd__nand2_2 _14531_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[15][1] ),
    .Y(_11708_));
 sky130_fd_sc_hd__or2_2 _14532_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[15][1] ),
    .X(_11709_));
 sky130_fd_sc_hd__and4_2 _14533_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[15][0] ),
    .C(_11708_),
    .D(_11709_),
    .X(_11710_));
 sky130_fd_sc_hd__inv_2 _14534_ (.A(_11710_),
    .Y(_11711_));
 sky130_fd_sc_hd__nor2_2 _14535_ (.A(_11258_),
    .B(\systolic_inst.load_acc ),
    .Y(_11712_));
 sky130_fd_sc_hd__or2_2 _14536_ (.A(_11258_),
    .B(\systolic_inst.load_acc ),
    .X(_11713_));
 sky130_fd_sc_hd__a22o_2 _14537_ (.A1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[15][0] ),
    .B1(_11708_),
    .B2(_11709_),
    .X(_11714_));
 sky130_fd_sc_hd__a32o_2 _14538_ (.A1(_11711_),
    .A2(_11712_),
    .A3(_11714_),
    .B1(\systolic_inst.acc_wires[15][1] ),
    .B2(_11258_),
    .X(_00979_));
 sky130_fd_sc_hd__nand2_2 _14539_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[15][2] ),
    .Y(_11715_));
 sky130_fd_sc_hd__or2_2 _14540_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[15][2] ),
    .X(_11716_));
 sky130_fd_sc_hd__a31o_2 _14541_ (.A1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[15][0] ),
    .A3(_11709_),
    .B1(_11707_),
    .X(_11717_));
 sky130_fd_sc_hd__a21o_2 _14542_ (.A1(_11715_),
    .A2(_11716_),
    .B1(_11717_),
    .X(_11718_));
 sky130_fd_sc_hd__and3_2 _14543_ (.A(_11715_),
    .B(_11716_),
    .C(_11717_),
    .X(_11719_));
 sky130_fd_sc_hd__inv_2 _14544_ (.A(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__a32o_2 _14545_ (.A1(_11712_),
    .A2(_11718_),
    .A3(_11720_),
    .B1(\systolic_inst.acc_wires[15][2] ),
    .B2(_11258_),
    .X(_00980_));
 sky130_fd_sc_hd__nand2_2 _14546_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[15][3] ),
    .Y(_11721_));
 sky130_fd_sc_hd__or2_2 _14547_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[15][3] ),
    .X(_11722_));
 sky130_fd_sc_hd__a21bo_2 _14548_ (.A1(_11716_),
    .A2(_11717_),
    .B1_N(_11715_),
    .X(_11723_));
 sky130_fd_sc_hd__a21o_2 _14549_ (.A1(_11721_),
    .A2(_11722_),
    .B1(_11723_),
    .X(_11724_));
 sky130_fd_sc_hd__and3_2 _14550_ (.A(_11721_),
    .B(_11722_),
    .C(_11723_),
    .X(_11725_));
 sky130_fd_sc_hd__inv_2 _14551_ (.A(_11725_),
    .Y(_11726_));
 sky130_fd_sc_hd__a32o_2 _14552_ (.A1(_11712_),
    .A2(_11724_),
    .A3(_11726_),
    .B1(\systolic_inst.acc_wires[15][3] ),
    .B2(_11258_),
    .X(_00981_));
 sky130_fd_sc_hd__nand2_2 _14553_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[15][4] ),
    .Y(_11727_));
 sky130_fd_sc_hd__or2_2 _14554_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[15][4] ),
    .X(_11728_));
 sky130_fd_sc_hd__a21bo_2 _14555_ (.A1(_11722_),
    .A2(_11723_),
    .B1_N(_11721_),
    .X(_11729_));
 sky130_fd_sc_hd__a21o_2 _14556_ (.A1(_11727_),
    .A2(_11728_),
    .B1(_11729_),
    .X(_11730_));
 sky130_fd_sc_hd__and3_2 _14557_ (.A(_11727_),
    .B(_11728_),
    .C(_11729_),
    .X(_11731_));
 sky130_fd_sc_hd__inv_2 _14558_ (.A(_11731_),
    .Y(_11732_));
 sky130_fd_sc_hd__a32o_2 _14559_ (.A1(_11712_),
    .A2(_11730_),
    .A3(_11732_),
    .B1(\systolic_inst.acc_wires[15][4] ),
    .B2(_11258_),
    .X(_00982_));
 sky130_fd_sc_hd__nand2_2 _14560_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[15][5] ),
    .Y(_11733_));
 sky130_fd_sc_hd__or2_2 _14561_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[15][5] ),
    .X(_11734_));
 sky130_fd_sc_hd__a21bo_2 _14562_ (.A1(_11728_),
    .A2(_11729_),
    .B1_N(_11727_),
    .X(_11735_));
 sky130_fd_sc_hd__a21o_2 _14563_ (.A1(_11733_),
    .A2(_11734_),
    .B1(_11735_),
    .X(_11736_));
 sky130_fd_sc_hd__and3_2 _14564_ (.A(_11733_),
    .B(_11734_),
    .C(_11735_),
    .X(_11737_));
 sky130_fd_sc_hd__inv_2 _14565_ (.A(_11737_),
    .Y(_11738_));
 sky130_fd_sc_hd__a32o_2 _14566_ (.A1(_11712_),
    .A2(_11736_),
    .A3(_11738_),
    .B1(\systolic_inst.acc_wires[15][5] ),
    .B2(_11258_),
    .X(_00983_));
 sky130_fd_sc_hd__nand2_2 _14567_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[15][6] ),
    .Y(_11739_));
 sky130_fd_sc_hd__or2_2 _14568_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[15][6] ),
    .X(_11740_));
 sky130_fd_sc_hd__a21bo_2 _14569_ (.A1(_11734_),
    .A2(_11735_),
    .B1_N(_11733_),
    .X(_11741_));
 sky130_fd_sc_hd__a21o_2 _14570_ (.A1(_11739_),
    .A2(_11740_),
    .B1(_11741_),
    .X(_11742_));
 sky130_fd_sc_hd__and3_2 _14571_ (.A(_11739_),
    .B(_11740_),
    .C(_11741_),
    .X(_11743_));
 sky130_fd_sc_hd__inv_2 _14572_ (.A(_11743_),
    .Y(_11744_));
 sky130_fd_sc_hd__a32o_2 _14573_ (.A1(_11712_),
    .A2(_11742_),
    .A3(_11744_),
    .B1(\systolic_inst.acc_wires[15][6] ),
    .B2(_11258_),
    .X(_00984_));
 sky130_fd_sc_hd__nand2_2 _14574_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[15][7] ),
    .Y(_11745_));
 sky130_fd_sc_hd__or2_2 _14575_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[15][7] ),
    .X(_11746_));
 sky130_fd_sc_hd__a21bo_2 _14576_ (.A1(_11740_),
    .A2(_11741_),
    .B1_N(_11739_),
    .X(_11747_));
 sky130_fd_sc_hd__a21o_2 _14577_ (.A1(_11745_),
    .A2(_11746_),
    .B1(_11747_),
    .X(_11748_));
 sky130_fd_sc_hd__nand3_2 _14578_ (.A(_11745_),
    .B(_11746_),
    .C(_11747_),
    .Y(_11749_));
 sky130_fd_sc_hd__a32o_2 _14579_ (.A1(_11712_),
    .A2(_11748_),
    .A3(_11749_),
    .B1(\systolic_inst.acc_wires[15][7] ),
    .B2(_11258_),
    .X(_00985_));
 sky130_fd_sc_hd__a21bo_2 _14580_ (.A1(_11746_),
    .A2(_11747_),
    .B1_N(_11745_),
    .X(_11750_));
 sky130_fd_sc_hd__xor2_2 _14581_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[15][8] ),
    .X(_11751_));
 sky130_fd_sc_hd__and2_2 _14582_ (.A(_11750_),
    .B(_11751_),
    .X(_11752_));
 sky130_fd_sc_hd__o21ai_2 _14583_ (.A1(_11750_),
    .A2(_11751_),
    .B1(_11712_),
    .Y(_11753_));
 sky130_fd_sc_hd__a2bb2o_2 _14584_ (.A1_N(_11753_),
    .A2_N(_11752_),
    .B1(\systolic_inst.acc_wires[15][8] ),
    .B2(_11258_),
    .X(_00986_));
 sky130_fd_sc_hd__xor2_2 _14585_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[15][9] ),
    .X(_11754_));
 sky130_fd_sc_hd__a211o_2 _14586_ (.A1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[15][8] ),
    .B1(_11752_),
    .C1(_11754_),
    .X(_11755_));
 sky130_fd_sc_hd__nand2_2 _14587_ (.A(_11751_),
    .B(_11754_),
    .Y(_11756_));
 sky130_fd_sc_hd__nand2_2 _14588_ (.A(_11752_),
    .B(_11754_),
    .Y(_11757_));
 sky130_fd_sc_hd__and3_2 _14589_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[15][8] ),
    .C(_11754_),
    .X(_11758_));
 sky130_fd_sc_hd__nor2_2 _14590_ (.A(_11713_),
    .B(_11758_),
    .Y(_11759_));
 sky130_fd_sc_hd__a32o_2 _14591_ (.A1(_11755_),
    .A2(_11757_),
    .A3(_11759_),
    .B1(\systolic_inst.acc_wires[15][9] ),
    .B2(_11258_),
    .X(_00987_));
 sky130_fd_sc_hd__nand2_2 _14592_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[15][10] ),
    .Y(_11760_));
 sky130_fd_sc_hd__or2_2 _14593_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[15][10] ),
    .X(_11761_));
 sky130_fd_sc_hd__and2_2 _14594_ (.A(_11760_),
    .B(_11761_),
    .X(_11762_));
 sky130_fd_sc_hd__a21oi_2 _14595_ (.A1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[15][9] ),
    .B1(_11758_),
    .Y(_11763_));
 sky130_fd_sc_hd__nand2_2 _14596_ (.A(_11757_),
    .B(_11763_),
    .Y(_11764_));
 sky130_fd_sc_hd__xor2_2 _14597_ (.A(_11762_),
    .B(_11764_),
    .X(_11765_));
 sky130_fd_sc_hd__a22o_2 _14598_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][10] ),
    .B1(_11712_),
    .B2(_11765_),
    .X(_00988_));
 sky130_fd_sc_hd__nor2_2 _14599_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[15][11] ),
    .Y(_11766_));
 sky130_fd_sc_hd__or2_2 _14600_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[15][11] ),
    .X(_11767_));
 sky130_fd_sc_hd__nand2_2 _14601_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[15][11] ),
    .Y(_11768_));
 sky130_fd_sc_hd__nand2_2 _14602_ (.A(_11767_),
    .B(_11768_),
    .Y(_11769_));
 sky130_fd_sc_hd__a21bo_2 _14603_ (.A1(_11762_),
    .A2(_11764_),
    .B1_N(_11760_),
    .X(_11770_));
 sky130_fd_sc_hd__xnor2_2 _14604_ (.A(_11769_),
    .B(_11770_),
    .Y(_11771_));
 sky130_fd_sc_hd__a22o_2 _14605_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][11] ),
    .B1(_11712_),
    .B2(_11771_),
    .X(_00989_));
 sky130_fd_sc_hd__nand3_2 _14606_ (.A(_11762_),
    .B(_11767_),
    .C(_11768_),
    .Y(_11772_));
 sky130_fd_sc_hd__nor2_2 _14607_ (.A(_11756_),
    .B(_11772_),
    .Y(_11773_));
 sky130_fd_sc_hd__o2bb2a_2 _14608_ (.A1_N(_11750_),
    .A2_N(_11773_),
    .B1(_11763_),
    .B2(_11772_),
    .X(_11774_));
 sky130_fd_sc_hd__o21a_2 _14609_ (.A1(_11760_),
    .A2(_11766_),
    .B1(_11768_),
    .X(_11775_));
 sky130_fd_sc_hd__xnor2_2 _14610_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[15][12] ),
    .Y(_11776_));
 sky130_fd_sc_hd__and3_2 _14611_ (.A(_11774_),
    .B(_11775_),
    .C(_11776_),
    .X(_11777_));
 sky130_fd_sc_hd__a21oi_2 _14612_ (.A1(_11774_),
    .A2(_11775_),
    .B1(_11776_),
    .Y(_11778_));
 sky130_fd_sc_hd__nor2_2 _14613_ (.A(_11777_),
    .B(_11778_),
    .Y(_11779_));
 sky130_fd_sc_hd__a22o_2 _14614_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][12] ),
    .B1(_11712_),
    .B2(_11779_),
    .X(_00990_));
 sky130_fd_sc_hd__xor2_2 _14615_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[15][13] ),
    .X(_11780_));
 sky130_fd_sc_hd__a211o_2 _14616_ (.A1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[15][12] ),
    .B1(_11778_),
    .C1(_11780_),
    .X(_11781_));
 sky130_fd_sc_hd__nand2b_2 _14617_ (.A_N(_11776_),
    .B(_11780_),
    .Y(_11782_));
 sky130_fd_sc_hd__a21o_2 _14618_ (.A1(_11774_),
    .A2(_11775_),
    .B1(_11782_),
    .X(_11783_));
 sky130_fd_sc_hd__and3_2 _14619_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[15][12] ),
    .C(_11780_),
    .X(_11784_));
 sky130_fd_sc_hd__nor2_2 _14620_ (.A(_11713_),
    .B(_11784_),
    .Y(_11785_));
 sky130_fd_sc_hd__a32o_2 _14621_ (.A1(_11781_),
    .A2(_11783_),
    .A3(_11785_),
    .B1(\systolic_inst.acc_wires[15][13] ),
    .B2(_11258_),
    .X(_00991_));
 sky130_fd_sc_hd__or2_2 _14622_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[15][14] ),
    .X(_11786_));
 sky130_fd_sc_hd__nand2_2 _14623_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[15][14] ),
    .Y(_11787_));
 sky130_fd_sc_hd__and2_2 _14624_ (.A(_11786_),
    .B(_11787_),
    .X(_11788_));
 sky130_fd_sc_hd__nand2_2 _14625_ (.A(_11786_),
    .B(_11787_),
    .Y(_11789_));
 sky130_fd_sc_hd__a21oi_2 _14626_ (.A1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[15][13] ),
    .B1(_11784_),
    .Y(_11790_));
 sky130_fd_sc_hd__nand2_2 _14627_ (.A(_11783_),
    .B(_11790_),
    .Y(_11791_));
 sky130_fd_sc_hd__nand2_2 _14628_ (.A(_11788_),
    .B(_11791_),
    .Y(_11792_));
 sky130_fd_sc_hd__or2_2 _14629_ (.A(_11788_),
    .B(_11791_),
    .X(_11793_));
 sky130_fd_sc_hd__a32o_2 _14630_ (.A1(_11712_),
    .A2(_11792_),
    .A3(_11793_),
    .B1(\systolic_inst.acc_wires[15][14] ),
    .B2(_11258_),
    .X(_00992_));
 sky130_fd_sc_hd__nor2_2 _14631_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][15] ),
    .Y(_11794_));
 sky130_fd_sc_hd__and2_2 _14632_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][15] ),
    .X(_11795_));
 sky130_fd_sc_hd__or2_2 _14633_ (.A(_11794_),
    .B(_11795_),
    .X(_11796_));
 sky130_fd_sc_hd__a21oi_2 _14634_ (.A1(_11787_),
    .A2(_11792_),
    .B1(_11796_),
    .Y(_11797_));
 sky130_fd_sc_hd__a31o_2 _14635_ (.A1(_11787_),
    .A2(_11792_),
    .A3(_11796_),
    .B1(_11713_),
    .X(_11798_));
 sky130_fd_sc_hd__a2bb2o_2 _14636_ (.A1_N(_11798_),
    .A2_N(_11797_),
    .B1(\systolic_inst.acc_wires[15][15] ),
    .B2(_11258_),
    .X(_00993_));
 sky130_fd_sc_hd__a211o_2 _14637_ (.A1(_11783_),
    .A2(_11790_),
    .B1(_11796_),
    .C1(_11789_),
    .X(_11799_));
 sky130_fd_sc_hd__o21ba_2 _14638_ (.A1(_11787_),
    .A2(_11794_),
    .B1_N(_11795_),
    .X(_11800_));
 sky130_fd_sc_hd__and2_2 _14639_ (.A(_11799_),
    .B(_11800_),
    .X(_11801_));
 sky130_fd_sc_hd__xnor2_2 _14640_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][16] ),
    .Y(_11802_));
 sky130_fd_sc_hd__nand2_2 _14641_ (.A(_11801_),
    .B(_11802_),
    .Y(_11803_));
 sky130_fd_sc_hd__nor2_2 _14642_ (.A(_11801_),
    .B(_11802_),
    .Y(_11804_));
 sky130_fd_sc_hd__nor2_2 _14643_ (.A(_11713_),
    .B(_11804_),
    .Y(_11805_));
 sky130_fd_sc_hd__a22o_2 _14644_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][16] ),
    .B1(_11803_),
    .B2(_11805_),
    .X(_00994_));
 sky130_fd_sc_hd__xor2_2 _14645_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][17] ),
    .X(_11806_));
 sky130_fd_sc_hd__inv_2 _14646_ (.A(_11806_),
    .Y(_11807_));
 sky130_fd_sc_hd__a21oi_2 _14647_ (.A1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[15][16] ),
    .B1(_11804_),
    .Y(_11808_));
 sky130_fd_sc_hd__xnor2_2 _14648_ (.A(_11806_),
    .B(_11808_),
    .Y(_11809_));
 sky130_fd_sc_hd__a22o_2 _14649_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][17] ),
    .B1(_11712_),
    .B2(_11809_),
    .X(_00995_));
 sky130_fd_sc_hd__or2_2 _14650_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][18] ),
    .X(_11810_));
 sky130_fd_sc_hd__nand2_2 _14651_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][18] ),
    .Y(_11811_));
 sky130_fd_sc_hd__nand2_2 _14652_ (.A(_11810_),
    .B(_11811_),
    .Y(_11812_));
 sky130_fd_sc_hd__o21a_2 _14653_ (.A1(\systolic_inst.acc_wires[15][16] ),
    .A2(\systolic_inst.acc_wires[15][17] ),
    .B1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .X(_11813_));
 sky130_fd_sc_hd__a21oi_2 _14654_ (.A1(_11804_),
    .A2(_11806_),
    .B1(_11813_),
    .Y(_11814_));
 sky130_fd_sc_hd__xor2_2 _14655_ (.A(_11812_),
    .B(_11814_),
    .X(_11815_));
 sky130_fd_sc_hd__a22o_2 _14656_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][18] ),
    .B1(_11712_),
    .B2(_11815_),
    .X(_00996_));
 sky130_fd_sc_hd__xnor2_2 _14657_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][19] ),
    .Y(_11816_));
 sky130_fd_sc_hd__o21ai_2 _14658_ (.A1(_11812_),
    .A2(_11814_),
    .B1(_11811_),
    .Y(_11817_));
 sky130_fd_sc_hd__xnor2_2 _14659_ (.A(_11816_),
    .B(_11817_),
    .Y(_11818_));
 sky130_fd_sc_hd__a22o_2 _14660_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][19] ),
    .B1(_11712_),
    .B2(_11818_),
    .X(_00997_));
 sky130_fd_sc_hd__or2_2 _14661_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][20] ),
    .X(_11819_));
 sky130_fd_sc_hd__nand2_2 _14662_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][20] ),
    .Y(_11820_));
 sky130_fd_sc_hd__and2_2 _14663_ (.A(_11819_),
    .B(_11820_),
    .X(_11821_));
 sky130_fd_sc_hd__or4_2 _14664_ (.A(_11802_),
    .B(_11807_),
    .C(_11812_),
    .D(_11816_),
    .X(_11822_));
 sky130_fd_sc_hd__nor2_2 _14665_ (.A(_11801_),
    .B(_11822_),
    .Y(_11823_));
 sky130_fd_sc_hd__o41a_2 _14666_ (.A1(\systolic_inst.acc_wires[15][16] ),
    .A2(\systolic_inst.acc_wires[15][17] ),
    .A3(\systolic_inst.acc_wires[15][18] ),
    .A4(\systolic_inst.acc_wires[15][19] ),
    .B1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .X(_11824_));
 sky130_fd_sc_hd__or3_2 _14667_ (.A(_11821_),
    .B(_11823_),
    .C(_11824_),
    .X(_11825_));
 sky130_fd_sc_hd__o21ai_2 _14668_ (.A1(_11823_),
    .A2(_11824_),
    .B1(_11821_),
    .Y(_11826_));
 sky130_fd_sc_hd__a32o_2 _14669_ (.A1(_11712_),
    .A2(_11825_),
    .A3(_11826_),
    .B1(\systolic_inst.acc_wires[15][20] ),
    .B2(_11258_),
    .X(_00998_));
 sky130_fd_sc_hd__xnor2_2 _14670_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][21] ),
    .Y(_11827_));
 sky130_fd_sc_hd__inv_2 _14671_ (.A(_11827_),
    .Y(_11828_));
 sky130_fd_sc_hd__a21oi_2 _14672_ (.A1(_11820_),
    .A2(_11826_),
    .B1(_11827_),
    .Y(_11829_));
 sky130_fd_sc_hd__a31o_2 _14673_ (.A1(_11820_),
    .A2(_11826_),
    .A3(_11827_),
    .B1(_11713_),
    .X(_11830_));
 sky130_fd_sc_hd__a2bb2o_2 _14674_ (.A1_N(_11830_),
    .A2_N(_11829_),
    .B1(\systolic_inst.acc_wires[15][21] ),
    .B2(_11258_),
    .X(_00999_));
 sky130_fd_sc_hd__or2_2 _14675_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][22] ),
    .X(_11831_));
 sky130_fd_sc_hd__nand2_2 _14676_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][22] ),
    .Y(_11832_));
 sky130_fd_sc_hd__and2_2 _14677_ (.A(_11831_),
    .B(_11832_),
    .X(_11833_));
 sky130_fd_sc_hd__o21a_2 _14678_ (.A1(\systolic_inst.acc_wires[15][20] ),
    .A2(\systolic_inst.acc_wires[15][21] ),
    .B1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .X(_11834_));
 sky130_fd_sc_hd__nor2_2 _14679_ (.A(_11826_),
    .B(_11827_),
    .Y(_11835_));
 sky130_fd_sc_hd__o21ai_2 _14680_ (.A1(_11834_),
    .A2(_11835_),
    .B1(_11833_),
    .Y(_11836_));
 sky130_fd_sc_hd__or3_2 _14681_ (.A(_11833_),
    .B(_11834_),
    .C(_11835_),
    .X(_11837_));
 sky130_fd_sc_hd__a32o_2 _14682_ (.A1(_11712_),
    .A2(_11836_),
    .A3(_11837_),
    .B1(\systolic_inst.acc_wires[15][22] ),
    .B2(_11258_),
    .X(_01000_));
 sky130_fd_sc_hd__xor2_2 _14683_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][23] ),
    .X(_11838_));
 sky130_fd_sc_hd__inv_2 _14684_ (.A(_11838_),
    .Y(_11839_));
 sky130_fd_sc_hd__nand3_2 _14685_ (.A(_11832_),
    .B(_11836_),
    .C(_11839_),
    .Y(_11840_));
 sky130_fd_sc_hd__a21o_2 _14686_ (.A1(_11832_),
    .A2(_11836_),
    .B1(_11839_),
    .X(_11841_));
 sky130_fd_sc_hd__a32o_2 _14687_ (.A1(_11712_),
    .A2(_11840_),
    .A3(_11841_),
    .B1(\systolic_inst.acc_wires[15][23] ),
    .B2(_11258_),
    .X(_01001_));
 sky130_fd_sc_hd__nand4_2 _14688_ (.A(_11821_),
    .B(_11828_),
    .C(_11833_),
    .D(_11838_),
    .Y(_11842_));
 sky130_fd_sc_hd__a211o_2 _14689_ (.A1(_11799_),
    .A2(_11800_),
    .B1(_11822_),
    .C1(_11842_),
    .X(_11843_));
 sky130_fd_sc_hd__o41a_2 _14690_ (.A1(\systolic_inst.acc_wires[15][20] ),
    .A2(\systolic_inst.acc_wires[15][21] ),
    .A3(\systolic_inst.acc_wires[15][22] ),
    .A4(\systolic_inst.acc_wires[15][23] ),
    .B1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .X(_11844_));
 sky130_fd_sc_hd__nor2_2 _14691_ (.A(_11824_),
    .B(_11844_),
    .Y(_11845_));
 sky130_fd_sc_hd__nor2_2 _14692_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][24] ),
    .Y(_11846_));
 sky130_fd_sc_hd__and2_2 _14693_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][24] ),
    .X(_11847_));
 sky130_fd_sc_hd__or2_2 _14694_ (.A(_11846_),
    .B(_11847_),
    .X(_11848_));
 sky130_fd_sc_hd__and3_2 _14695_ (.A(_11843_),
    .B(_11845_),
    .C(_11848_),
    .X(_11849_));
 sky130_fd_sc_hd__a21oi_2 _14696_ (.A1(_11843_),
    .A2(_11845_),
    .B1(_11848_),
    .Y(_11850_));
 sky130_fd_sc_hd__nor2_2 _14697_ (.A(_11849_),
    .B(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__a22o_2 _14698_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][24] ),
    .B1(_11712_),
    .B2(_11851_),
    .X(_01002_));
 sky130_fd_sc_hd__xor2_2 _14699_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][25] ),
    .X(_11852_));
 sky130_fd_sc_hd__or3_2 _14700_ (.A(_11847_),
    .B(_11850_),
    .C(_11852_),
    .X(_11853_));
 sky130_fd_sc_hd__o21ai_2 _14701_ (.A1(_11847_),
    .A2(_11850_),
    .B1(_11852_),
    .Y(_11854_));
 sky130_fd_sc_hd__a32o_2 _14702_ (.A1(_11712_),
    .A2(_11853_),
    .A3(_11854_),
    .B1(\systolic_inst.acc_wires[15][25] ),
    .B2(_11258_),
    .X(_01003_));
 sky130_fd_sc_hd__or2_2 _14703_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][26] ),
    .X(_11855_));
 sky130_fd_sc_hd__nand2_2 _14704_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][26] ),
    .Y(_11856_));
 sky130_fd_sc_hd__nand2_2 _14705_ (.A(_11855_),
    .B(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__o21a_2 _14706_ (.A1(\systolic_inst.acc_wires[15][24] ),
    .A2(\systolic_inst.acc_wires[15][25] ),
    .B1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .X(_11858_));
 sky130_fd_sc_hd__a21o_2 _14707_ (.A1(_11850_),
    .A2(_11852_),
    .B1(_11858_),
    .X(_11859_));
 sky130_fd_sc_hd__xnor2_2 _14708_ (.A(_11857_),
    .B(_11859_),
    .Y(_11860_));
 sky130_fd_sc_hd__a22o_2 _14709_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][26] ),
    .B1(_11712_),
    .B2(_11860_),
    .X(_01004_));
 sky130_fd_sc_hd__xnor2_2 _14710_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][27] ),
    .Y(_11861_));
 sky130_fd_sc_hd__a21bo_2 _14711_ (.A1(_11855_),
    .A2(_11859_),
    .B1_N(_11856_),
    .X(_11862_));
 sky130_fd_sc_hd__xnor2_2 _14712_ (.A(_11861_),
    .B(_11862_),
    .Y(_11863_));
 sky130_fd_sc_hd__a22o_2 _14713_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][27] ),
    .B1(_11712_),
    .B2(_11863_),
    .X(_01005_));
 sky130_fd_sc_hd__nor2_2 _14714_ (.A(_11857_),
    .B(_11861_),
    .Y(_11864_));
 sky130_fd_sc_hd__o21a_2 _14715_ (.A1(\systolic_inst.acc_wires[15][26] ),
    .A2(\systolic_inst.acc_wires[15][27] ),
    .B1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .X(_11865_));
 sky130_fd_sc_hd__a311oi_2 _14716_ (.A1(_11850_),
    .A2(_11852_),
    .A3(_11864_),
    .B1(_11865_),
    .C1(_11858_),
    .Y(_11866_));
 sky130_fd_sc_hd__or2_2 _14717_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][28] ),
    .X(_11867_));
 sky130_fd_sc_hd__nand2_2 _14718_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][28] ),
    .Y(_11868_));
 sky130_fd_sc_hd__nand2_2 _14719_ (.A(_11867_),
    .B(_11868_),
    .Y(_11869_));
 sky130_fd_sc_hd__or2_2 _14720_ (.A(_11866_),
    .B(_11869_),
    .X(_11870_));
 sky130_fd_sc_hd__nand2_2 _14721_ (.A(_11866_),
    .B(_11869_),
    .Y(_11871_));
 sky130_fd_sc_hd__a32o_2 _14722_ (.A1(_11712_),
    .A2(_11870_),
    .A3(_11871_),
    .B1(\systolic_inst.acc_wires[15][28] ),
    .B2(_11258_),
    .X(_01006_));
 sky130_fd_sc_hd__xor2_2 _14723_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][29] ),
    .X(_11872_));
 sky130_fd_sc_hd__inv_2 _14724_ (.A(_11872_),
    .Y(_11873_));
 sky130_fd_sc_hd__o21a_2 _14725_ (.A1(_11866_),
    .A2(_11869_),
    .B1(_11868_),
    .X(_11874_));
 sky130_fd_sc_hd__xnor2_2 _14726_ (.A(_11872_),
    .B(_11874_),
    .Y(_11875_));
 sky130_fd_sc_hd__a22o_2 _14727_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[15][29] ),
    .B1(_11712_),
    .B2(_11875_),
    .X(_01007_));
 sky130_fd_sc_hd__o21ai_2 _14728_ (.A1(\systolic_inst.acc_wires[15][28] ),
    .A2(\systolic_inst.acc_wires[15][29] ),
    .B1(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .Y(_11876_));
 sky130_fd_sc_hd__o31a_2 _14729_ (.A1(_11866_),
    .A2(_11869_),
    .A3(_11873_),
    .B1(_11876_),
    .X(_11877_));
 sky130_fd_sc_hd__nand2_2 _14730_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][30] ),
    .Y(_11878_));
 sky130_fd_sc_hd__or2_2 _14731_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][30] ),
    .X(_11879_));
 sky130_fd_sc_hd__nand2_2 _14732_ (.A(_11878_),
    .B(_11879_),
    .Y(_11880_));
 sky130_fd_sc_hd__nand2_2 _14733_ (.A(_11877_),
    .B(_11880_),
    .Y(_11881_));
 sky130_fd_sc_hd__or2_2 _14734_ (.A(_11877_),
    .B(_11880_),
    .X(_11882_));
 sky130_fd_sc_hd__a32o_2 _14735_ (.A1(_11712_),
    .A2(_11881_),
    .A3(_11882_),
    .B1(\systolic_inst.acc_wires[15][30] ),
    .B2(_11258_),
    .X(_01008_));
 sky130_fd_sc_hd__xnor2_2 _14736_ (.A(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[15][31] ),
    .Y(_11883_));
 sky130_fd_sc_hd__a21oi_2 _14737_ (.A1(_11878_),
    .A2(_11882_),
    .B1(_11883_),
    .Y(_11884_));
 sky130_fd_sc_hd__a31o_2 _14738_ (.A1(_11878_),
    .A2(_11882_),
    .A3(_11883_),
    .B1(_11713_),
    .X(_11885_));
 sky130_fd_sc_hd__a2bb2o_2 _14739_ (.A1_N(_11885_),
    .A2_N(_11884_),
    .B1(\systolic_inst.acc_wires[15][31] ),
    .B2(_11258_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _14740_ (.A0(\systolic_inst.A_outs[14][0] ),
    .A1(\systolic_inst.A_outs[13][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _14741_ (.A0(\systolic_inst.A_outs[14][1] ),
    .A1(\systolic_inst.A_outs[13][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _14742_ (.A0(\systolic_inst.A_outs[14][2] ),
    .A1(\systolic_inst.A_outs[13][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _14743_ (.A0(\systolic_inst.A_outs[14][3] ),
    .A1(\systolic_inst.A_outs[13][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _14744_ (.A0(\systolic_inst.A_outs[14][4] ),
    .A1(\systolic_inst.A_outs[13][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _14745_ (.A0(\systolic_inst.A_outs[14][5] ),
    .A1(\systolic_inst.A_outs[13][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _14746_ (.A0(\systolic_inst.A_outs[14][6] ),
    .A1(\systolic_inst.A_outs[13][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _14747_ (.A0(\systolic_inst.A_outs[14][7] ),
    .A1(\systolic_inst.A_outs[13][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _14748_ (.A0(\systolic_inst.B_outs[13][0] ),
    .A1(\systolic_inst.B_outs[9][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _14749_ (.A0(\systolic_inst.B_outs[13][1] ),
    .A1(\systolic_inst.B_outs[9][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _14750_ (.A0(\systolic_inst.B_outs[13][2] ),
    .A1(\systolic_inst.B_outs[9][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _14751_ (.A0(\systolic_inst.B_outs[13][3] ),
    .A1(\systolic_inst.B_outs[9][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _14752_ (.A0(\systolic_inst.B_outs[13][4] ),
    .A1(\systolic_inst.B_outs[9][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _14753_ (.A0(\systolic_inst.B_outs[13][5] ),
    .A1(\systolic_inst.B_outs[9][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _14754_ (.A0(\systolic_inst.B_outs[13][6] ),
    .A1(\systolic_inst.B_outs[9][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _14755_ (.A0(\systolic_inst.B_outs[13][7] ),
    .A1(\systolic_inst.B_outs[9][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01025_));
 sky130_fd_sc_hd__and3_2 _14756_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[14][0] ),
    .C(\systolic_inst.A_outs[14][0] ),
    .X(_11886_));
 sky130_fd_sc_hd__a21o_2 _14757_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[0] ),
    .B1(_11886_),
    .X(_01026_));
 sky130_fd_sc_hd__and4_2 _14758_ (.A(\systolic_inst.B_outs[14][0] ),
    .B(\systolic_inst.A_outs[14][0] ),
    .C(\systolic_inst.B_outs[14][1] ),
    .D(\systolic_inst.A_outs[14][1] ),
    .X(_11887_));
 sky130_fd_sc_hd__inv_2 _14759_ (.A(_11887_),
    .Y(_11888_));
 sky130_fd_sc_hd__a22o_2 _14760_ (.A1(\systolic_inst.A_outs[14][0] ),
    .A2(\systolic_inst.B_outs[14][1] ),
    .B1(\systolic_inst.A_outs[14][1] ),
    .B2(\systolic_inst.B_outs[14][0] ),
    .X(_11889_));
 sky130_fd_sc_hd__and2_2 _14761_ (.A(\systolic_inst.ce_local ),
    .B(_11889_),
    .X(_11890_));
 sky130_fd_sc_hd__a22o_2 _14762_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[1] ),
    .B1(_11888_),
    .B2(_11890_),
    .X(_01027_));
 sky130_fd_sc_hd__nand2_2 _14763_ (.A(\systolic_inst.B_outs[14][1] ),
    .B(\systolic_inst.A_outs[14][1] ),
    .Y(_11891_));
 sky130_fd_sc_hd__nand2_2 _14764_ (.A(\systolic_inst.B_outs[14][0] ),
    .B(\systolic_inst.A_outs[14][2] ),
    .Y(_11892_));
 sky130_fd_sc_hd__and4_2 _14765_ (.A(\systolic_inst.B_outs[14][0] ),
    .B(\systolic_inst.B_outs[14][1] ),
    .C(\systolic_inst.A_outs[14][1] ),
    .D(\systolic_inst.A_outs[14][2] ),
    .X(_11893_));
 sky130_fd_sc_hd__a21o_2 _14766_ (.A1(_11891_),
    .A2(_11892_),
    .B1(_11893_),
    .X(_11894_));
 sky130_fd_sc_hd__xnor2_2 _14767_ (.A(_11887_),
    .B(_11894_),
    .Y(_11895_));
 sky130_fd_sc_hd__and2_2 _14768_ (.A(\systolic_inst.A_outs[14][0] ),
    .B(\systolic_inst.B_outs[14][2] ),
    .X(_11896_));
 sky130_fd_sc_hd__nand2_2 _14769_ (.A(_11895_),
    .B(_11896_),
    .Y(_11897_));
 sky130_fd_sc_hd__o21a_2 _14770_ (.A1(_11895_),
    .A2(_11896_),
    .B1(\systolic_inst.ce_local ),
    .X(_11898_));
 sky130_fd_sc_hd__a22o_2 _14771_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[2] ),
    .B1(_11897_),
    .B2(_11898_),
    .X(_01028_));
 sky130_fd_sc_hd__a22oi_2 _14772_ (.A1(\systolic_inst.A_outs[14][1] ),
    .A2(\systolic_inst.B_outs[14][2] ),
    .B1(\systolic_inst.B_outs[14][3] ),
    .B2(\systolic_inst.A_outs[14][0] ),
    .Y(_11899_));
 sky130_fd_sc_hd__and4_2 _14773_ (.A(\systolic_inst.A_outs[14][0] ),
    .B(\systolic_inst.A_outs[14][1] ),
    .C(\systolic_inst.B_outs[14][2] ),
    .D(\systolic_inst.B_outs[14][3] ),
    .X(_11900_));
 sky130_fd_sc_hd__or2_2 _14774_ (.A(_11899_),
    .B(_11900_),
    .X(_11901_));
 sky130_fd_sc_hd__nand2_2 _14775_ (.A(\systolic_inst.B_outs[14][1] ),
    .B(\systolic_inst.A_outs[14][3] ),
    .Y(_11902_));
 sky130_fd_sc_hd__or2_2 _14776_ (.A(_11892_),
    .B(_11902_),
    .X(_11903_));
 sky130_fd_sc_hd__a22o_2 _14777_ (.A1(\systolic_inst.B_outs[14][1] ),
    .A2(\systolic_inst.A_outs[14][2] ),
    .B1(\systolic_inst.A_outs[14][3] ),
    .B2(\systolic_inst.B_outs[14][0] ),
    .X(_11904_));
 sky130_fd_sc_hd__nand3_2 _14778_ (.A(_11893_),
    .B(_11903_),
    .C(_11904_),
    .Y(_11905_));
 sky130_fd_sc_hd__a21o_2 _14779_ (.A1(_11903_),
    .A2(_11904_),
    .B1(_11893_),
    .X(_11906_));
 sky130_fd_sc_hd__nand2_2 _14780_ (.A(_11905_),
    .B(_11906_),
    .Y(_11907_));
 sky130_fd_sc_hd__or2_2 _14781_ (.A(_11901_),
    .B(_11907_),
    .X(_11908_));
 sky130_fd_sc_hd__xnor2_2 _14782_ (.A(_11901_),
    .B(_11907_),
    .Y(_11909_));
 sky130_fd_sc_hd__o21ai_2 _14783_ (.A1(_11888_),
    .A2(_11894_),
    .B1(_11897_),
    .Y(_11910_));
 sky130_fd_sc_hd__and2b_2 _14784_ (.A_N(_11909_),
    .B(_11910_),
    .X(_11911_));
 sky130_fd_sc_hd__xnor2_2 _14785_ (.A(_11909_),
    .B(_11910_),
    .Y(_11912_));
 sky130_fd_sc_hd__mux2_1 _14786_ (.A0(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[3] ),
    .A1(_11912_),
    .S(\systolic_inst.ce_local ),
    .X(_01029_));
 sky130_fd_sc_hd__and2_2 _14787_ (.A(\systolic_inst.B_outs[14][2] ),
    .B(\systolic_inst.A_outs[14][2] ),
    .X(_11913_));
 sky130_fd_sc_hd__nand4_2 _14788_ (.A(\systolic_inst.A_outs[14][0] ),
    .B(\systolic_inst.A_outs[14][1] ),
    .C(\systolic_inst.B_outs[14][3] ),
    .D(\systolic_inst.B_outs[14][4] ),
    .Y(_11914_));
 sky130_fd_sc_hd__a22o_2 _14789_ (.A1(\systolic_inst.A_outs[14][1] ),
    .A2(\systolic_inst.B_outs[14][3] ),
    .B1(\systolic_inst.B_outs[14][4] ),
    .B2(\systolic_inst.A_outs[14][0] ),
    .X(_11915_));
 sky130_fd_sc_hd__nand2_2 _14790_ (.A(_11914_),
    .B(_11915_),
    .Y(_11916_));
 sky130_fd_sc_hd__xnor2_2 _14791_ (.A(_11913_),
    .B(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__inv_2 _14792_ (.A(_11917_),
    .Y(_11918_));
 sky130_fd_sc_hd__nand2_2 _14793_ (.A(\systolic_inst.B_outs[14][0] ),
    .B(\systolic_inst.A_outs[14][4] ),
    .Y(_11919_));
 sky130_fd_sc_hd__and4_2 _14794_ (.A(\systolic_inst.B_outs[14][0] ),
    .B(\systolic_inst.B_outs[14][1] ),
    .C(\systolic_inst.A_outs[14][3] ),
    .D(\systolic_inst.A_outs[14][4] ),
    .X(_11920_));
 sky130_fd_sc_hd__a21oi_2 _14795_ (.A1(_11902_),
    .A2(_11919_),
    .B1(_11920_),
    .Y(_11921_));
 sky130_fd_sc_hd__xnor2_2 _14796_ (.A(_11900_),
    .B(_11921_),
    .Y(_11922_));
 sky130_fd_sc_hd__nor2_2 _14797_ (.A(_11903_),
    .B(_11922_),
    .Y(_11923_));
 sky130_fd_sc_hd__xnor2_2 _14798_ (.A(_11903_),
    .B(_11922_),
    .Y(_11924_));
 sky130_fd_sc_hd__nor2_2 _14799_ (.A(_11918_),
    .B(_11924_),
    .Y(_11925_));
 sky130_fd_sc_hd__xnor2_2 _14800_ (.A(_11918_),
    .B(_11924_),
    .Y(_11926_));
 sky130_fd_sc_hd__a21o_2 _14801_ (.A1(_11905_),
    .A2(_11908_),
    .B1(_11926_),
    .X(_11927_));
 sky130_fd_sc_hd__inv_2 _14802_ (.A(_11927_),
    .Y(_11928_));
 sky130_fd_sc_hd__nand3_2 _14803_ (.A(_11905_),
    .B(_11908_),
    .C(_11926_),
    .Y(_11929_));
 sky130_fd_sc_hd__a21oi_2 _14804_ (.A1(_11927_),
    .A2(_11929_),
    .B1(_11911_),
    .Y(_11930_));
 sky130_fd_sc_hd__and3_2 _14805_ (.A(_11911_),
    .B(_11927_),
    .C(_11929_),
    .X(_11931_));
 sky130_fd_sc_hd__or3_2 _14806_ (.A(_11258_),
    .B(_11930_),
    .C(_11931_),
    .X(_11932_));
 sky130_fd_sc_hd__a21bo_2 _14807_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[4] ),
    .B1_N(_11932_),
    .X(_01030_));
 sky130_fd_sc_hd__a21oi_2 _14808_ (.A1(_11900_),
    .A2(_11921_),
    .B1(_11923_),
    .Y(_11933_));
 sky130_fd_sc_hd__a21bo_2 _14809_ (.A1(_11913_),
    .A2(_11915_),
    .B1_N(_11914_),
    .X(_11934_));
 sky130_fd_sc_hd__a22oi_2 _14810_ (.A1(\systolic_inst.B_outs[14][1] ),
    .A2(\systolic_inst.A_outs[14][4] ),
    .B1(\systolic_inst.A_outs[14][5] ),
    .B2(\systolic_inst.B_outs[14][0] ),
    .Y(_11935_));
 sky130_fd_sc_hd__and4_2 _14811_ (.A(\systolic_inst.B_outs[14][0] ),
    .B(\systolic_inst.B_outs[14][1] ),
    .C(\systolic_inst.A_outs[14][4] ),
    .D(\systolic_inst.A_outs[14][5] ),
    .X(_11936_));
 sky130_fd_sc_hd__or2_2 _14812_ (.A(_11935_),
    .B(_11936_),
    .X(_11937_));
 sky130_fd_sc_hd__nand2b_2 _14813_ (.A_N(_11937_),
    .B(_11934_),
    .Y(_11938_));
 sky130_fd_sc_hd__xnor2_2 _14814_ (.A(_11934_),
    .B(_11937_),
    .Y(_11939_));
 sky130_fd_sc_hd__nand2_2 _14815_ (.A(_11920_),
    .B(_11939_),
    .Y(_11940_));
 sky130_fd_sc_hd__xnor2_2 _14816_ (.A(_11920_),
    .B(_11939_),
    .Y(_11941_));
 sky130_fd_sc_hd__nand2_2 _14817_ (.A(\systolic_inst.A_outs[14][0] ),
    .B(\systolic_inst.B_outs[14][5] ),
    .Y(_11942_));
 sky130_fd_sc_hd__nand2_2 _14818_ (.A(\systolic_inst.B_outs[14][2] ),
    .B(\systolic_inst.A_outs[14][3] ),
    .Y(_11943_));
 sky130_fd_sc_hd__and4_2 _14819_ (.A(\systolic_inst.A_outs[14][1] ),
    .B(\systolic_inst.A_outs[14][2] ),
    .C(\systolic_inst.B_outs[14][3] ),
    .D(\systolic_inst.B_outs[14][4] ),
    .X(_11944_));
 sky130_fd_sc_hd__a22o_2 _14820_ (.A1(\systolic_inst.A_outs[14][2] ),
    .A2(\systolic_inst.B_outs[14][3] ),
    .B1(\systolic_inst.B_outs[14][4] ),
    .B2(\systolic_inst.A_outs[14][1] ),
    .X(_11945_));
 sky130_fd_sc_hd__and2b_2 _14821_ (.A_N(_11944_),
    .B(_11945_),
    .X(_11946_));
 sky130_fd_sc_hd__xnor2_2 _14822_ (.A(_11943_),
    .B(_11946_),
    .Y(_11947_));
 sky130_fd_sc_hd__nand2b_2 _14823_ (.A_N(_11942_),
    .B(_11947_),
    .Y(_11948_));
 sky130_fd_sc_hd__xor2_2 _14824_ (.A(_11942_),
    .B(_11947_),
    .X(_11949_));
 sky130_fd_sc_hd__nor2_2 _14825_ (.A(_11941_),
    .B(_11949_),
    .Y(_11950_));
 sky130_fd_sc_hd__inv_2 _14826_ (.A(_11950_),
    .Y(_11951_));
 sky130_fd_sc_hd__xor2_2 _14827_ (.A(_11941_),
    .B(_11949_),
    .X(_11952_));
 sky130_fd_sc_hd__nand2_2 _14828_ (.A(_11925_),
    .B(_11952_),
    .Y(_11953_));
 sky130_fd_sc_hd__or2_2 _14829_ (.A(_11925_),
    .B(_11952_),
    .X(_11954_));
 sky130_fd_sc_hd__and2_2 _14830_ (.A(_11953_),
    .B(_11954_),
    .X(_11955_));
 sky130_fd_sc_hd__nand2b_2 _14831_ (.A_N(_11933_),
    .B(_11955_),
    .Y(_11956_));
 sky130_fd_sc_hd__xnor2_2 _14832_ (.A(_11933_),
    .B(_11955_),
    .Y(_11957_));
 sky130_fd_sc_hd__nor2_2 _14833_ (.A(_11928_),
    .B(_11931_),
    .Y(_11958_));
 sky130_fd_sc_hd__nand2b_2 _14834_ (.A_N(_11958_),
    .B(_11957_),
    .Y(_11959_));
 sky130_fd_sc_hd__o31a_2 _14835_ (.A1(_11928_),
    .A2(_11931_),
    .A3(_11957_),
    .B1(\systolic_inst.ce_local ),
    .X(_11960_));
 sky130_fd_sc_hd__a22o_2 _14836_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[5] ),
    .B1(_11959_),
    .B2(_11960_),
    .X(_01031_));
 sky130_fd_sc_hd__a31o_2 _14837_ (.A1(\systolic_inst.B_outs[14][2] ),
    .A2(\systolic_inst.A_outs[14][3] ),
    .A3(_11945_),
    .B1(_11944_),
    .X(_11961_));
 sky130_fd_sc_hd__a22oi_2 _14838_ (.A1(\systolic_inst.B_outs[14][1] ),
    .A2(\systolic_inst.A_outs[14][5] ),
    .B1(\systolic_inst.A_outs[14][6] ),
    .B2(\systolic_inst.B_outs[14][0] ),
    .Y(_11962_));
 sky130_fd_sc_hd__and4_2 _14839_ (.A(\systolic_inst.B_outs[14][0] ),
    .B(\systolic_inst.B_outs[14][1] ),
    .C(\systolic_inst.A_outs[14][5] ),
    .D(\systolic_inst.A_outs[14][6] ),
    .X(_11963_));
 sky130_fd_sc_hd__nor2_2 _14840_ (.A(_11962_),
    .B(_11963_),
    .Y(_11964_));
 sky130_fd_sc_hd__xor2_2 _14841_ (.A(_11961_),
    .B(_11964_),
    .X(_11965_));
 sky130_fd_sc_hd__and2_2 _14842_ (.A(_11936_),
    .B(_11965_),
    .X(_11966_));
 sky130_fd_sc_hd__nor2_2 _14843_ (.A(_11936_),
    .B(_11965_),
    .Y(_11967_));
 sky130_fd_sc_hd__or2_2 _14844_ (.A(_11966_),
    .B(_11967_),
    .X(_11968_));
 sky130_fd_sc_hd__nand2_2 _14845_ (.A(\systolic_inst.B_outs[14][2] ),
    .B(\systolic_inst.A_outs[14][4] ),
    .Y(_11969_));
 sky130_fd_sc_hd__and4_2 _14846_ (.A(\systolic_inst.A_outs[14][2] ),
    .B(\systolic_inst.B_outs[14][3] ),
    .C(\systolic_inst.A_outs[14][3] ),
    .D(\systolic_inst.B_outs[14][4] ),
    .X(_11970_));
 sky130_fd_sc_hd__a22oi_2 _14847_ (.A1(\systolic_inst.B_outs[14][3] ),
    .A2(\systolic_inst.A_outs[14][3] ),
    .B1(\systolic_inst.B_outs[14][4] ),
    .B2(\systolic_inst.A_outs[14][2] ),
    .Y(_11971_));
 sky130_fd_sc_hd__or2_2 _14848_ (.A(_11970_),
    .B(_11971_),
    .X(_11972_));
 sky130_fd_sc_hd__xnor2_2 _14849_ (.A(_11969_),
    .B(_11972_),
    .Y(_11973_));
 sky130_fd_sc_hd__a22oi_2 _14850_ (.A1(\systolic_inst.A_outs[14][1] ),
    .A2(\systolic_inst.B_outs[14][5] ),
    .B1(\systolic_inst.B_outs[14][6] ),
    .B2(\systolic_inst.A_outs[14][0] ),
    .Y(_11974_));
 sky130_fd_sc_hd__nand2_2 _14851_ (.A(\systolic_inst.A_outs[14][1] ),
    .B(\systolic_inst.B_outs[14][6] ),
    .Y(_11975_));
 sky130_fd_sc_hd__nor2_2 _14852_ (.A(_11942_),
    .B(_11975_),
    .Y(_11976_));
 sky130_fd_sc_hd__nor2_2 _14853_ (.A(_11974_),
    .B(_11976_),
    .Y(_11977_));
 sky130_fd_sc_hd__or3_2 _14854_ (.A(_11973_),
    .B(_11974_),
    .C(_11976_),
    .X(_11978_));
 sky130_fd_sc_hd__xor2_2 _14855_ (.A(_11973_),
    .B(_11977_),
    .X(_11979_));
 sky130_fd_sc_hd__xnor2_2 _14856_ (.A(_11948_),
    .B(_11979_),
    .Y(_11980_));
 sky130_fd_sc_hd__xnor2_2 _14857_ (.A(_11968_),
    .B(_11980_),
    .Y(_11981_));
 sky130_fd_sc_hd__xnor2_2 _14858_ (.A(_11951_),
    .B(_11981_),
    .Y(_11982_));
 sky130_fd_sc_hd__a21oi_2 _14859_ (.A1(_11938_),
    .A2(_11940_),
    .B1(_11982_),
    .Y(_11983_));
 sky130_fd_sc_hd__and3_2 _14860_ (.A(_11938_),
    .B(_11940_),
    .C(_11982_),
    .X(_11984_));
 sky130_fd_sc_hd__a211oi_2 _14861_ (.A1(_11953_),
    .A2(_11956_),
    .B1(_11983_),
    .C1(_11984_),
    .Y(_11985_));
 sky130_fd_sc_hd__o211a_2 _14862_ (.A1(_11983_),
    .A2(_11984_),
    .B1(_11953_),
    .C1(_11956_),
    .X(_11986_));
 sky130_fd_sc_hd__o21ai_2 _14863_ (.A1(_11985_),
    .A2(_11986_),
    .B1(_11959_),
    .Y(_11987_));
 sky130_fd_sc_hd__nor3_2 _14864_ (.A(_11959_),
    .B(_11985_),
    .C(_11986_),
    .Y(_11988_));
 sky130_fd_sc_hd__nor2_2 _14865_ (.A(_11258_),
    .B(_11988_),
    .Y(_11989_));
 sky130_fd_sc_hd__a22o_2 _14866_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[6] ),
    .B1(_11987_),
    .B2(_11989_),
    .X(_01032_));
 sky130_fd_sc_hd__o21ba_2 _14867_ (.A1(_11951_),
    .A2(_11981_),
    .B1_N(_11983_),
    .X(_11990_));
 sky130_fd_sc_hd__a21oi_2 _14868_ (.A1(_11961_),
    .A2(_11964_),
    .B1(_11966_),
    .Y(_11991_));
 sky130_fd_sc_hd__o21ba_2 _14869_ (.A1(_11969_),
    .A2(_11971_),
    .B1_N(_11970_),
    .X(_11992_));
 sky130_fd_sc_hd__a22o_2 _14870_ (.A1(\systolic_inst.B_outs[14][1] ),
    .A2(\systolic_inst.A_outs[14][6] ),
    .B1(\systolic_inst.A_outs[14][7] ),
    .B2(\systolic_inst.B_outs[14][0] ),
    .X(_11993_));
 sky130_fd_sc_hd__nand4_2 _14871_ (.A(\systolic_inst.B_outs[14][0] ),
    .B(\systolic_inst.B_outs[14][1] ),
    .C(\systolic_inst.A_outs[14][6] ),
    .D(\systolic_inst.A_outs[14][7] ),
    .Y(_11994_));
 sky130_fd_sc_hd__nand2_2 _14872_ (.A(_11993_),
    .B(_11994_),
    .Y(_11995_));
 sky130_fd_sc_hd__xnor2_2 _14873_ (.A(_11264_),
    .B(_11995_),
    .Y(_11996_));
 sky130_fd_sc_hd__nor2_2 _14874_ (.A(_11992_),
    .B(_11996_),
    .Y(_11997_));
 sky130_fd_sc_hd__and2_2 _14875_ (.A(_11992_),
    .B(_11996_),
    .X(_11998_));
 sky130_fd_sc_hd__nor2_2 _14876_ (.A(_11997_),
    .B(_11998_),
    .Y(_11999_));
 sky130_fd_sc_hd__xnor2_2 _14877_ (.A(_11963_),
    .B(_11999_),
    .Y(_12000_));
 sky130_fd_sc_hd__nand2_2 _14878_ (.A(\systolic_inst.B_outs[14][2] ),
    .B(\systolic_inst.A_outs[14][5] ),
    .Y(_12001_));
 sky130_fd_sc_hd__and4_2 _14879_ (.A(\systolic_inst.B_outs[14][3] ),
    .B(\systolic_inst.A_outs[14][3] ),
    .C(\systolic_inst.B_outs[14][4] ),
    .D(\systolic_inst.A_outs[14][4] ),
    .X(_12002_));
 sky130_fd_sc_hd__a22oi_2 _14880_ (.A1(\systolic_inst.A_outs[14][3] ),
    .A2(\systolic_inst.B_outs[14][4] ),
    .B1(\systolic_inst.A_outs[14][4] ),
    .B2(\systolic_inst.B_outs[14][3] ),
    .Y(_12003_));
 sky130_fd_sc_hd__or2_2 _14881_ (.A(_12002_),
    .B(_12003_),
    .X(_12004_));
 sky130_fd_sc_hd__xnor2_2 _14882_ (.A(_12001_),
    .B(_12004_),
    .Y(_12005_));
 sky130_fd_sc_hd__nand2_2 _14883_ (.A(\systolic_inst.A_outs[14][2] ),
    .B(\systolic_inst.B_outs[14][5] ),
    .Y(_12006_));
 sky130_fd_sc_hd__and2b_2 _14884_ (.A_N(\systolic_inst.A_outs[14][0] ),
    .B(\systolic_inst.B_outs[14][7] ),
    .X(_12007_));
 sky130_fd_sc_hd__and3_2 _14885_ (.A(\systolic_inst.A_outs[14][1] ),
    .B(\systolic_inst.B_outs[14][6] ),
    .C(_12007_),
    .X(_12008_));
 sky130_fd_sc_hd__xnor2_2 _14886_ (.A(_11975_),
    .B(_12007_),
    .Y(_12009_));
 sky130_fd_sc_hd__xnor2_2 _14887_ (.A(_12006_),
    .B(_12009_),
    .Y(_12010_));
 sky130_fd_sc_hd__xnor2_2 _14888_ (.A(_11976_),
    .B(_12010_),
    .Y(_12011_));
 sky130_fd_sc_hd__nor2_2 _14889_ (.A(_12005_),
    .B(_12011_),
    .Y(_12012_));
 sky130_fd_sc_hd__xnor2_2 _14890_ (.A(_12005_),
    .B(_12011_),
    .Y(_12013_));
 sky130_fd_sc_hd__or2_2 _14891_ (.A(_11978_),
    .B(_12013_),
    .X(_12014_));
 sky130_fd_sc_hd__and2_2 _14892_ (.A(_11978_),
    .B(_12013_),
    .X(_12015_));
 sky130_fd_sc_hd__xor2_2 _14893_ (.A(_11978_),
    .B(_12013_),
    .X(_12016_));
 sky130_fd_sc_hd__xnor2_2 _14894_ (.A(_12000_),
    .B(_12016_),
    .Y(_12017_));
 sky130_fd_sc_hd__o32a_2 _14895_ (.A1(_11966_),
    .A2(_11967_),
    .A3(_11980_),
    .B1(_11979_),
    .B2(_11948_),
    .X(_12018_));
 sky130_fd_sc_hd__nand2b_2 _14896_ (.A_N(_12018_),
    .B(_12017_),
    .Y(_12019_));
 sky130_fd_sc_hd__xnor2_2 _14897_ (.A(_12017_),
    .B(_12018_),
    .Y(_12020_));
 sky130_fd_sc_hd__nand2b_2 _14898_ (.A_N(_11991_),
    .B(_12020_),
    .Y(_12021_));
 sky130_fd_sc_hd__xnor2_2 _14899_ (.A(_11991_),
    .B(_12020_),
    .Y(_12022_));
 sky130_fd_sc_hd__nand2b_2 _14900_ (.A_N(_11990_),
    .B(_12022_),
    .Y(_12023_));
 sky130_fd_sc_hd__xnor2_2 _14901_ (.A(_11990_),
    .B(_12022_),
    .Y(_12024_));
 sky130_fd_sc_hd__o21ai_2 _14902_ (.A1(_11985_),
    .A2(_11988_),
    .B1(_12024_),
    .Y(_12025_));
 sky130_fd_sc_hd__o31a_2 _14903_ (.A1(_11985_),
    .A2(_11988_),
    .A3(_12024_),
    .B1(\systolic_inst.ce_local ),
    .X(_12026_));
 sky130_fd_sc_hd__a22o_2 _14904_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[7] ),
    .B1(_12025_),
    .B2(_12026_),
    .X(_01033_));
 sky130_fd_sc_hd__a21o_2 _14905_ (.A1(_11963_),
    .A2(_11999_),
    .B1(_11997_),
    .X(_12027_));
 sky130_fd_sc_hd__a21bo_2 _14906_ (.A1(\systolic_inst.B_outs[14][7] ),
    .A2(_11993_),
    .B1_N(_11994_),
    .X(_12028_));
 sky130_fd_sc_hd__o21bai_2 _14907_ (.A1(_12001_),
    .A2(_12003_),
    .B1_N(_12002_),
    .Y(_12029_));
 sky130_fd_sc_hd__o21a_2 _14908_ (.A1(\systolic_inst.B_outs[14][0] ),
    .A2(\systolic_inst.B_outs[14][1] ),
    .B1(\systolic_inst.A_outs[14][7] ),
    .X(_12030_));
 sky130_fd_sc_hd__o21ai_2 _14909_ (.A1(\systolic_inst.B_outs[14][0] ),
    .A2(\systolic_inst.B_outs[14][1] ),
    .B1(\systolic_inst.A_outs[14][7] ),
    .Y(_12031_));
 sky130_fd_sc_hd__a21o_2 _14910_ (.A1(\systolic_inst.B_outs[14][0] ),
    .A2(\systolic_inst.B_outs[14][1] ),
    .B1(_12031_),
    .X(_12032_));
 sky130_fd_sc_hd__and2b_2 _14911_ (.A_N(_12032_),
    .B(_12029_),
    .X(_12033_));
 sky130_fd_sc_hd__xnor2_2 _14912_ (.A(_12029_),
    .B(_12032_),
    .Y(_12034_));
 sky130_fd_sc_hd__xnor2_2 _14913_ (.A(_12028_),
    .B(_12034_),
    .Y(_12035_));
 sky130_fd_sc_hd__and4_2 _14914_ (.A(\systolic_inst.B_outs[14][3] ),
    .B(\systolic_inst.B_outs[14][4] ),
    .C(\systolic_inst.A_outs[14][4] ),
    .D(\systolic_inst.A_outs[14][5] ),
    .X(_12036_));
 sky130_fd_sc_hd__a22oi_2 _14915_ (.A1(\systolic_inst.B_outs[14][4] ),
    .A2(\systolic_inst.A_outs[14][4] ),
    .B1(\systolic_inst.A_outs[14][5] ),
    .B2(\systolic_inst.B_outs[14][3] ),
    .Y(_12037_));
 sky130_fd_sc_hd__nor2_2 _14916_ (.A(_12036_),
    .B(_12037_),
    .Y(_12038_));
 sky130_fd_sc_hd__nand2_2 _14917_ (.A(\systolic_inst.B_outs[14][2] ),
    .B(\systolic_inst.A_outs[14][6] ),
    .Y(_12039_));
 sky130_fd_sc_hd__xnor2_2 _14918_ (.A(_12038_),
    .B(_12039_),
    .Y(_12040_));
 sky130_fd_sc_hd__nand2_2 _14919_ (.A(\systolic_inst.A_outs[14][3] ),
    .B(\systolic_inst.B_outs[14][5] ),
    .Y(_12041_));
 sky130_fd_sc_hd__and4b_2 _14920_ (.A_N(\systolic_inst.A_outs[14][1] ),
    .B(\systolic_inst.A_outs[14][2] ),
    .C(\systolic_inst.B_outs[14][6] ),
    .D(\systolic_inst.B_outs[14][7] ),
    .X(_12042_));
 sky130_fd_sc_hd__o2bb2a_2 _14921_ (.A1_N(\systolic_inst.A_outs[14][2] ),
    .A2_N(\systolic_inst.B_outs[14][6] ),
    .B1(_11264_),
    .B2(\systolic_inst.A_outs[14][1] ),
    .X(_12043_));
 sky130_fd_sc_hd__nor2_2 _14922_ (.A(_12042_),
    .B(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__xnor2_2 _14923_ (.A(_12041_),
    .B(_12044_),
    .Y(_12045_));
 sky130_fd_sc_hd__a31oi_2 _14924_ (.A1(\systolic_inst.A_outs[14][2] ),
    .A2(\systolic_inst.B_outs[14][5] ),
    .A3(_12009_),
    .B1(_12008_),
    .Y(_12046_));
 sky130_fd_sc_hd__nand2b_2 _14925_ (.A_N(_12046_),
    .B(_12045_),
    .Y(_12047_));
 sky130_fd_sc_hd__xnor2_2 _14926_ (.A(_12045_),
    .B(_12046_),
    .Y(_12048_));
 sky130_fd_sc_hd__nand2_2 _14927_ (.A(_12040_),
    .B(_12048_),
    .Y(_12049_));
 sky130_fd_sc_hd__xnor2_2 _14928_ (.A(_12040_),
    .B(_12048_),
    .Y(_12050_));
 sky130_fd_sc_hd__a21oi_2 _14929_ (.A1(_11976_),
    .A2(_12010_),
    .B1(_12012_),
    .Y(_12051_));
 sky130_fd_sc_hd__xnor2_2 _14930_ (.A(_12050_),
    .B(_12051_),
    .Y(_12052_));
 sky130_fd_sc_hd__or2_2 _14931_ (.A(_12035_),
    .B(_12052_),
    .X(_12053_));
 sky130_fd_sc_hd__xor2_2 _14932_ (.A(_12035_),
    .B(_12052_),
    .X(_12054_));
 sky130_fd_sc_hd__o21a_2 _14933_ (.A1(_12000_),
    .A2(_12015_),
    .B1(_12014_),
    .X(_12055_));
 sky130_fd_sc_hd__nand2b_2 _14934_ (.A_N(_12055_),
    .B(_12054_),
    .Y(_12056_));
 sky130_fd_sc_hd__xor2_2 _14935_ (.A(_12054_),
    .B(_12055_),
    .X(_12057_));
 sky130_fd_sc_hd__nand2b_2 _14936_ (.A_N(_12057_),
    .B(_12027_),
    .Y(_12058_));
 sky130_fd_sc_hd__xor2_2 _14937_ (.A(_12027_),
    .B(_12057_),
    .X(_12059_));
 sky130_fd_sc_hd__and2_2 _14938_ (.A(_12019_),
    .B(_12021_),
    .X(_12060_));
 sky130_fd_sc_hd__or2_2 _14939_ (.A(_12059_),
    .B(_12060_),
    .X(_12061_));
 sky130_fd_sc_hd__inv_2 _14940_ (.A(_12061_),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_2 _14941_ (.A(_12059_),
    .B(_12060_),
    .Y(_12063_));
 sky130_fd_sc_hd__and2_2 _14942_ (.A(_12061_),
    .B(_12063_),
    .X(_12064_));
 sky130_fd_sc_hd__and2_2 _14943_ (.A(_12023_),
    .B(_12025_),
    .X(_12065_));
 sky130_fd_sc_hd__and2b_2 _14944_ (.A_N(_12065_),
    .B(_12064_),
    .X(_12066_));
 sky130_fd_sc_hd__nand2b_2 _14945_ (.A_N(_12065_),
    .B(_12064_),
    .Y(_12067_));
 sky130_fd_sc_hd__nand2b_2 _14946_ (.A_N(_12064_),
    .B(_12065_),
    .Y(_12068_));
 sky130_fd_sc_hd__and2_2 _14947_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[8] ),
    .X(_12069_));
 sky130_fd_sc_hd__a31o_2 _14948_ (.A1(\systolic_inst.ce_local ),
    .A2(_12067_),
    .A3(_12068_),
    .B1(_12069_),
    .X(_01034_));
 sky130_fd_sc_hd__a21o_2 _14949_ (.A1(_12028_),
    .A2(_12034_),
    .B1(_12033_),
    .X(_12070_));
 sky130_fd_sc_hd__o21ba_2 _14950_ (.A1(_12037_),
    .A2(_12039_),
    .B1_N(_12036_),
    .X(_12071_));
 sky130_fd_sc_hd__nor2_2 _14951_ (.A(_12031_),
    .B(_12071_),
    .Y(_12072_));
 sky130_fd_sc_hd__and2_2 _14952_ (.A(_12031_),
    .B(_12071_),
    .X(_12073_));
 sky130_fd_sc_hd__or2_2 _14953_ (.A(_12072_),
    .B(_12073_),
    .X(_12074_));
 sky130_fd_sc_hd__nand2_2 _14954_ (.A(\systolic_inst.B_outs[14][2] ),
    .B(\systolic_inst.A_outs[14][7] ),
    .Y(_12075_));
 sky130_fd_sc_hd__a22oi_2 _14955_ (.A1(\systolic_inst.B_outs[14][4] ),
    .A2(\systolic_inst.A_outs[14][5] ),
    .B1(\systolic_inst.A_outs[14][6] ),
    .B2(\systolic_inst.B_outs[14][3] ),
    .Y(_12076_));
 sky130_fd_sc_hd__and4_2 _14956_ (.A(\systolic_inst.B_outs[14][3] ),
    .B(\systolic_inst.B_outs[14][4] ),
    .C(\systolic_inst.A_outs[14][5] ),
    .D(\systolic_inst.A_outs[14][6] ),
    .X(_12077_));
 sky130_fd_sc_hd__nor2_2 _14957_ (.A(_12076_),
    .B(_12077_),
    .Y(_12078_));
 sky130_fd_sc_hd__xnor2_2 _14958_ (.A(_12075_),
    .B(_12078_),
    .Y(_12079_));
 sky130_fd_sc_hd__nand2_2 _14959_ (.A(\systolic_inst.A_outs[14][4] ),
    .B(\systolic_inst.B_outs[14][5] ),
    .Y(_12080_));
 sky130_fd_sc_hd__and4b_2 _14960_ (.A_N(\systolic_inst.A_outs[14][2] ),
    .B(\systolic_inst.A_outs[14][3] ),
    .C(\systolic_inst.B_outs[14][6] ),
    .D(\systolic_inst.B_outs[14][7] ),
    .X(_12081_));
 sky130_fd_sc_hd__o2bb2a_2 _14961_ (.A1_N(\systolic_inst.A_outs[14][3] ),
    .A2_N(\systolic_inst.B_outs[14][6] ),
    .B1(_11264_),
    .B2(\systolic_inst.A_outs[14][2] ),
    .X(_12082_));
 sky130_fd_sc_hd__nor2_2 _14962_ (.A(_12081_),
    .B(_12082_),
    .Y(_12083_));
 sky130_fd_sc_hd__xnor2_2 _14963_ (.A(_12080_),
    .B(_12083_),
    .Y(_12084_));
 sky130_fd_sc_hd__o21ba_2 _14964_ (.A1(_12041_),
    .A2(_12043_),
    .B1_N(_12042_),
    .X(_12085_));
 sky130_fd_sc_hd__nand2b_2 _14965_ (.A_N(_12085_),
    .B(_12084_),
    .Y(_12086_));
 sky130_fd_sc_hd__xnor2_2 _14966_ (.A(_12084_),
    .B(_12085_),
    .Y(_12087_));
 sky130_fd_sc_hd__xnor2_2 _14967_ (.A(_12079_),
    .B(_12087_),
    .Y(_12088_));
 sky130_fd_sc_hd__a21o_2 _14968_ (.A1(_12047_),
    .A2(_12049_),
    .B1(_12088_),
    .X(_12089_));
 sky130_fd_sc_hd__nand3_2 _14969_ (.A(_12047_),
    .B(_12049_),
    .C(_12088_),
    .Y(_12090_));
 sky130_fd_sc_hd__nand2_2 _14970_ (.A(_12089_),
    .B(_12090_),
    .Y(_12091_));
 sky130_fd_sc_hd__xor2_2 _14971_ (.A(_12074_),
    .B(_12091_),
    .X(_12092_));
 sky130_fd_sc_hd__o21a_2 _14972_ (.A1(_12050_),
    .A2(_12051_),
    .B1(_12053_),
    .X(_12093_));
 sky130_fd_sc_hd__nand2b_2 _14973_ (.A_N(_12093_),
    .B(_12092_),
    .Y(_12094_));
 sky130_fd_sc_hd__xnor2_2 _14974_ (.A(_12092_),
    .B(_12093_),
    .Y(_12095_));
 sky130_fd_sc_hd__xnor2_2 _14975_ (.A(_12070_),
    .B(_12095_),
    .Y(_12096_));
 sky130_fd_sc_hd__and3_2 _14976_ (.A(_12056_),
    .B(_12058_),
    .C(_12096_),
    .X(_12097_));
 sky130_fd_sc_hd__inv_2 _14977_ (.A(_12097_),
    .Y(_12098_));
 sky130_fd_sc_hd__a21o_2 _14978_ (.A1(_12056_),
    .A2(_12058_),
    .B1(_12096_),
    .X(_12099_));
 sky130_fd_sc_hd__inv_2 _14979_ (.A(_12099_),
    .Y(_12100_));
 sky130_fd_sc_hd__nand2_2 _14980_ (.A(_12098_),
    .B(_12099_),
    .Y(_12101_));
 sky130_fd_sc_hd__a21oi_2 _14981_ (.A1(_12061_),
    .A2(_12067_),
    .B1(_12101_),
    .Y(_12102_));
 sky130_fd_sc_hd__a31o_2 _14982_ (.A1(_12061_),
    .A2(_12067_),
    .A3(_12101_),
    .B1(_11258_),
    .X(_12103_));
 sky130_fd_sc_hd__a2bb2o_2 _14983_ (.A1_N(_12103_),
    .A2_N(_12102_),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[9] ),
    .B2(_11258_),
    .X(_01035_));
 sky130_fd_sc_hd__o21ba_2 _14984_ (.A1(_12075_),
    .A2(_12076_),
    .B1_N(_12077_),
    .X(_12104_));
 sky130_fd_sc_hd__nor2_2 _14985_ (.A(_12031_),
    .B(_12104_),
    .Y(_12105_));
 sky130_fd_sc_hd__and2_2 _14986_ (.A(_12031_),
    .B(_12104_),
    .X(_12106_));
 sky130_fd_sc_hd__or2_2 _14987_ (.A(_12105_),
    .B(_12106_),
    .X(_12107_));
 sky130_fd_sc_hd__a22o_2 _14988_ (.A1(\systolic_inst.B_outs[14][4] ),
    .A2(\systolic_inst.A_outs[14][6] ),
    .B1(\systolic_inst.A_outs[14][7] ),
    .B2(\systolic_inst.B_outs[14][3] ),
    .X(_12108_));
 sky130_fd_sc_hd__and3_2 _14989_ (.A(\systolic_inst.B_outs[14][3] ),
    .B(\systolic_inst.B_outs[14][4] ),
    .C(\systolic_inst.A_outs[14][7] ),
    .X(_12109_));
 sky130_fd_sc_hd__a21bo_2 _14990_ (.A1(\systolic_inst.A_outs[14][6] ),
    .A2(_12109_),
    .B1_N(_12108_),
    .X(_12110_));
 sky130_fd_sc_hd__xor2_2 _14991_ (.A(_12075_),
    .B(_12110_),
    .X(_12111_));
 sky130_fd_sc_hd__nand2_2 _14992_ (.A(\systolic_inst.B_outs[14][5] ),
    .B(\systolic_inst.A_outs[14][5] ),
    .Y(_12112_));
 sky130_fd_sc_hd__and4b_2 _14993_ (.A_N(\systolic_inst.A_outs[14][3] ),
    .B(\systolic_inst.A_outs[14][4] ),
    .C(\systolic_inst.B_outs[14][6] ),
    .D(\systolic_inst.B_outs[14][7] ),
    .X(_12113_));
 sky130_fd_sc_hd__o2bb2a_2 _14994_ (.A1_N(\systolic_inst.A_outs[14][4] ),
    .A2_N(\systolic_inst.B_outs[14][6] ),
    .B1(_11264_),
    .B2(\systolic_inst.A_outs[14][3] ),
    .X(_12114_));
 sky130_fd_sc_hd__nor2_2 _14995_ (.A(_12113_),
    .B(_12114_),
    .Y(_12115_));
 sky130_fd_sc_hd__xnor2_2 _14996_ (.A(_12112_),
    .B(_12115_),
    .Y(_12116_));
 sky130_fd_sc_hd__o21ba_2 _14997_ (.A1(_12080_),
    .A2(_12082_),
    .B1_N(_12081_),
    .X(_12117_));
 sky130_fd_sc_hd__nand2b_2 _14998_ (.A_N(_12117_),
    .B(_12116_),
    .Y(_12118_));
 sky130_fd_sc_hd__xnor2_2 _14999_ (.A(_12116_),
    .B(_12117_),
    .Y(_12119_));
 sky130_fd_sc_hd__nand2_2 _15000_ (.A(_12111_),
    .B(_12119_),
    .Y(_12120_));
 sky130_fd_sc_hd__or2_2 _15001_ (.A(_12111_),
    .B(_12119_),
    .X(_12121_));
 sky130_fd_sc_hd__nand2_2 _15002_ (.A(_12120_),
    .B(_12121_),
    .Y(_12122_));
 sky130_fd_sc_hd__a21bo_2 _15003_ (.A1(_12079_),
    .A2(_12087_),
    .B1_N(_12086_),
    .X(_12123_));
 sky130_fd_sc_hd__nand2b_2 _15004_ (.A_N(_12122_),
    .B(_12123_),
    .Y(_12124_));
 sky130_fd_sc_hd__xor2_2 _15005_ (.A(_12122_),
    .B(_12123_),
    .X(_12125_));
 sky130_fd_sc_hd__xor2_2 _15006_ (.A(_12107_),
    .B(_12125_),
    .X(_12126_));
 sky130_fd_sc_hd__o21a_2 _15007_ (.A1(_12074_),
    .A2(_12091_),
    .B1(_12089_),
    .X(_12127_));
 sky130_fd_sc_hd__nand2b_2 _15008_ (.A_N(_12127_),
    .B(_12126_),
    .Y(_12128_));
 sky130_fd_sc_hd__xnor2_2 _15009_ (.A(_12126_),
    .B(_12127_),
    .Y(_12129_));
 sky130_fd_sc_hd__nand2_2 _15010_ (.A(_12072_),
    .B(_12129_),
    .Y(_12130_));
 sky130_fd_sc_hd__or2_2 _15011_ (.A(_12072_),
    .B(_12129_),
    .X(_12131_));
 sky130_fd_sc_hd__nand2_2 _15012_ (.A(_12130_),
    .B(_12131_),
    .Y(_12132_));
 sky130_fd_sc_hd__a21boi_2 _15013_ (.A1(_12070_),
    .A2(_12095_),
    .B1_N(_12094_),
    .Y(_12133_));
 sky130_fd_sc_hd__nor2_2 _15014_ (.A(_12132_),
    .B(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__xor2_2 _15015_ (.A(_12132_),
    .B(_12133_),
    .X(_12135_));
 sky130_fd_sc_hd__a31o_2 _15016_ (.A1(_12061_),
    .A2(_12067_),
    .A3(_12099_),
    .B1(_12097_),
    .X(_12136_));
 sky130_fd_sc_hd__and2b_2 _15017_ (.A_N(_12135_),
    .B(_12136_),
    .X(_12137_));
 sky130_fd_sc_hd__o311a_2 _15018_ (.A1(_12062_),
    .A2(_12066_),
    .A3(_12100_),
    .B1(_12135_),
    .C1(_12098_),
    .X(_12138_));
 sky130_fd_sc_hd__nor2_2 _15019_ (.A(_12137_),
    .B(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__mux2_1 _15020_ (.A0(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[10] ),
    .A1(_12139_),
    .S(\systolic_inst.ce_local ),
    .X(_01036_));
 sky130_fd_sc_hd__o2bb2a_2 _15021_ (.A1_N(\systolic_inst.A_outs[14][6] ),
    .A2_N(_12109_),
    .B1(_12110_),
    .B2(_12075_),
    .X(_12140_));
 sky130_fd_sc_hd__or2_2 _15022_ (.A(_12031_),
    .B(_12140_),
    .X(_12141_));
 sky130_fd_sc_hd__nand2_2 _15023_ (.A(_12031_),
    .B(_12140_),
    .Y(_12142_));
 sky130_fd_sc_hd__nand2_2 _15024_ (.A(_12141_),
    .B(_12142_),
    .Y(_12143_));
 sky130_fd_sc_hd__or2_2 _15025_ (.A(\systolic_inst.B_outs[14][3] ),
    .B(\systolic_inst.B_outs[14][4] ),
    .X(_12144_));
 sky130_fd_sc_hd__and3b_2 _15026_ (.A_N(_12109_),
    .B(_12144_),
    .C(\systolic_inst.A_outs[14][7] ),
    .X(_12145_));
 sky130_fd_sc_hd__xnor2_2 _15027_ (.A(_12075_),
    .B(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__nand2_2 _15028_ (.A(\systolic_inst.B_outs[14][5] ),
    .B(\systolic_inst.A_outs[14][6] ),
    .Y(_12147_));
 sky130_fd_sc_hd__and4b_2 _15029_ (.A_N(\systolic_inst.A_outs[14][4] ),
    .B(\systolic_inst.A_outs[14][5] ),
    .C(\systolic_inst.B_outs[14][6] ),
    .D(\systolic_inst.B_outs[14][7] ),
    .X(_12148_));
 sky130_fd_sc_hd__o2bb2a_2 _15030_ (.A1_N(\systolic_inst.A_outs[14][5] ),
    .A2_N(\systolic_inst.B_outs[14][6] ),
    .B1(_11264_),
    .B2(\systolic_inst.A_outs[14][4] ),
    .X(_12149_));
 sky130_fd_sc_hd__nor2_2 _15031_ (.A(_12148_),
    .B(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__xnor2_2 _15032_ (.A(_12147_),
    .B(_12150_),
    .Y(_12151_));
 sky130_fd_sc_hd__o21ba_2 _15033_ (.A1(_12112_),
    .A2(_12114_),
    .B1_N(_12113_),
    .X(_12152_));
 sky130_fd_sc_hd__nand2b_2 _15034_ (.A_N(_12152_),
    .B(_12151_),
    .Y(_12153_));
 sky130_fd_sc_hd__xnor2_2 _15035_ (.A(_12151_),
    .B(_12152_),
    .Y(_12154_));
 sky130_fd_sc_hd__nand2_2 _15036_ (.A(_12146_),
    .B(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__xnor2_2 _15037_ (.A(_12146_),
    .B(_12154_),
    .Y(_12156_));
 sky130_fd_sc_hd__a21o_2 _15038_ (.A1(_12118_),
    .A2(_12120_),
    .B1(_12156_),
    .X(_12157_));
 sky130_fd_sc_hd__nand3_2 _15039_ (.A(_12118_),
    .B(_12120_),
    .C(_12156_),
    .Y(_12158_));
 sky130_fd_sc_hd__nand2_2 _15040_ (.A(_12157_),
    .B(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__xor2_2 _15041_ (.A(_12143_),
    .B(_12159_),
    .X(_12160_));
 sky130_fd_sc_hd__o21a_2 _15042_ (.A1(_12107_),
    .A2(_12125_),
    .B1(_12124_),
    .X(_12161_));
 sky130_fd_sc_hd__and2b_2 _15043_ (.A_N(_12161_),
    .B(_12160_),
    .X(_12162_));
 sky130_fd_sc_hd__and2b_2 _15044_ (.A_N(_12160_),
    .B(_12161_),
    .X(_12163_));
 sky130_fd_sc_hd__nor2_2 _15045_ (.A(_12162_),
    .B(_12163_),
    .Y(_12164_));
 sky130_fd_sc_hd__xnor2_2 _15046_ (.A(_12105_),
    .B(_12164_),
    .Y(_12165_));
 sky130_fd_sc_hd__nand3_2 _15047_ (.A(_12128_),
    .B(_12130_),
    .C(_12165_),
    .Y(_12166_));
 sky130_fd_sc_hd__inv_2 _15048_ (.A(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__a21oi_2 _15049_ (.A1(_12128_),
    .A2(_12130_),
    .B1(_12165_),
    .Y(_12168_));
 sky130_fd_sc_hd__nor2_2 _15050_ (.A(_12167_),
    .B(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__or3_2 _15051_ (.A(_12134_),
    .B(_12138_),
    .C(_12169_),
    .X(_12170_));
 sky130_fd_sc_hd__o21ai_2 _15052_ (.A1(_12134_),
    .A2(_12138_),
    .B1(_12169_),
    .Y(_12171_));
 sky130_fd_sc_hd__and2_2 _15053_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[11] ),
    .X(_12172_));
 sky130_fd_sc_hd__a31o_2 _15054_ (.A1(\systolic_inst.ce_local ),
    .A2(_12170_),
    .A3(_12171_),
    .B1(_12172_),
    .X(_01037_));
 sky130_fd_sc_hd__a31o_2 _15055_ (.A1(\systolic_inst.B_outs[14][2] ),
    .A2(\systolic_inst.A_outs[14][7] ),
    .A3(_12144_),
    .B1(_12109_),
    .X(_12173_));
 sky130_fd_sc_hd__or2_2 _15056_ (.A(_12030_),
    .B(_12173_),
    .X(_12174_));
 sky130_fd_sc_hd__nand2_2 _15057_ (.A(_12030_),
    .B(_12173_),
    .Y(_12175_));
 sky130_fd_sc_hd__nand2_2 _15058_ (.A(_12174_),
    .B(_12175_),
    .Y(_12176_));
 sky130_fd_sc_hd__inv_2 _15059_ (.A(_12176_),
    .Y(_12177_));
 sky130_fd_sc_hd__o2bb2a_2 _15060_ (.A1_N(\systolic_inst.B_outs[14][6] ),
    .A2_N(\systolic_inst.A_outs[14][6] ),
    .B1(_11264_),
    .B2(\systolic_inst.A_outs[14][5] ),
    .X(_12178_));
 sky130_fd_sc_hd__and4b_2 _15061_ (.A_N(\systolic_inst.A_outs[14][5] ),
    .B(\systolic_inst.B_outs[14][6] ),
    .C(\systolic_inst.A_outs[14][6] ),
    .D(\systolic_inst.B_outs[14][7] ),
    .X(_12179_));
 sky130_fd_sc_hd__nor2_2 _15062_ (.A(_12178_),
    .B(_12179_),
    .Y(_12180_));
 sky130_fd_sc_hd__nand2_2 _15063_ (.A(\systolic_inst.B_outs[14][5] ),
    .B(\systolic_inst.A_outs[14][7] ),
    .Y(_12181_));
 sky130_fd_sc_hd__and3_2 _15064_ (.A(\systolic_inst.B_outs[14][5] ),
    .B(\systolic_inst.A_outs[14][7] ),
    .C(_12180_),
    .X(_12182_));
 sky130_fd_sc_hd__xnor2_2 _15065_ (.A(_12180_),
    .B(_12181_),
    .Y(_12183_));
 sky130_fd_sc_hd__o21ba_2 _15066_ (.A1(_12147_),
    .A2(_12149_),
    .B1_N(_12148_),
    .X(_12184_));
 sky130_fd_sc_hd__nand2b_2 _15067_ (.A_N(_12184_),
    .B(_12183_),
    .Y(_12185_));
 sky130_fd_sc_hd__xnor2_2 _15068_ (.A(_12183_),
    .B(_12184_),
    .Y(_12186_));
 sky130_fd_sc_hd__xnor2_2 _15069_ (.A(_12146_),
    .B(_12186_),
    .Y(_12187_));
 sky130_fd_sc_hd__a21o_2 _15070_ (.A1(_12153_),
    .A2(_12155_),
    .B1(_12187_),
    .X(_12188_));
 sky130_fd_sc_hd__nand3_2 _15071_ (.A(_12153_),
    .B(_12155_),
    .C(_12187_),
    .Y(_12189_));
 sky130_fd_sc_hd__nand2_2 _15072_ (.A(_12188_),
    .B(_12189_),
    .Y(_12190_));
 sky130_fd_sc_hd__xnor2_2 _15073_ (.A(_12177_),
    .B(_12190_),
    .Y(_12191_));
 sky130_fd_sc_hd__o21a_2 _15074_ (.A1(_12143_),
    .A2(_12159_),
    .B1(_12157_),
    .X(_12192_));
 sky130_fd_sc_hd__and2b_2 _15075_ (.A_N(_12192_),
    .B(_12191_),
    .X(_12193_));
 sky130_fd_sc_hd__and2b_2 _15076_ (.A_N(_12191_),
    .B(_12192_),
    .X(_12194_));
 sky130_fd_sc_hd__nor2_2 _15077_ (.A(_12193_),
    .B(_12194_),
    .Y(_12195_));
 sky130_fd_sc_hd__and2b_2 _15078_ (.A_N(_12141_),
    .B(_12195_),
    .X(_12196_));
 sky130_fd_sc_hd__xor2_2 _15079_ (.A(_12141_),
    .B(_12195_),
    .X(_12197_));
 sky130_fd_sc_hd__a21oi_2 _15080_ (.A1(_12105_),
    .A2(_12164_),
    .B1(_12162_),
    .Y(_12198_));
 sky130_fd_sc_hd__nor2_2 _15081_ (.A(_12197_),
    .B(_12198_),
    .Y(_12199_));
 sky130_fd_sc_hd__and2_2 _15082_ (.A(_12197_),
    .B(_12198_),
    .X(_12200_));
 sky130_fd_sc_hd__nor2_2 _15083_ (.A(_12199_),
    .B(_12200_),
    .Y(_12201_));
 sky130_fd_sc_hd__o31a_2 _15084_ (.A1(_12134_),
    .A2(_12138_),
    .A3(_12168_),
    .B1(_12166_),
    .X(_12202_));
 sky130_fd_sc_hd__o311a_2 _15085_ (.A1(_12134_),
    .A2(_12138_),
    .A3(_12168_),
    .B1(_12201_),
    .C1(_12166_),
    .X(_12203_));
 sky130_fd_sc_hd__xor2_2 _15086_ (.A(_12201_),
    .B(_12202_),
    .X(_12204_));
 sky130_fd_sc_hd__mux2_1 _15087_ (.A0(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[12] ),
    .A1(_12204_),
    .S(\systolic_inst.ce_local ),
    .X(_01038_));
 sky130_fd_sc_hd__nand2_2 _15088_ (.A(\systolic_inst.B_outs[14][6] ),
    .B(\systolic_inst.A_outs[14][7] ),
    .Y(_12205_));
 sky130_fd_sc_hd__or2_2 _15089_ (.A(\systolic_inst.A_outs[14][6] ),
    .B(_11264_),
    .X(_12206_));
 sky130_fd_sc_hd__and2_2 _15090_ (.A(_12205_),
    .B(_12206_),
    .X(_12207_));
 sky130_fd_sc_hd__nor2_2 _15091_ (.A(_12205_),
    .B(_12206_),
    .Y(_12208_));
 sky130_fd_sc_hd__nor2_2 _15092_ (.A(_12207_),
    .B(_12208_),
    .Y(_12209_));
 sky130_fd_sc_hd__xnor2_2 _15093_ (.A(_12181_),
    .B(_12209_),
    .Y(_12210_));
 sky130_fd_sc_hd__o21ai_2 _15094_ (.A1(_12179_),
    .A2(_12182_),
    .B1(_12210_),
    .Y(_12211_));
 sky130_fd_sc_hd__or3_2 _15095_ (.A(_12179_),
    .B(_12182_),
    .C(_12210_),
    .X(_12212_));
 sky130_fd_sc_hd__and2_2 _15096_ (.A(_12211_),
    .B(_12212_),
    .X(_12213_));
 sky130_fd_sc_hd__nand2_2 _15097_ (.A(_12146_),
    .B(_12213_),
    .Y(_12214_));
 sky130_fd_sc_hd__or2_2 _15098_ (.A(_12146_),
    .B(_12213_),
    .X(_12215_));
 sky130_fd_sc_hd__nand2_2 _15099_ (.A(_12214_),
    .B(_12215_),
    .Y(_12216_));
 sky130_fd_sc_hd__a21bo_2 _15100_ (.A1(_12146_),
    .A2(_12186_),
    .B1_N(_12185_),
    .X(_12217_));
 sky130_fd_sc_hd__nand2b_2 _15101_ (.A_N(_12216_),
    .B(_12217_),
    .Y(_12218_));
 sky130_fd_sc_hd__xor2_2 _15102_ (.A(_12216_),
    .B(_12217_),
    .X(_12219_));
 sky130_fd_sc_hd__xnor2_2 _15103_ (.A(_12177_),
    .B(_12219_),
    .Y(_12220_));
 sky130_fd_sc_hd__o21a_2 _15104_ (.A1(_12176_),
    .A2(_12190_),
    .B1(_12188_),
    .X(_12221_));
 sky130_fd_sc_hd__and2b_2 _15105_ (.A_N(_12221_),
    .B(_12220_),
    .X(_12222_));
 sky130_fd_sc_hd__and2b_2 _15106_ (.A_N(_12220_),
    .B(_12221_),
    .X(_12223_));
 sky130_fd_sc_hd__nor2_2 _15107_ (.A(_12222_),
    .B(_12223_),
    .Y(_12224_));
 sky130_fd_sc_hd__xnor2_2 _15108_ (.A(_12175_),
    .B(_12224_),
    .Y(_12225_));
 sky130_fd_sc_hd__o21a_2 _15109_ (.A1(_12193_),
    .A2(_12196_),
    .B1(_12225_),
    .X(_12226_));
 sky130_fd_sc_hd__or3_2 _15110_ (.A(_12193_),
    .B(_12196_),
    .C(_12225_),
    .X(_12227_));
 sky130_fd_sc_hd__and2b_2 _15111_ (.A_N(_12226_),
    .B(_12227_),
    .X(_12228_));
 sky130_fd_sc_hd__nor2_2 _15112_ (.A(_12199_),
    .B(_12203_),
    .Y(_12229_));
 sky130_fd_sc_hd__xnor2_2 _15113_ (.A(_12228_),
    .B(_12229_),
    .Y(_12230_));
 sky130_fd_sc_hd__mux2_1 _15114_ (.A0(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[13] ),
    .A1(_12230_),
    .S(\systolic_inst.ce_local ),
    .X(_01039_));
 sky130_fd_sc_hd__a31o_2 _15115_ (.A1(\systolic_inst.B_outs[14][5] ),
    .A2(\systolic_inst.A_outs[14][7] ),
    .A3(_12209_),
    .B1(_12208_),
    .X(_12231_));
 sky130_fd_sc_hd__nand3_2 _15116_ (.A(\systolic_inst.B_outs[14][5] ),
    .B(\systolic_inst.B_outs[14][6] ),
    .C(\systolic_inst.A_outs[14][7] ),
    .Y(_12232_));
 sky130_fd_sc_hd__o211a_2 _15117_ (.A1(_11264_),
    .A2(\systolic_inst.A_outs[14][7] ),
    .B1(_12181_),
    .C1(_12205_),
    .X(_12233_));
 sky130_fd_sc_hd__a21oi_2 _15118_ (.A1(_12231_),
    .A2(_12232_),
    .B1(_12233_),
    .Y(_12234_));
 sky130_fd_sc_hd__nor2_2 _15119_ (.A(_12146_),
    .B(_12234_),
    .Y(_12235_));
 sky130_fd_sc_hd__and2_2 _15120_ (.A(_12146_),
    .B(_12234_),
    .X(_12236_));
 sky130_fd_sc_hd__or2_2 _15121_ (.A(_12235_),
    .B(_12236_),
    .X(_12237_));
 sky130_fd_sc_hd__a21oi_2 _15122_ (.A1(_12211_),
    .A2(_12214_),
    .B1(_12237_),
    .Y(_12238_));
 sky130_fd_sc_hd__and3_2 _15123_ (.A(_12211_),
    .B(_12214_),
    .C(_12237_),
    .X(_12239_));
 sky130_fd_sc_hd__nor2_2 _15124_ (.A(_12238_),
    .B(_12239_),
    .Y(_12240_));
 sky130_fd_sc_hd__xnor2_2 _15125_ (.A(_12176_),
    .B(_12240_),
    .Y(_12241_));
 sky130_fd_sc_hd__o21a_2 _15126_ (.A1(_12176_),
    .A2(_12219_),
    .B1(_12218_),
    .X(_12242_));
 sky130_fd_sc_hd__and2b_2 _15127_ (.A_N(_12242_),
    .B(_12241_),
    .X(_12243_));
 sky130_fd_sc_hd__and2b_2 _15128_ (.A_N(_12241_),
    .B(_12242_),
    .X(_12244_));
 sky130_fd_sc_hd__nor2_2 _15129_ (.A(_12243_),
    .B(_12244_),
    .Y(_12245_));
 sky130_fd_sc_hd__xnor2_2 _15130_ (.A(_12175_),
    .B(_12245_),
    .Y(_12246_));
 sky130_fd_sc_hd__o21ba_2 _15131_ (.A1(_12175_),
    .A2(_12223_),
    .B1_N(_12222_),
    .X(_12247_));
 sky130_fd_sc_hd__and2b_2 _15132_ (.A_N(_12247_),
    .B(_12246_),
    .X(_12248_));
 sky130_fd_sc_hd__xnor2_2 _15133_ (.A(_12246_),
    .B(_12247_),
    .Y(_12249_));
 sky130_fd_sc_hd__o31a_2 _15134_ (.A1(_12199_),
    .A2(_12203_),
    .A3(_12226_),
    .B1(_12227_),
    .X(_12250_));
 sky130_fd_sc_hd__or2_2 _15135_ (.A(_12249_),
    .B(_12250_),
    .X(_12251_));
 sky130_fd_sc_hd__o311a_2 _15136_ (.A1(_12199_),
    .A2(_12203_),
    .A3(_12226_),
    .B1(_12227_),
    .C1(_12249_),
    .X(_12252_));
 sky130_fd_sc_hd__nor2_2 _15137_ (.A(_11258_),
    .B(_12252_),
    .Y(_12253_));
 sky130_fd_sc_hd__a22o_2 _15138_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[14] ),
    .B1(_12251_),
    .B2(_12253_),
    .X(_01040_));
 sky130_fd_sc_hd__a31o_2 _15139_ (.A1(_12030_),
    .A2(_12173_),
    .A3(_12245_),
    .B1(_12243_),
    .X(_12254_));
 sky130_fd_sc_hd__a21oi_2 _15140_ (.A1(_12177_),
    .A2(_12240_),
    .B1(_12238_),
    .Y(_12255_));
 sky130_fd_sc_hd__xnor2_2 _15141_ (.A(_12174_),
    .B(_12235_),
    .Y(_12256_));
 sky130_fd_sc_hd__xnor2_2 _15142_ (.A(_12255_),
    .B(_12256_),
    .Y(_12257_));
 sky130_fd_sc_hd__xnor2_2 _15143_ (.A(_12254_),
    .B(_12257_),
    .Y(_12258_));
 sky130_fd_sc_hd__or3_2 _15144_ (.A(_11258_),
    .B(_12248_),
    .C(_12258_),
    .X(_12259_));
 sky130_fd_sc_hd__a2bb2o_2 _15145_ (.A1_N(_12259_),
    .A2_N(_12252_),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B2(_11258_),
    .X(_01041_));
 sky130_fd_sc_hd__a21o_2 _15146_ (.A1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[14][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_12260_));
 sky130_fd_sc_hd__a21oi_2 _15147_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[14][0] ),
    .Y(_12261_));
 sky130_fd_sc_hd__a21oi_2 _15148_ (.A1(\systolic_inst.ce_local ),
    .A2(_12260_),
    .B1(_12261_),
    .Y(_01042_));
 sky130_fd_sc_hd__and2_2 _15149_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[14][1] ),
    .X(_12262_));
 sky130_fd_sc_hd__nand2_2 _15150_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[14][1] ),
    .Y(_12263_));
 sky130_fd_sc_hd__or2_2 _15151_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[14][1] ),
    .X(_12264_));
 sky130_fd_sc_hd__and4_2 _15152_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[14][0] ),
    .C(_12263_),
    .D(_12264_),
    .X(_12265_));
 sky130_fd_sc_hd__inv_2 _15153_ (.A(_12265_),
    .Y(_12266_));
 sky130_fd_sc_hd__a22o_2 _15154_ (.A1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[14][0] ),
    .B1(_12263_),
    .B2(_12264_),
    .X(_12267_));
 sky130_fd_sc_hd__a32o_2 _15155_ (.A1(_11712_),
    .A2(_12266_),
    .A3(_12267_),
    .B1(\systolic_inst.acc_wires[14][1] ),
    .B2(_11258_),
    .X(_01043_));
 sky130_fd_sc_hd__and2_2 _15156_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[14][2] ),
    .X(_12268_));
 sky130_fd_sc_hd__nand2_2 _15157_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[14][2] ),
    .Y(_12269_));
 sky130_fd_sc_hd__or2_2 _15158_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[14][2] ),
    .X(_12270_));
 sky130_fd_sc_hd__a211o_2 _15159_ (.A1(_12269_),
    .A2(_12270_),
    .B1(_12262_),
    .C1(_12265_),
    .X(_12271_));
 sky130_fd_sc_hd__o211a_2 _15160_ (.A1(_12262_),
    .A2(_12265_),
    .B1(_12269_),
    .C1(_12270_),
    .X(_12272_));
 sky130_fd_sc_hd__inv_2 _15161_ (.A(_12272_),
    .Y(_12273_));
 sky130_fd_sc_hd__a32o_2 _15162_ (.A1(_11712_),
    .A2(_12271_),
    .A3(_12273_),
    .B1(\systolic_inst.acc_wires[14][2] ),
    .B2(_11258_),
    .X(_01044_));
 sky130_fd_sc_hd__and2_2 _15163_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[14][3] ),
    .X(_12274_));
 sky130_fd_sc_hd__nand2_2 _15164_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[14][3] ),
    .Y(_12275_));
 sky130_fd_sc_hd__or2_2 _15165_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[14][3] ),
    .X(_12276_));
 sky130_fd_sc_hd__a211o_2 _15166_ (.A1(_12275_),
    .A2(_12276_),
    .B1(_12268_),
    .C1(_12272_),
    .X(_12277_));
 sky130_fd_sc_hd__o211a_2 _15167_ (.A1(_12268_),
    .A2(_12272_),
    .B1(_12275_),
    .C1(_12276_),
    .X(_12278_));
 sky130_fd_sc_hd__inv_2 _15168_ (.A(_12278_),
    .Y(_12279_));
 sky130_fd_sc_hd__a32o_2 _15169_ (.A1(_11712_),
    .A2(_12277_),
    .A3(_12279_),
    .B1(\systolic_inst.acc_wires[14][3] ),
    .B2(_11258_),
    .X(_01045_));
 sky130_fd_sc_hd__and2_2 _15170_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[14][4] ),
    .X(_12280_));
 sky130_fd_sc_hd__nand2_2 _15171_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[14][4] ),
    .Y(_12281_));
 sky130_fd_sc_hd__or2_2 _15172_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[14][4] ),
    .X(_12282_));
 sky130_fd_sc_hd__a211o_2 _15173_ (.A1(_12281_),
    .A2(_12282_),
    .B1(_12274_),
    .C1(_12278_),
    .X(_12283_));
 sky130_fd_sc_hd__o211a_2 _15174_ (.A1(_12274_),
    .A2(_12278_),
    .B1(_12281_),
    .C1(_12282_),
    .X(_12284_));
 sky130_fd_sc_hd__inv_2 _15175_ (.A(_12284_),
    .Y(_12285_));
 sky130_fd_sc_hd__a32o_2 _15176_ (.A1(_11712_),
    .A2(_12283_),
    .A3(_12285_),
    .B1(\systolic_inst.acc_wires[14][4] ),
    .B2(_11258_),
    .X(_01046_));
 sky130_fd_sc_hd__and2_2 _15177_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[14][5] ),
    .X(_12286_));
 sky130_fd_sc_hd__nand2_2 _15178_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[14][5] ),
    .Y(_12287_));
 sky130_fd_sc_hd__or2_2 _15179_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[14][5] ),
    .X(_12288_));
 sky130_fd_sc_hd__a211o_2 _15180_ (.A1(_12287_),
    .A2(_12288_),
    .B1(_12280_),
    .C1(_12284_),
    .X(_12289_));
 sky130_fd_sc_hd__o211a_2 _15181_ (.A1(_12280_),
    .A2(_12284_),
    .B1(_12287_),
    .C1(_12288_),
    .X(_12290_));
 sky130_fd_sc_hd__inv_2 _15182_ (.A(_12290_),
    .Y(_12291_));
 sky130_fd_sc_hd__a32o_2 _15183_ (.A1(_11712_),
    .A2(_12289_),
    .A3(_12291_),
    .B1(\systolic_inst.acc_wires[14][5] ),
    .B2(_11258_),
    .X(_01047_));
 sky130_fd_sc_hd__and2_2 _15184_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[14][6] ),
    .X(_12292_));
 sky130_fd_sc_hd__nand2_2 _15185_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[14][6] ),
    .Y(_12293_));
 sky130_fd_sc_hd__or2_2 _15186_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[14][6] ),
    .X(_12294_));
 sky130_fd_sc_hd__a211o_2 _15187_ (.A1(_12293_),
    .A2(_12294_),
    .B1(_12286_),
    .C1(_12290_),
    .X(_12295_));
 sky130_fd_sc_hd__o211a_2 _15188_ (.A1(_12286_),
    .A2(_12290_),
    .B1(_12293_),
    .C1(_12294_),
    .X(_12296_));
 sky130_fd_sc_hd__inv_2 _15189_ (.A(_12296_),
    .Y(_12297_));
 sky130_fd_sc_hd__a32o_2 _15190_ (.A1(_11712_),
    .A2(_12295_),
    .A3(_12297_),
    .B1(\systolic_inst.acc_wires[14][6] ),
    .B2(_11258_),
    .X(_01048_));
 sky130_fd_sc_hd__nand2_2 _15191_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[14][7] ),
    .Y(_12298_));
 sky130_fd_sc_hd__or2_2 _15192_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[14][7] ),
    .X(_12299_));
 sky130_fd_sc_hd__a211o_2 _15193_ (.A1(_12298_),
    .A2(_12299_),
    .B1(_12292_),
    .C1(_12296_),
    .X(_12300_));
 sky130_fd_sc_hd__o211ai_2 _15194_ (.A1(_12292_),
    .A2(_12296_),
    .B1(_12298_),
    .C1(_12299_),
    .Y(_12301_));
 sky130_fd_sc_hd__a32o_2 _15195_ (.A1(_11712_),
    .A2(_12300_),
    .A3(_12301_),
    .B1(\systolic_inst.acc_wires[14][7] ),
    .B2(_11258_),
    .X(_01049_));
 sky130_fd_sc_hd__and2_2 _15196_ (.A(_12298_),
    .B(_12301_),
    .X(_12302_));
 sky130_fd_sc_hd__nand2_2 _15197_ (.A(_12298_),
    .B(_12301_),
    .Y(_12303_));
 sky130_fd_sc_hd__nor2_2 _15198_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[14][8] ),
    .Y(_12304_));
 sky130_fd_sc_hd__and2_2 _15199_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[14][8] ),
    .X(_12305_));
 sky130_fd_sc_hd__nor2_2 _15200_ (.A(_12304_),
    .B(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__xnor2_2 _15201_ (.A(_12302_),
    .B(_12306_),
    .Y(_12307_));
 sky130_fd_sc_hd__a22o_2 _15202_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][8] ),
    .B1(_11712_),
    .B2(_12307_),
    .X(_01050_));
 sky130_fd_sc_hd__xor2_2 _15203_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[14][9] ),
    .X(_12308_));
 sky130_fd_sc_hd__a211o_2 _15204_ (.A1(_12303_),
    .A2(_12306_),
    .B1(_12308_),
    .C1(_12305_),
    .X(_12309_));
 sky130_fd_sc_hd__nand2_2 _15205_ (.A(_12306_),
    .B(_12308_),
    .Y(_12310_));
 sky130_fd_sc_hd__or2_2 _15206_ (.A(_12302_),
    .B(_12310_),
    .X(_12311_));
 sky130_fd_sc_hd__and2_2 _15207_ (.A(_12305_),
    .B(_12308_),
    .X(_12312_));
 sky130_fd_sc_hd__nor2_2 _15208_ (.A(_11713_),
    .B(_12312_),
    .Y(_12313_));
 sky130_fd_sc_hd__a32o_2 _15209_ (.A1(_12309_),
    .A2(_12311_),
    .A3(_12313_),
    .B1(\systolic_inst.acc_wires[14][9] ),
    .B2(_11258_),
    .X(_01051_));
 sky130_fd_sc_hd__nand2_2 _15210_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[14][10] ),
    .Y(_12314_));
 sky130_fd_sc_hd__or2_2 _15211_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[14][10] ),
    .X(_12315_));
 sky130_fd_sc_hd__and2_2 _15212_ (.A(_12314_),
    .B(_12315_),
    .X(_12316_));
 sky130_fd_sc_hd__a21oi_2 _15213_ (.A1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[14][9] ),
    .B1(_12312_),
    .Y(_12317_));
 sky130_fd_sc_hd__nand2_2 _15214_ (.A(_12311_),
    .B(_12317_),
    .Y(_12318_));
 sky130_fd_sc_hd__xor2_2 _15215_ (.A(_12316_),
    .B(_12318_),
    .X(_12319_));
 sky130_fd_sc_hd__a22o_2 _15216_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][10] ),
    .B1(_11712_),
    .B2(_12319_),
    .X(_01052_));
 sky130_fd_sc_hd__nor2_2 _15217_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[14][11] ),
    .Y(_12320_));
 sky130_fd_sc_hd__or2_2 _15218_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[14][11] ),
    .X(_12321_));
 sky130_fd_sc_hd__nand2_2 _15219_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[14][11] ),
    .Y(_12322_));
 sky130_fd_sc_hd__nand2_2 _15220_ (.A(_12321_),
    .B(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__a21bo_2 _15221_ (.A1(_12316_),
    .A2(_12318_),
    .B1_N(_12314_),
    .X(_12324_));
 sky130_fd_sc_hd__xnor2_2 _15222_ (.A(_12323_),
    .B(_12324_),
    .Y(_12325_));
 sky130_fd_sc_hd__a22o_2 _15223_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][11] ),
    .B1(_11712_),
    .B2(_12325_),
    .X(_01053_));
 sky130_fd_sc_hd__nand3_2 _15224_ (.A(_12316_),
    .B(_12321_),
    .C(_12322_),
    .Y(_12326_));
 sky130_fd_sc_hd__a211o_2 _15225_ (.A1(_12298_),
    .A2(_12301_),
    .B1(_12310_),
    .C1(_12326_),
    .X(_12327_));
 sky130_fd_sc_hd__o21a_2 _15226_ (.A1(_12314_),
    .A2(_12320_),
    .B1(_12322_),
    .X(_12328_));
 sky130_fd_sc_hd__o211a_2 _15227_ (.A1(_12317_),
    .A2(_12326_),
    .B1(_12327_),
    .C1(_12328_),
    .X(_12329_));
 sky130_fd_sc_hd__xnor2_2 _15228_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[14][12] ),
    .Y(_12330_));
 sky130_fd_sc_hd__inv_2 _15229_ (.A(_12330_),
    .Y(_12331_));
 sky130_fd_sc_hd__nand2_2 _15230_ (.A(_12329_),
    .B(_12330_),
    .Y(_12332_));
 sky130_fd_sc_hd__nor2_2 _15231_ (.A(_12329_),
    .B(_12330_),
    .Y(_12333_));
 sky130_fd_sc_hd__nor2_2 _15232_ (.A(_11713_),
    .B(_12333_),
    .Y(_12334_));
 sky130_fd_sc_hd__a22o_2 _15233_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][12] ),
    .B1(_12332_),
    .B2(_12334_),
    .X(_01054_));
 sky130_fd_sc_hd__xor2_2 _15234_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[14][13] ),
    .X(_12335_));
 sky130_fd_sc_hd__a211o_2 _15235_ (.A1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[14][12] ),
    .B1(_12333_),
    .C1(_12335_),
    .X(_12336_));
 sky130_fd_sc_hd__nand2_2 _15236_ (.A(_12331_),
    .B(_12335_),
    .Y(_12337_));
 sky130_fd_sc_hd__and3_2 _15237_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[14][12] ),
    .C(_12335_),
    .X(_12338_));
 sky130_fd_sc_hd__a21oi_2 _15238_ (.A1(_12333_),
    .A2(_12335_),
    .B1(_12338_),
    .Y(_12339_));
 sky130_fd_sc_hd__a32o_2 _15239_ (.A1(_11712_),
    .A2(_12336_),
    .A3(_12339_),
    .B1(\systolic_inst.acc_wires[14][13] ),
    .B2(_11258_),
    .X(_01055_));
 sky130_fd_sc_hd__or2_2 _15240_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[14][14] ),
    .X(_12340_));
 sky130_fd_sc_hd__nand2_2 _15241_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[14][14] ),
    .Y(_12341_));
 sky130_fd_sc_hd__and2_2 _15242_ (.A(_12340_),
    .B(_12341_),
    .X(_12342_));
 sky130_fd_sc_hd__a21oi_2 _15243_ (.A1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[14][13] ),
    .B1(_12338_),
    .Y(_12343_));
 sky130_fd_sc_hd__o21ai_2 _15244_ (.A1(_12329_),
    .A2(_12337_),
    .B1(_12343_),
    .Y(_12344_));
 sky130_fd_sc_hd__nand2_2 _15245_ (.A(_12342_),
    .B(_12344_),
    .Y(_12345_));
 sky130_fd_sc_hd__or2_2 _15246_ (.A(_12342_),
    .B(_12344_),
    .X(_12346_));
 sky130_fd_sc_hd__a32o_2 _15247_ (.A1(_11712_),
    .A2(_12345_),
    .A3(_12346_),
    .B1(\systolic_inst.acc_wires[14][14] ),
    .B2(_11258_),
    .X(_01056_));
 sky130_fd_sc_hd__nor2_2 _15248_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][15] ),
    .Y(_12347_));
 sky130_fd_sc_hd__and2_2 _15249_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][15] ),
    .X(_12348_));
 sky130_fd_sc_hd__o211ai_2 _15250_ (.A1(_12347_),
    .A2(_12348_),
    .B1(_12341_),
    .C1(_12345_),
    .Y(_12349_));
 sky130_fd_sc_hd__a211o_2 _15251_ (.A1(_12341_),
    .A2(_12345_),
    .B1(_12347_),
    .C1(_12348_),
    .X(_12350_));
 sky130_fd_sc_hd__a32o_2 _15252_ (.A1(_11712_),
    .A2(_12349_),
    .A3(_12350_),
    .B1(\systolic_inst.acc_wires[14][15] ),
    .B2(_11258_),
    .X(_01057_));
 sky130_fd_sc_hd__or3b_2 _15253_ (.A(_12347_),
    .B(_12348_),
    .C_N(_12342_),
    .X(_12351_));
 sky130_fd_sc_hd__or2_2 _15254_ (.A(_12343_),
    .B(_12351_),
    .X(_12352_));
 sky130_fd_sc_hd__o31a_2 _15255_ (.A1(_12329_),
    .A2(_12337_),
    .A3(_12351_),
    .B1(_12352_),
    .X(_12353_));
 sky130_fd_sc_hd__o21ba_2 _15256_ (.A1(_12341_),
    .A2(_12347_),
    .B1_N(_12348_),
    .X(_12354_));
 sky130_fd_sc_hd__and2_2 _15257_ (.A(_12353_),
    .B(_12354_),
    .X(_12355_));
 sky130_fd_sc_hd__xnor2_2 _15258_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][16] ),
    .Y(_12356_));
 sky130_fd_sc_hd__nand2_2 _15259_ (.A(_12355_),
    .B(_12356_),
    .Y(_12357_));
 sky130_fd_sc_hd__nor2_2 _15260_ (.A(_12355_),
    .B(_12356_),
    .Y(_12358_));
 sky130_fd_sc_hd__nor2_2 _15261_ (.A(_11713_),
    .B(_12358_),
    .Y(_12359_));
 sky130_fd_sc_hd__a22o_2 _15262_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][16] ),
    .B1(_12357_),
    .B2(_12359_),
    .X(_01058_));
 sky130_fd_sc_hd__xor2_2 _15263_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][17] ),
    .X(_12360_));
 sky130_fd_sc_hd__inv_2 _15264_ (.A(_12360_),
    .Y(_12361_));
 sky130_fd_sc_hd__a21oi_2 _15265_ (.A1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[14][16] ),
    .B1(_12358_),
    .Y(_12362_));
 sky130_fd_sc_hd__xnor2_2 _15266_ (.A(_12360_),
    .B(_12362_),
    .Y(_12363_));
 sky130_fd_sc_hd__a22o_2 _15267_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][17] ),
    .B1(_11712_),
    .B2(_12363_),
    .X(_01059_));
 sky130_fd_sc_hd__or2_2 _15268_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][18] ),
    .X(_12364_));
 sky130_fd_sc_hd__nand2_2 _15269_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][18] ),
    .Y(_12365_));
 sky130_fd_sc_hd__nand2_2 _15270_ (.A(_12364_),
    .B(_12365_),
    .Y(_12366_));
 sky130_fd_sc_hd__o21a_2 _15271_ (.A1(\systolic_inst.acc_wires[14][16] ),
    .A2(\systolic_inst.acc_wires[14][17] ),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .X(_12367_));
 sky130_fd_sc_hd__a21oi_2 _15272_ (.A1(_12358_),
    .A2(_12360_),
    .B1(_12367_),
    .Y(_12368_));
 sky130_fd_sc_hd__xor2_2 _15273_ (.A(_12366_),
    .B(_12368_),
    .X(_12369_));
 sky130_fd_sc_hd__a22o_2 _15274_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][18] ),
    .B1(_11712_),
    .B2(_12369_),
    .X(_01060_));
 sky130_fd_sc_hd__xnor2_2 _15275_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][19] ),
    .Y(_12370_));
 sky130_fd_sc_hd__o21ai_2 _15276_ (.A1(_12366_),
    .A2(_12368_),
    .B1(_12365_),
    .Y(_12371_));
 sky130_fd_sc_hd__xnor2_2 _15277_ (.A(_12370_),
    .B(_12371_),
    .Y(_12372_));
 sky130_fd_sc_hd__a22o_2 _15278_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][19] ),
    .B1(_11712_),
    .B2(_12372_),
    .X(_01061_));
 sky130_fd_sc_hd__or2_2 _15279_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][20] ),
    .X(_12373_));
 sky130_fd_sc_hd__nand2_2 _15280_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][20] ),
    .Y(_12374_));
 sky130_fd_sc_hd__and2_2 _15281_ (.A(_12373_),
    .B(_12374_),
    .X(_12375_));
 sky130_fd_sc_hd__or4_2 _15282_ (.A(_12356_),
    .B(_12361_),
    .C(_12366_),
    .D(_12370_),
    .X(_12376_));
 sky130_fd_sc_hd__nor2_2 _15283_ (.A(_12355_),
    .B(_12376_),
    .Y(_12377_));
 sky130_fd_sc_hd__o41a_2 _15284_ (.A1(\systolic_inst.acc_wires[14][16] ),
    .A2(\systolic_inst.acc_wires[14][17] ),
    .A3(\systolic_inst.acc_wires[14][18] ),
    .A4(\systolic_inst.acc_wires[14][19] ),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .X(_12378_));
 sky130_fd_sc_hd__o21ai_2 _15285_ (.A1(_12377_),
    .A2(_12378_),
    .B1(_12375_),
    .Y(_12379_));
 sky130_fd_sc_hd__or3_2 _15286_ (.A(_12375_),
    .B(_12377_),
    .C(_12378_),
    .X(_12380_));
 sky130_fd_sc_hd__a32o_2 _15287_ (.A1(_11712_),
    .A2(_12379_),
    .A3(_12380_),
    .B1(\systolic_inst.acc_wires[14][20] ),
    .B2(_11258_),
    .X(_01062_));
 sky130_fd_sc_hd__xnor2_2 _15288_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][21] ),
    .Y(_12381_));
 sky130_fd_sc_hd__inv_2 _15289_ (.A(_12381_),
    .Y(_12382_));
 sky130_fd_sc_hd__a21oi_2 _15290_ (.A1(_12374_),
    .A2(_12379_),
    .B1(_12381_),
    .Y(_12383_));
 sky130_fd_sc_hd__a31o_2 _15291_ (.A1(_12374_),
    .A2(_12379_),
    .A3(_12381_),
    .B1(_11713_),
    .X(_12384_));
 sky130_fd_sc_hd__a2bb2o_2 _15292_ (.A1_N(_12384_),
    .A2_N(_12383_),
    .B1(\systolic_inst.acc_wires[14][21] ),
    .B2(_11258_),
    .X(_01063_));
 sky130_fd_sc_hd__or2_2 _15293_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][22] ),
    .X(_12385_));
 sky130_fd_sc_hd__nand2_2 _15294_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][22] ),
    .Y(_12386_));
 sky130_fd_sc_hd__and2_2 _15295_ (.A(_12385_),
    .B(_12386_),
    .X(_12387_));
 sky130_fd_sc_hd__o21a_2 _15296_ (.A1(\systolic_inst.acc_wires[14][20] ),
    .A2(\systolic_inst.acc_wires[14][21] ),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .X(_12388_));
 sky130_fd_sc_hd__nor2_2 _15297_ (.A(_12379_),
    .B(_12381_),
    .Y(_12389_));
 sky130_fd_sc_hd__o21ai_2 _15298_ (.A1(_12388_),
    .A2(_12389_),
    .B1(_12387_),
    .Y(_12390_));
 sky130_fd_sc_hd__or3_2 _15299_ (.A(_12387_),
    .B(_12388_),
    .C(_12389_),
    .X(_12391_));
 sky130_fd_sc_hd__a32o_2 _15300_ (.A1(_11712_),
    .A2(_12390_),
    .A3(_12391_),
    .B1(\systolic_inst.acc_wires[14][22] ),
    .B2(_11258_),
    .X(_01064_));
 sky130_fd_sc_hd__xor2_2 _15301_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][23] ),
    .X(_12392_));
 sky130_fd_sc_hd__inv_2 _15302_ (.A(_12392_),
    .Y(_12393_));
 sky130_fd_sc_hd__nand3_2 _15303_ (.A(_12386_),
    .B(_12390_),
    .C(_12393_),
    .Y(_12394_));
 sky130_fd_sc_hd__a21o_2 _15304_ (.A1(_12386_),
    .A2(_12390_),
    .B1(_12393_),
    .X(_12395_));
 sky130_fd_sc_hd__a32o_2 _15305_ (.A1(_11712_),
    .A2(_12394_),
    .A3(_12395_),
    .B1(\systolic_inst.acc_wires[14][23] ),
    .B2(_11258_),
    .X(_01065_));
 sky130_fd_sc_hd__nand4_2 _15306_ (.A(_12375_),
    .B(_12382_),
    .C(_12387_),
    .D(_12392_),
    .Y(_12396_));
 sky130_fd_sc_hd__a211o_2 _15307_ (.A1(_12353_),
    .A2(_12354_),
    .B1(_12376_),
    .C1(_12396_),
    .X(_12397_));
 sky130_fd_sc_hd__o41a_2 _15308_ (.A1(\systolic_inst.acc_wires[14][20] ),
    .A2(\systolic_inst.acc_wires[14][21] ),
    .A3(\systolic_inst.acc_wires[14][22] ),
    .A4(\systolic_inst.acc_wires[14][23] ),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .X(_12398_));
 sky130_fd_sc_hd__nor2_2 _15309_ (.A(_12378_),
    .B(_12398_),
    .Y(_12399_));
 sky130_fd_sc_hd__nor2_2 _15310_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][24] ),
    .Y(_12400_));
 sky130_fd_sc_hd__and2_2 _15311_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][24] ),
    .X(_12401_));
 sky130_fd_sc_hd__or2_2 _15312_ (.A(_12400_),
    .B(_12401_),
    .X(_12402_));
 sky130_fd_sc_hd__a21oi_2 _15313_ (.A1(_12397_),
    .A2(_12399_),
    .B1(_12402_),
    .Y(_12403_));
 sky130_fd_sc_hd__a31o_2 _15314_ (.A1(_12397_),
    .A2(_12399_),
    .A3(_12402_),
    .B1(_11713_),
    .X(_12404_));
 sky130_fd_sc_hd__a2bb2o_2 _15315_ (.A1_N(_12404_),
    .A2_N(_12403_),
    .B1(\systolic_inst.acc_wires[14][24] ),
    .B2(_11258_),
    .X(_01066_));
 sky130_fd_sc_hd__xor2_2 _15316_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][25] ),
    .X(_12405_));
 sky130_fd_sc_hd__or3_2 _15317_ (.A(_12401_),
    .B(_12403_),
    .C(_12405_),
    .X(_12406_));
 sky130_fd_sc_hd__o21ai_2 _15318_ (.A1(_12401_),
    .A2(_12403_),
    .B1(_12405_),
    .Y(_12407_));
 sky130_fd_sc_hd__a32o_2 _15319_ (.A1(_11712_),
    .A2(_12406_),
    .A3(_12407_),
    .B1(\systolic_inst.acc_wires[14][25] ),
    .B2(_11258_),
    .X(_01067_));
 sky130_fd_sc_hd__or2_2 _15320_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][26] ),
    .X(_12408_));
 sky130_fd_sc_hd__nand2_2 _15321_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][26] ),
    .Y(_12409_));
 sky130_fd_sc_hd__nand2_2 _15322_ (.A(_12408_),
    .B(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__o21a_2 _15323_ (.A1(\systolic_inst.acc_wires[14][24] ),
    .A2(\systolic_inst.acc_wires[14][25] ),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .X(_12411_));
 sky130_fd_sc_hd__a21o_2 _15324_ (.A1(_12403_),
    .A2(_12405_),
    .B1(_12411_),
    .X(_12412_));
 sky130_fd_sc_hd__xnor2_2 _15325_ (.A(_12410_),
    .B(_12412_),
    .Y(_12413_));
 sky130_fd_sc_hd__a22o_2 _15326_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][26] ),
    .B1(_11712_),
    .B2(_12413_),
    .X(_01068_));
 sky130_fd_sc_hd__xnor2_2 _15327_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][27] ),
    .Y(_12414_));
 sky130_fd_sc_hd__a21bo_2 _15328_ (.A1(_12408_),
    .A2(_12412_),
    .B1_N(_12409_),
    .X(_12415_));
 sky130_fd_sc_hd__xnor2_2 _15329_ (.A(_12414_),
    .B(_12415_),
    .Y(_12416_));
 sky130_fd_sc_hd__a22o_2 _15330_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][27] ),
    .B1(_11712_),
    .B2(_12416_),
    .X(_01069_));
 sky130_fd_sc_hd__nor2_2 _15331_ (.A(_12410_),
    .B(_12414_),
    .Y(_12417_));
 sky130_fd_sc_hd__o21a_2 _15332_ (.A1(\systolic_inst.acc_wires[14][26] ),
    .A2(\systolic_inst.acc_wires[14][27] ),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .X(_12418_));
 sky130_fd_sc_hd__a311oi_2 _15333_ (.A1(_12403_),
    .A2(_12405_),
    .A3(_12417_),
    .B1(_12418_),
    .C1(_12411_),
    .Y(_12419_));
 sky130_fd_sc_hd__or2_2 _15334_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][28] ),
    .X(_12420_));
 sky130_fd_sc_hd__nand2_2 _15335_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][28] ),
    .Y(_12421_));
 sky130_fd_sc_hd__nand2_2 _15336_ (.A(_12420_),
    .B(_12421_),
    .Y(_12422_));
 sky130_fd_sc_hd__xor2_2 _15337_ (.A(_12419_),
    .B(_12422_),
    .X(_12423_));
 sky130_fd_sc_hd__a22o_2 _15338_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][28] ),
    .B1(_11712_),
    .B2(_12423_),
    .X(_01070_));
 sky130_fd_sc_hd__xor2_2 _15339_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][29] ),
    .X(_12424_));
 sky130_fd_sc_hd__inv_2 _15340_ (.A(_12424_),
    .Y(_12425_));
 sky130_fd_sc_hd__o21a_2 _15341_ (.A1(_12419_),
    .A2(_12422_),
    .B1(_12421_),
    .X(_12426_));
 sky130_fd_sc_hd__xnor2_2 _15342_ (.A(_12424_),
    .B(_12426_),
    .Y(_12427_));
 sky130_fd_sc_hd__a22o_2 _15343_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[14][29] ),
    .B1(_11712_),
    .B2(_12427_),
    .X(_01071_));
 sky130_fd_sc_hd__o21ai_2 _15344_ (.A1(\systolic_inst.acc_wires[14][28] ),
    .A2(\systolic_inst.acc_wires[14][29] ),
    .B1(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .Y(_12428_));
 sky130_fd_sc_hd__o31a_2 _15345_ (.A1(_12419_),
    .A2(_12422_),
    .A3(_12425_),
    .B1(_12428_),
    .X(_12429_));
 sky130_fd_sc_hd__nand2_2 _15346_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][30] ),
    .Y(_12430_));
 sky130_fd_sc_hd__or2_2 _15347_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][30] ),
    .X(_12431_));
 sky130_fd_sc_hd__nand2_2 _15348_ (.A(_12430_),
    .B(_12431_),
    .Y(_12432_));
 sky130_fd_sc_hd__nand2_2 _15349_ (.A(_12429_),
    .B(_12432_),
    .Y(_12433_));
 sky130_fd_sc_hd__or2_2 _15350_ (.A(_12429_),
    .B(_12432_),
    .X(_12434_));
 sky130_fd_sc_hd__a32o_2 _15351_ (.A1(_11712_),
    .A2(_12433_),
    .A3(_12434_),
    .B1(\systolic_inst.acc_wires[14][30] ),
    .B2(_11258_),
    .X(_01072_));
 sky130_fd_sc_hd__xnor2_2 _15352_ (.A(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[14][31] ),
    .Y(_12435_));
 sky130_fd_sc_hd__a21oi_2 _15353_ (.A1(_12430_),
    .A2(_12434_),
    .B1(_12435_),
    .Y(_12436_));
 sky130_fd_sc_hd__a31o_2 _15354_ (.A1(_12430_),
    .A2(_12434_),
    .A3(_12435_),
    .B1(_11713_),
    .X(_12437_));
 sky130_fd_sc_hd__a2bb2o_2 _15355_ (.A1_N(_12437_),
    .A2_N(_12436_),
    .B1(\systolic_inst.acc_wires[14][31] ),
    .B2(_11258_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _15356_ (.A0(\systolic_inst.A_outs[13][0] ),
    .A1(\systolic_inst.A_outs[12][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _15357_ (.A0(\systolic_inst.A_outs[13][1] ),
    .A1(\systolic_inst.A_outs[12][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _15358_ (.A0(\systolic_inst.A_outs[13][2] ),
    .A1(\systolic_inst.A_outs[12][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _15359_ (.A0(\systolic_inst.A_outs[13][3] ),
    .A1(\systolic_inst.A_outs[12][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _15360_ (.A0(\systolic_inst.A_outs[13][4] ),
    .A1(\systolic_inst.A_outs[12][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _15361_ (.A0(\systolic_inst.A_outs[13][5] ),
    .A1(\systolic_inst.A_outs[12][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _15362_ (.A0(\systolic_inst.A_outs[13][6] ),
    .A1(\systolic_inst.A_outs[12][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _15363_ (.A0(\systolic_inst.A_outs[13][7] ),
    .A1(\systolic_inst.A_outs[12][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _15364_ (.A0(\systolic_inst.B_outs[12][0] ),
    .A1(\systolic_inst.B_outs[8][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _15365_ (.A0(\systolic_inst.B_outs[12][1] ),
    .A1(\systolic_inst.B_outs[8][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _15366_ (.A0(\systolic_inst.B_outs[12][2] ),
    .A1(\systolic_inst.B_outs[8][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _15367_ (.A0(\systolic_inst.B_outs[12][3] ),
    .A1(\systolic_inst.B_outs[8][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _15368_ (.A0(\systolic_inst.B_outs[12][4] ),
    .A1(\systolic_inst.B_outs[8][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _15369_ (.A0(\systolic_inst.B_outs[12][5] ),
    .A1(\systolic_inst.B_outs[8][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _15370_ (.A0(\systolic_inst.B_outs[12][6] ),
    .A1(\systolic_inst.B_outs[8][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _15371_ (.A0(\systolic_inst.B_outs[12][7] ),
    .A1(\systolic_inst.B_outs[8][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01089_));
 sky130_fd_sc_hd__and3_2 _15372_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[13][0] ),
    .C(\systolic_inst.A_outs[13][0] ),
    .X(_12438_));
 sky130_fd_sc_hd__a21o_2 _15373_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[0] ),
    .B1(_12438_),
    .X(_01090_));
 sky130_fd_sc_hd__and4_2 _15374_ (.A(\systolic_inst.B_outs[13][0] ),
    .B(\systolic_inst.A_outs[13][0] ),
    .C(\systolic_inst.B_outs[13][1] ),
    .D(\systolic_inst.A_outs[13][1] ),
    .X(_12439_));
 sky130_fd_sc_hd__a22o_2 _15375_ (.A1(\systolic_inst.A_outs[13][0] ),
    .A2(\systolic_inst.B_outs[13][1] ),
    .B1(\systolic_inst.A_outs[13][1] ),
    .B2(\systolic_inst.B_outs[13][0] ),
    .X(_12440_));
 sky130_fd_sc_hd__nand2_2 _15376_ (.A(\systolic_inst.ce_local ),
    .B(_12440_),
    .Y(_12441_));
 sky130_fd_sc_hd__a2bb2o_2 _15377_ (.A1_N(_12441_),
    .A2_N(_12439_),
    .B1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01091_));
 sky130_fd_sc_hd__and2_2 _15378_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[2] ),
    .X(_12442_));
 sky130_fd_sc_hd__a22oi_2 _15379_ (.A1(\systolic_inst.B_outs[13][1] ),
    .A2(\systolic_inst.A_outs[13][1] ),
    .B1(\systolic_inst.A_outs[13][2] ),
    .B2(\systolic_inst.B_outs[13][0] ),
    .Y(_12443_));
 sky130_fd_sc_hd__and4_2 _15380_ (.A(\systolic_inst.B_outs[13][0] ),
    .B(\systolic_inst.B_outs[13][1] ),
    .C(\systolic_inst.A_outs[13][1] ),
    .D(\systolic_inst.A_outs[13][2] ),
    .X(_12444_));
 sky130_fd_sc_hd__or2_2 _15381_ (.A(_12443_),
    .B(_12444_),
    .X(_12445_));
 sky130_fd_sc_hd__or3b_2 _15382_ (.A(_12443_),
    .B(_12444_),
    .C_N(_12439_),
    .X(_12446_));
 sky130_fd_sc_hd__xnor2_2 _15383_ (.A(_12439_),
    .B(_12445_),
    .Y(_12447_));
 sky130_fd_sc_hd__nand3_2 _15384_ (.A(\systolic_inst.A_outs[13][0] ),
    .B(\systolic_inst.B_outs[13][2] ),
    .C(_12447_),
    .Y(_12448_));
 sky130_fd_sc_hd__a21o_2 _15385_ (.A1(\systolic_inst.A_outs[13][0] ),
    .A2(\systolic_inst.B_outs[13][2] ),
    .B1(_12447_),
    .X(_12449_));
 sky130_fd_sc_hd__a31o_2 _15386_ (.A1(\systolic_inst.ce_local ),
    .A2(_12448_),
    .A3(_12449_),
    .B1(_12442_),
    .X(_01092_));
 sky130_fd_sc_hd__a22oi_2 _15387_ (.A1(\systolic_inst.A_outs[13][1] ),
    .A2(\systolic_inst.B_outs[13][2] ),
    .B1(\systolic_inst.B_outs[13][3] ),
    .B2(\systolic_inst.A_outs[13][0] ),
    .Y(_12450_));
 sky130_fd_sc_hd__and4_2 _15388_ (.A(\systolic_inst.A_outs[13][0] ),
    .B(\systolic_inst.A_outs[13][1] ),
    .C(\systolic_inst.B_outs[13][2] ),
    .D(\systolic_inst.B_outs[13][3] ),
    .X(_12451_));
 sky130_fd_sc_hd__nor2_2 _15389_ (.A(_12450_),
    .B(_12451_),
    .Y(_12452_));
 sky130_fd_sc_hd__nand4_2 _15390_ (.A(\systolic_inst.B_outs[13][0] ),
    .B(\systolic_inst.B_outs[13][1] ),
    .C(\systolic_inst.A_outs[13][2] ),
    .D(\systolic_inst.A_outs[13][3] ),
    .Y(_12453_));
 sky130_fd_sc_hd__a22o_2 _15391_ (.A1(\systolic_inst.B_outs[13][1] ),
    .A2(\systolic_inst.A_outs[13][2] ),
    .B1(\systolic_inst.A_outs[13][3] ),
    .B2(\systolic_inst.B_outs[13][0] ),
    .X(_12454_));
 sky130_fd_sc_hd__nand3_2 _15392_ (.A(_12444_),
    .B(_12453_),
    .C(_12454_),
    .Y(_12455_));
 sky130_fd_sc_hd__a21o_2 _15393_ (.A1(_12453_),
    .A2(_12454_),
    .B1(_12444_),
    .X(_12456_));
 sky130_fd_sc_hd__and2_2 _15394_ (.A(_12455_),
    .B(_12456_),
    .X(_12457_));
 sky130_fd_sc_hd__nand2_2 _15395_ (.A(_12452_),
    .B(_12457_),
    .Y(_12458_));
 sky130_fd_sc_hd__xnor2_2 _15396_ (.A(_12452_),
    .B(_12457_),
    .Y(_12459_));
 sky130_fd_sc_hd__and3_2 _15397_ (.A(_12446_),
    .B(_12448_),
    .C(_12459_),
    .X(_12460_));
 sky130_fd_sc_hd__a21oi_2 _15398_ (.A1(_12446_),
    .A2(_12448_),
    .B1(_12459_),
    .Y(_12461_));
 sky130_fd_sc_hd__nand2_2 _15399_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[3] ),
    .Y(_12462_));
 sky130_fd_sc_hd__o31ai_2 _15400_ (.A1(_11258_),
    .A2(_12460_),
    .A3(_12461_),
    .B1(_12462_),
    .Y(_01093_));
 sky130_fd_sc_hd__and2_2 _15401_ (.A(\systolic_inst.B_outs[13][2] ),
    .B(\systolic_inst.A_outs[13][2] ),
    .X(_12463_));
 sky130_fd_sc_hd__nand4_2 _15402_ (.A(\systolic_inst.A_outs[13][0] ),
    .B(\systolic_inst.A_outs[13][1] ),
    .C(\systolic_inst.B_outs[13][3] ),
    .D(\systolic_inst.B_outs[13][4] ),
    .Y(_12464_));
 sky130_fd_sc_hd__a22o_2 _15403_ (.A1(\systolic_inst.A_outs[13][1] ),
    .A2(\systolic_inst.B_outs[13][3] ),
    .B1(\systolic_inst.B_outs[13][4] ),
    .B2(\systolic_inst.A_outs[13][0] ),
    .X(_12465_));
 sky130_fd_sc_hd__nand2_2 _15404_ (.A(_12464_),
    .B(_12465_),
    .Y(_12466_));
 sky130_fd_sc_hd__xnor2_2 _15405_ (.A(_12463_),
    .B(_12466_),
    .Y(_12467_));
 sky130_fd_sc_hd__a22o_2 _15406_ (.A1(\systolic_inst.B_outs[13][1] ),
    .A2(\systolic_inst.A_outs[13][3] ),
    .B1(\systolic_inst.A_outs[13][4] ),
    .B2(\systolic_inst.B_outs[13][0] ),
    .X(_12468_));
 sky130_fd_sc_hd__and3_2 _15407_ (.A(\systolic_inst.B_outs[13][0] ),
    .B(\systolic_inst.B_outs[13][1] ),
    .C(\systolic_inst.A_outs[13][3] ),
    .X(_12469_));
 sky130_fd_sc_hd__nand2_2 _15408_ (.A(\systolic_inst.A_outs[13][4] ),
    .B(_12469_),
    .Y(_12470_));
 sky130_fd_sc_hd__and3_2 _15409_ (.A(_12451_),
    .B(_12468_),
    .C(_12470_),
    .X(_12471_));
 sky130_fd_sc_hd__a21oi_2 _15410_ (.A1(_12468_),
    .A2(_12470_),
    .B1(_12451_),
    .Y(_12472_));
 sky130_fd_sc_hd__o21ai_2 _15411_ (.A1(_12471_),
    .A2(_12472_),
    .B1(_12453_),
    .Y(_12473_));
 sky130_fd_sc_hd__or3_2 _15412_ (.A(_12453_),
    .B(_12471_),
    .C(_12472_),
    .X(_12474_));
 sky130_fd_sc_hd__and3_2 _15413_ (.A(_12467_),
    .B(_12473_),
    .C(_12474_),
    .X(_12475_));
 sky130_fd_sc_hd__a21oi_2 _15414_ (.A1(_12473_),
    .A2(_12474_),
    .B1(_12467_),
    .Y(_12476_));
 sky130_fd_sc_hd__a211o_2 _15415_ (.A1(_12455_),
    .A2(_12458_),
    .B1(_12475_),
    .C1(_12476_),
    .X(_12477_));
 sky130_fd_sc_hd__o211ai_2 _15416_ (.A1(_12475_),
    .A2(_12476_),
    .B1(_12455_),
    .C1(_12458_),
    .Y(_12478_));
 sky130_fd_sc_hd__a21oi_2 _15417_ (.A1(_12477_),
    .A2(_12478_),
    .B1(_12461_),
    .Y(_12479_));
 sky130_fd_sc_hd__and3_2 _15418_ (.A(_12461_),
    .B(_12477_),
    .C(_12478_),
    .X(_12480_));
 sky130_fd_sc_hd__or3_2 _15419_ (.A(_11258_),
    .B(_12479_),
    .C(_12480_),
    .X(_12481_));
 sky130_fd_sc_hd__a21bo_2 _15420_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[4] ),
    .B1_N(_12481_),
    .X(_01094_));
 sky130_fd_sc_hd__and2b_2 _15421_ (.A_N(_12471_),
    .B(_12474_),
    .X(_12482_));
 sky130_fd_sc_hd__a21bo_2 _15422_ (.A1(_12463_),
    .A2(_12465_),
    .B1_N(_12464_),
    .X(_12483_));
 sky130_fd_sc_hd__a22oi_2 _15423_ (.A1(\systolic_inst.B_outs[13][1] ),
    .A2(\systolic_inst.A_outs[13][4] ),
    .B1(\systolic_inst.A_outs[13][5] ),
    .B2(\systolic_inst.B_outs[13][0] ),
    .Y(_12484_));
 sky130_fd_sc_hd__and4_2 _15424_ (.A(\systolic_inst.B_outs[13][0] ),
    .B(\systolic_inst.B_outs[13][1] ),
    .C(\systolic_inst.A_outs[13][4] ),
    .D(\systolic_inst.A_outs[13][5] ),
    .X(_12485_));
 sky130_fd_sc_hd__nor2_2 _15425_ (.A(_12484_),
    .B(_12485_),
    .Y(_12486_));
 sky130_fd_sc_hd__xor2_2 _15426_ (.A(_12483_),
    .B(_12486_),
    .X(_12487_));
 sky130_fd_sc_hd__xor2_2 _15427_ (.A(_12470_),
    .B(_12487_),
    .X(_12488_));
 sky130_fd_sc_hd__and4_2 _15428_ (.A(\systolic_inst.A_outs[13][1] ),
    .B(\systolic_inst.A_outs[13][2] ),
    .C(\systolic_inst.B_outs[13][3] ),
    .D(\systolic_inst.B_outs[13][4] ),
    .X(_12489_));
 sky130_fd_sc_hd__a22oi_2 _15429_ (.A1(\systolic_inst.A_outs[13][2] ),
    .A2(\systolic_inst.B_outs[13][3] ),
    .B1(\systolic_inst.B_outs[13][4] ),
    .B2(\systolic_inst.A_outs[13][1] ),
    .Y(_12490_));
 sky130_fd_sc_hd__a22o_2 _15430_ (.A1(\systolic_inst.A_outs[13][2] ),
    .A2(\systolic_inst.B_outs[13][3] ),
    .B1(\systolic_inst.B_outs[13][4] ),
    .B2(\systolic_inst.A_outs[13][1] ),
    .X(_12491_));
 sky130_fd_sc_hd__and4b_2 _15431_ (.A_N(_12489_),
    .B(_12491_),
    .C(\systolic_inst.B_outs[13][2] ),
    .D(\systolic_inst.A_outs[13][3] ),
    .X(_12492_));
 sky130_fd_sc_hd__o2bb2a_2 _15432_ (.A1_N(\systolic_inst.B_outs[13][2] ),
    .A2_N(\systolic_inst.A_outs[13][3] ),
    .B1(_12489_),
    .B2(_12490_),
    .X(_12493_));
 sky130_fd_sc_hd__and4bb_2 _15433_ (.A_N(_12492_),
    .B_N(_12493_),
    .C(\systolic_inst.A_outs[13][0] ),
    .D(\systolic_inst.B_outs[13][5] ),
    .X(_12494_));
 sky130_fd_sc_hd__o2bb2a_2 _15434_ (.A1_N(\systolic_inst.A_outs[13][0] ),
    .A2_N(\systolic_inst.B_outs[13][5] ),
    .B1(_12492_),
    .B2(_12493_),
    .X(_12495_));
 sky130_fd_sc_hd__or2_2 _15435_ (.A(_12494_),
    .B(_12495_),
    .X(_12496_));
 sky130_fd_sc_hd__nor2_2 _15436_ (.A(_12488_),
    .B(_12496_),
    .Y(_12497_));
 sky130_fd_sc_hd__xor2_2 _15437_ (.A(_12488_),
    .B(_12496_),
    .X(_12498_));
 sky130_fd_sc_hd__nand2_2 _15438_ (.A(_12475_),
    .B(_12498_),
    .Y(_12499_));
 sky130_fd_sc_hd__xor2_2 _15439_ (.A(_12475_),
    .B(_12498_),
    .X(_12500_));
 sky130_fd_sc_hd__nand2b_2 _15440_ (.A_N(_12482_),
    .B(_12500_),
    .Y(_12501_));
 sky130_fd_sc_hd__xnor2_2 _15441_ (.A(_12482_),
    .B(_12500_),
    .Y(_12502_));
 sky130_fd_sc_hd__a21bo_2 _15442_ (.A1(_12461_),
    .A2(_12478_),
    .B1_N(_12477_),
    .X(_12503_));
 sky130_fd_sc_hd__nand2_2 _15443_ (.A(_12502_),
    .B(_12503_),
    .Y(_12504_));
 sky130_fd_sc_hd__o21a_2 _15444_ (.A1(_12502_),
    .A2(_12503_),
    .B1(\systolic_inst.ce_local ),
    .X(_12505_));
 sky130_fd_sc_hd__a22o_2 _15445_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[5] ),
    .B1(_12504_),
    .B2(_12505_),
    .X(_01095_));
 sky130_fd_sc_hd__a32o_2 _15446_ (.A1(\systolic_inst.A_outs[13][4] ),
    .A2(_12469_),
    .A3(_12487_),
    .B1(_12486_),
    .B2(_12483_),
    .X(_12506_));
 sky130_fd_sc_hd__inv_2 _15447_ (.A(_12506_),
    .Y(_12507_));
 sky130_fd_sc_hd__a31o_2 _15448_ (.A1(\systolic_inst.B_outs[13][2] ),
    .A2(\systolic_inst.A_outs[13][3] ),
    .A3(_12491_),
    .B1(_12489_),
    .X(_12508_));
 sky130_fd_sc_hd__a22oi_2 _15449_ (.A1(\systolic_inst.B_outs[13][1] ),
    .A2(\systolic_inst.A_outs[13][5] ),
    .B1(\systolic_inst.A_outs[13][6] ),
    .B2(\systolic_inst.B_outs[13][0] ),
    .Y(_12509_));
 sky130_fd_sc_hd__and4_2 _15450_ (.A(\systolic_inst.B_outs[13][0] ),
    .B(\systolic_inst.B_outs[13][1] ),
    .C(\systolic_inst.A_outs[13][5] ),
    .D(\systolic_inst.A_outs[13][6] ),
    .X(_12510_));
 sky130_fd_sc_hd__or2_2 _15451_ (.A(_12509_),
    .B(_12510_),
    .X(_12511_));
 sky130_fd_sc_hd__and2b_2 _15452_ (.A_N(_12511_),
    .B(_12508_),
    .X(_12512_));
 sky130_fd_sc_hd__xnor2_2 _15453_ (.A(_12508_),
    .B(_12511_),
    .Y(_12513_));
 sky130_fd_sc_hd__xor2_2 _15454_ (.A(_12485_),
    .B(_12513_),
    .X(_12514_));
 sky130_fd_sc_hd__nand4_2 _15455_ (.A(\systolic_inst.A_outs[13][2] ),
    .B(\systolic_inst.B_outs[13][3] ),
    .C(\systolic_inst.A_outs[13][3] ),
    .D(\systolic_inst.B_outs[13][4] ),
    .Y(_12515_));
 sky130_fd_sc_hd__a22o_2 _15456_ (.A1(\systolic_inst.B_outs[13][3] ),
    .A2(\systolic_inst.A_outs[13][3] ),
    .B1(\systolic_inst.B_outs[13][4] ),
    .B2(\systolic_inst.A_outs[13][2] ),
    .X(_12516_));
 sky130_fd_sc_hd__nand4_2 _15457_ (.A(\systolic_inst.B_outs[13][2] ),
    .B(\systolic_inst.A_outs[13][4] ),
    .C(_12515_),
    .D(_12516_),
    .Y(_12517_));
 sky130_fd_sc_hd__a22o_2 _15458_ (.A1(\systolic_inst.B_outs[13][2] ),
    .A2(\systolic_inst.A_outs[13][4] ),
    .B1(_12515_),
    .B2(_12516_),
    .X(_12518_));
 sky130_fd_sc_hd__a22oi_2 _15459_ (.A1(\systolic_inst.A_outs[13][1] ),
    .A2(\systolic_inst.B_outs[13][5] ),
    .B1(\systolic_inst.B_outs[13][6] ),
    .B2(\systolic_inst.A_outs[13][0] ),
    .Y(_12519_));
 sky130_fd_sc_hd__nand2_2 _15460_ (.A(\systolic_inst.A_outs[13][1] ),
    .B(\systolic_inst.B_outs[13][6] ),
    .Y(_12520_));
 sky130_fd_sc_hd__and4_2 _15461_ (.A(\systolic_inst.A_outs[13][0] ),
    .B(\systolic_inst.A_outs[13][1] ),
    .C(\systolic_inst.B_outs[13][5] ),
    .D(\systolic_inst.B_outs[13][6] ),
    .X(_12521_));
 sky130_fd_sc_hd__nor2_2 _15462_ (.A(_12519_),
    .B(_12521_),
    .Y(_12522_));
 sky130_fd_sc_hd__nand3_2 _15463_ (.A(_12517_),
    .B(_12518_),
    .C(_12522_),
    .Y(_12523_));
 sky130_fd_sc_hd__a21o_2 _15464_ (.A1(_12517_),
    .A2(_12518_),
    .B1(_12522_),
    .X(_12524_));
 sky130_fd_sc_hd__and3_2 _15465_ (.A(_12494_),
    .B(_12523_),
    .C(_12524_),
    .X(_12525_));
 sky130_fd_sc_hd__a21oi_2 _15466_ (.A1(_12523_),
    .A2(_12524_),
    .B1(_12494_),
    .Y(_12526_));
 sky130_fd_sc_hd__or3b_2 _15467_ (.A(_12525_),
    .B(_12526_),
    .C_N(_12514_),
    .X(_12527_));
 sky130_fd_sc_hd__o21bai_2 _15468_ (.A1(_12525_),
    .A2(_12526_),
    .B1_N(_12514_),
    .Y(_12528_));
 sky130_fd_sc_hd__and3_2 _15469_ (.A(_12497_),
    .B(_12527_),
    .C(_12528_),
    .X(_12529_));
 sky130_fd_sc_hd__a21oi_2 _15470_ (.A1(_12527_),
    .A2(_12528_),
    .B1(_12497_),
    .Y(_12530_));
 sky130_fd_sc_hd__nor3_2 _15471_ (.A(_12507_),
    .B(_12529_),
    .C(_12530_),
    .Y(_12531_));
 sky130_fd_sc_hd__o21a_2 _15472_ (.A1(_12529_),
    .A2(_12530_),
    .B1(_12507_),
    .X(_12532_));
 sky130_fd_sc_hd__a211oi_2 _15473_ (.A1(_12499_),
    .A2(_12501_),
    .B1(_12531_),
    .C1(_12532_),
    .Y(_12533_));
 sky130_fd_sc_hd__o211a_2 _15474_ (.A1(_12531_),
    .A2(_12532_),
    .B1(_12499_),
    .C1(_12501_),
    .X(_12534_));
 sky130_fd_sc_hd__nor2_2 _15475_ (.A(_12533_),
    .B(_12534_),
    .Y(_12535_));
 sky130_fd_sc_hd__xnor2_2 _15476_ (.A(_12504_),
    .B(_12535_),
    .Y(_12536_));
 sky130_fd_sc_hd__mux2_1 _15477_ (.A0(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[6] ),
    .A1(_12536_),
    .S(\systolic_inst.ce_local ),
    .X(_01096_));
 sky130_fd_sc_hd__nor2_2 _15478_ (.A(_12529_),
    .B(_12531_),
    .Y(_12537_));
 sky130_fd_sc_hd__a21oi_2 _15479_ (.A1(_12485_),
    .A2(_12513_),
    .B1(_12512_),
    .Y(_12538_));
 sky130_fd_sc_hd__nand2_2 _15480_ (.A(_12515_),
    .B(_12517_),
    .Y(_12539_));
 sky130_fd_sc_hd__a22o_2 _15481_ (.A1(\systolic_inst.B_outs[13][1] ),
    .A2(\systolic_inst.A_outs[13][6] ),
    .B1(\systolic_inst.A_outs[13][7] ),
    .B2(\systolic_inst.B_outs[13][0] ),
    .X(_12540_));
 sky130_fd_sc_hd__nand4_2 _15482_ (.A(\systolic_inst.B_outs[13][0] ),
    .B(\systolic_inst.B_outs[13][1] ),
    .C(\systolic_inst.A_outs[13][6] ),
    .D(\systolic_inst.A_outs[13][7] ),
    .Y(_12541_));
 sky130_fd_sc_hd__nand2_2 _15483_ (.A(_12540_),
    .B(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__xnor2_2 _15484_ (.A(_11272_),
    .B(_12542_),
    .Y(_12543_));
 sky130_fd_sc_hd__nand2b_2 _15485_ (.A_N(_12543_),
    .B(_12539_),
    .Y(_12544_));
 sky130_fd_sc_hd__xnor2_2 _15486_ (.A(_12539_),
    .B(_12543_),
    .Y(_12545_));
 sky130_fd_sc_hd__xnor2_2 _15487_ (.A(_12510_),
    .B(_12545_),
    .Y(_12546_));
 sky130_fd_sc_hd__nand2_2 _15488_ (.A(\systolic_inst.B_outs[13][2] ),
    .B(\systolic_inst.A_outs[13][5] ),
    .Y(_12547_));
 sky130_fd_sc_hd__and4_2 _15489_ (.A(\systolic_inst.B_outs[13][3] ),
    .B(\systolic_inst.A_outs[13][3] ),
    .C(\systolic_inst.B_outs[13][4] ),
    .D(\systolic_inst.A_outs[13][4] ),
    .X(_12548_));
 sky130_fd_sc_hd__a22oi_2 _15490_ (.A1(\systolic_inst.A_outs[13][3] ),
    .A2(\systolic_inst.B_outs[13][4] ),
    .B1(\systolic_inst.A_outs[13][4] ),
    .B2(\systolic_inst.B_outs[13][3] ),
    .Y(_12549_));
 sky130_fd_sc_hd__or2_2 _15491_ (.A(_12548_),
    .B(_12549_),
    .X(_12550_));
 sky130_fd_sc_hd__xnor2_2 _15492_ (.A(_12547_),
    .B(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__nand2_2 _15493_ (.A(\systolic_inst.A_outs[13][2] ),
    .B(\systolic_inst.B_outs[13][5] ),
    .Y(_12552_));
 sky130_fd_sc_hd__and2b_2 _15494_ (.A_N(\systolic_inst.A_outs[13][0] ),
    .B(\systolic_inst.B_outs[13][7] ),
    .X(_12553_));
 sky130_fd_sc_hd__and3_2 _15495_ (.A(\systolic_inst.A_outs[13][1] ),
    .B(\systolic_inst.B_outs[13][6] ),
    .C(_12553_),
    .X(_12554_));
 sky130_fd_sc_hd__xnor2_2 _15496_ (.A(_12520_),
    .B(_12553_),
    .Y(_12555_));
 sky130_fd_sc_hd__xnor2_2 _15497_ (.A(_12552_),
    .B(_12555_),
    .Y(_12556_));
 sky130_fd_sc_hd__xnor2_2 _15498_ (.A(_12521_),
    .B(_12556_),
    .Y(_12557_));
 sky130_fd_sc_hd__nor2_2 _15499_ (.A(_12551_),
    .B(_12557_),
    .Y(_12558_));
 sky130_fd_sc_hd__xnor2_2 _15500_ (.A(_12551_),
    .B(_12557_),
    .Y(_12559_));
 sky130_fd_sc_hd__or2_2 _15501_ (.A(_12523_),
    .B(_12559_),
    .X(_12560_));
 sky130_fd_sc_hd__and2_2 _15502_ (.A(_12523_),
    .B(_12559_),
    .X(_12561_));
 sky130_fd_sc_hd__xor2_2 _15503_ (.A(_12523_),
    .B(_12559_),
    .X(_12562_));
 sky130_fd_sc_hd__xnor2_2 _15504_ (.A(_12546_),
    .B(_12562_),
    .Y(_12563_));
 sky130_fd_sc_hd__and2b_2 _15505_ (.A_N(_12525_),
    .B(_12527_),
    .X(_12564_));
 sky130_fd_sc_hd__nand2b_2 _15506_ (.A_N(_12564_),
    .B(_12563_),
    .Y(_12565_));
 sky130_fd_sc_hd__xnor2_2 _15507_ (.A(_12563_),
    .B(_12564_),
    .Y(_12566_));
 sky130_fd_sc_hd__nand2b_2 _15508_ (.A_N(_12538_),
    .B(_12566_),
    .Y(_12567_));
 sky130_fd_sc_hd__xnor2_2 _15509_ (.A(_12538_),
    .B(_12566_),
    .Y(_12568_));
 sky130_fd_sc_hd__and2b_2 _15510_ (.A_N(_12537_),
    .B(_12568_),
    .X(_12569_));
 sky130_fd_sc_hd__xnor2_2 _15511_ (.A(_12537_),
    .B(_12568_),
    .Y(_12570_));
 sky130_fd_sc_hd__a31o_2 _15512_ (.A1(_12502_),
    .A2(_12503_),
    .A3(_12535_),
    .B1(_12533_),
    .X(_12571_));
 sky130_fd_sc_hd__xor2_2 _15513_ (.A(_12570_),
    .B(_12571_),
    .X(_12572_));
 sky130_fd_sc_hd__mux2_1 _15514_ (.A0(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[7] ),
    .A1(_12572_),
    .S(\systolic_inst.ce_local ),
    .X(_01097_));
 sky130_fd_sc_hd__a21bo_2 _15515_ (.A1(_12510_),
    .A2(_12545_),
    .B1_N(_12544_),
    .X(_12573_));
 sky130_fd_sc_hd__a21bo_2 _15516_ (.A1(\systolic_inst.B_outs[13][7] ),
    .A2(_12540_),
    .B1_N(_12541_),
    .X(_12574_));
 sky130_fd_sc_hd__o21bai_2 _15517_ (.A1(_12547_),
    .A2(_12549_),
    .B1_N(_12548_),
    .Y(_12575_));
 sky130_fd_sc_hd__o21a_2 _15518_ (.A1(\systolic_inst.B_outs[13][0] ),
    .A2(\systolic_inst.B_outs[13][1] ),
    .B1(\systolic_inst.A_outs[13][7] ),
    .X(_12576_));
 sky130_fd_sc_hd__o21ai_2 _15519_ (.A1(\systolic_inst.B_outs[13][0] ),
    .A2(\systolic_inst.B_outs[13][1] ),
    .B1(\systolic_inst.A_outs[13][7] ),
    .Y(_12577_));
 sky130_fd_sc_hd__a21o_2 _15520_ (.A1(\systolic_inst.B_outs[13][0] ),
    .A2(\systolic_inst.B_outs[13][1] ),
    .B1(_12577_),
    .X(_12578_));
 sky130_fd_sc_hd__and2b_2 _15521_ (.A_N(_12578_),
    .B(_12575_),
    .X(_12579_));
 sky130_fd_sc_hd__xnor2_2 _15522_ (.A(_12575_),
    .B(_12578_),
    .Y(_12580_));
 sky130_fd_sc_hd__xnor2_2 _15523_ (.A(_12574_),
    .B(_12580_),
    .Y(_12581_));
 sky130_fd_sc_hd__and4_2 _15524_ (.A(\systolic_inst.B_outs[13][3] ),
    .B(\systolic_inst.B_outs[13][4] ),
    .C(\systolic_inst.A_outs[13][4] ),
    .D(\systolic_inst.A_outs[13][5] ),
    .X(_12582_));
 sky130_fd_sc_hd__a22oi_2 _15525_ (.A1(\systolic_inst.B_outs[13][4] ),
    .A2(\systolic_inst.A_outs[13][4] ),
    .B1(\systolic_inst.A_outs[13][5] ),
    .B2(\systolic_inst.B_outs[13][3] ),
    .Y(_12583_));
 sky130_fd_sc_hd__nor2_2 _15526_ (.A(_12582_),
    .B(_12583_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand2_2 _15527_ (.A(\systolic_inst.B_outs[13][2] ),
    .B(\systolic_inst.A_outs[13][6] ),
    .Y(_12585_));
 sky130_fd_sc_hd__xnor2_2 _15528_ (.A(_12584_),
    .B(_12585_),
    .Y(_12586_));
 sky130_fd_sc_hd__nand2_2 _15529_ (.A(\systolic_inst.A_outs[13][3] ),
    .B(\systolic_inst.B_outs[13][5] ),
    .Y(_12587_));
 sky130_fd_sc_hd__and4b_2 _15530_ (.A_N(\systolic_inst.A_outs[13][1] ),
    .B(\systolic_inst.A_outs[13][2] ),
    .C(\systolic_inst.B_outs[13][6] ),
    .D(\systolic_inst.B_outs[13][7] ),
    .X(_12588_));
 sky130_fd_sc_hd__a2bb2o_2 _15531_ (.A1_N(\systolic_inst.A_outs[13][1] ),
    .A2_N(_11272_),
    .B1(\systolic_inst.B_outs[13][6] ),
    .B2(\systolic_inst.A_outs[13][2] ),
    .X(_12589_));
 sky130_fd_sc_hd__and2b_2 _15532_ (.A_N(_12588_),
    .B(_12589_),
    .X(_12590_));
 sky130_fd_sc_hd__xnor2_2 _15533_ (.A(_12587_),
    .B(_12590_),
    .Y(_12591_));
 sky130_fd_sc_hd__a31o_2 _15534_ (.A1(\systolic_inst.A_outs[13][2] ),
    .A2(\systolic_inst.B_outs[13][5] ),
    .A3(_12555_),
    .B1(_12554_),
    .X(_12592_));
 sky130_fd_sc_hd__and2_2 _15535_ (.A(_12591_),
    .B(_12592_),
    .X(_12593_));
 sky130_fd_sc_hd__xor2_2 _15536_ (.A(_12591_),
    .B(_12592_),
    .X(_12594_));
 sky130_fd_sc_hd__xor2_2 _15537_ (.A(_12586_),
    .B(_12594_),
    .X(_12595_));
 sky130_fd_sc_hd__a21oi_2 _15538_ (.A1(_12521_),
    .A2(_12556_),
    .B1(_12558_),
    .Y(_12596_));
 sky130_fd_sc_hd__and2b_2 _15539_ (.A_N(_12596_),
    .B(_12595_),
    .X(_12597_));
 sky130_fd_sc_hd__xor2_2 _15540_ (.A(_12595_),
    .B(_12596_),
    .X(_12598_));
 sky130_fd_sc_hd__xor2_2 _15541_ (.A(_12581_),
    .B(_12598_),
    .X(_12599_));
 sky130_fd_sc_hd__o21a_2 _15542_ (.A1(_12546_),
    .A2(_12561_),
    .B1(_12560_),
    .X(_12600_));
 sky130_fd_sc_hd__and2b_2 _15543_ (.A_N(_12600_),
    .B(_12599_),
    .X(_12601_));
 sky130_fd_sc_hd__xnor2_2 _15544_ (.A(_12599_),
    .B(_12600_),
    .Y(_12602_));
 sky130_fd_sc_hd__xnor2_2 _15545_ (.A(_12573_),
    .B(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__and2_2 _15546_ (.A(_12565_),
    .B(_12567_),
    .X(_12604_));
 sky130_fd_sc_hd__nor2_2 _15547_ (.A(_12603_),
    .B(_12604_),
    .Y(_12605_));
 sky130_fd_sc_hd__xor2_2 _15548_ (.A(_12603_),
    .B(_12604_),
    .X(_12606_));
 sky130_fd_sc_hd__a21oi_2 _15549_ (.A1(_12570_),
    .A2(_12571_),
    .B1(_12569_),
    .Y(_12607_));
 sky130_fd_sc_hd__and2b_2 _15550_ (.A_N(_12607_),
    .B(_12606_),
    .X(_12608_));
 sky130_fd_sc_hd__xnor2_2 _15551_ (.A(_12606_),
    .B(_12607_),
    .Y(_12609_));
 sky130_fd_sc_hd__mux2_1 _15552_ (.A0(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[8] ),
    .A1(_12609_),
    .S(\systolic_inst.ce_local ),
    .X(_01098_));
 sky130_fd_sc_hd__a21o_2 _15553_ (.A1(_12573_),
    .A2(_12602_),
    .B1(_12601_),
    .X(_12610_));
 sky130_fd_sc_hd__a21o_2 _15554_ (.A1(_12574_),
    .A2(_12580_),
    .B1(_12579_),
    .X(_12611_));
 sky130_fd_sc_hd__o21ba_2 _15555_ (.A1(_12583_),
    .A2(_12585_),
    .B1_N(_12582_),
    .X(_12612_));
 sky130_fd_sc_hd__nor2_2 _15556_ (.A(_12577_),
    .B(_12612_),
    .Y(_12613_));
 sky130_fd_sc_hd__and2_2 _15557_ (.A(_12577_),
    .B(_12612_),
    .X(_12614_));
 sky130_fd_sc_hd__or2_2 _15558_ (.A(_12613_),
    .B(_12614_),
    .X(_12615_));
 sky130_fd_sc_hd__nand2_2 _15559_ (.A(\systolic_inst.B_outs[13][2] ),
    .B(\systolic_inst.A_outs[13][7] ),
    .Y(_12616_));
 sky130_fd_sc_hd__a22oi_2 _15560_ (.A1(\systolic_inst.B_outs[13][4] ),
    .A2(\systolic_inst.A_outs[13][5] ),
    .B1(\systolic_inst.A_outs[13][6] ),
    .B2(\systolic_inst.B_outs[13][3] ),
    .Y(_12617_));
 sky130_fd_sc_hd__and4_2 _15561_ (.A(\systolic_inst.B_outs[13][3] ),
    .B(\systolic_inst.B_outs[13][4] ),
    .C(\systolic_inst.A_outs[13][5] ),
    .D(\systolic_inst.A_outs[13][6] ),
    .X(_12618_));
 sky130_fd_sc_hd__nor2_2 _15562_ (.A(_12617_),
    .B(_12618_),
    .Y(_12619_));
 sky130_fd_sc_hd__xnor2_2 _15563_ (.A(_12616_),
    .B(_12619_),
    .Y(_12620_));
 sky130_fd_sc_hd__nand2_2 _15564_ (.A(\systolic_inst.A_outs[13][4] ),
    .B(\systolic_inst.B_outs[13][5] ),
    .Y(_12621_));
 sky130_fd_sc_hd__and4b_2 _15565_ (.A_N(\systolic_inst.A_outs[13][2] ),
    .B(\systolic_inst.A_outs[13][3] ),
    .C(\systolic_inst.B_outs[13][6] ),
    .D(\systolic_inst.B_outs[13][7] ),
    .X(_12622_));
 sky130_fd_sc_hd__o2bb2a_2 _15566_ (.A1_N(\systolic_inst.A_outs[13][3] ),
    .A2_N(\systolic_inst.B_outs[13][6] ),
    .B1(_11272_),
    .B2(\systolic_inst.A_outs[13][2] ),
    .X(_12623_));
 sky130_fd_sc_hd__nor2_2 _15567_ (.A(_12622_),
    .B(_12623_),
    .Y(_12624_));
 sky130_fd_sc_hd__xnor2_2 _15568_ (.A(_12621_),
    .B(_12624_),
    .Y(_12625_));
 sky130_fd_sc_hd__a31oi_2 _15569_ (.A1(\systolic_inst.A_outs[13][3] ),
    .A2(\systolic_inst.B_outs[13][5] ),
    .A3(_12589_),
    .B1(_12588_),
    .Y(_12626_));
 sky130_fd_sc_hd__nand2b_2 _15570_ (.A_N(_12626_),
    .B(_12625_),
    .Y(_12627_));
 sky130_fd_sc_hd__xnor2_2 _15571_ (.A(_12625_),
    .B(_12626_),
    .Y(_12628_));
 sky130_fd_sc_hd__xnor2_2 _15572_ (.A(_12620_),
    .B(_12628_),
    .Y(_12629_));
 sky130_fd_sc_hd__a21o_2 _15573_ (.A1(_12586_),
    .A2(_12594_),
    .B1(_12593_),
    .X(_12630_));
 sky130_fd_sc_hd__and2b_2 _15574_ (.A_N(_12629_),
    .B(_12630_),
    .X(_12631_));
 sky130_fd_sc_hd__xor2_2 _15575_ (.A(_12629_),
    .B(_12630_),
    .X(_12632_));
 sky130_fd_sc_hd__xor2_2 _15576_ (.A(_12615_),
    .B(_12632_),
    .X(_12633_));
 sky130_fd_sc_hd__o21ba_2 _15577_ (.A1(_12581_),
    .A2(_12598_),
    .B1_N(_12597_),
    .X(_12634_));
 sky130_fd_sc_hd__nand2b_2 _15578_ (.A_N(_12634_),
    .B(_12633_),
    .Y(_12635_));
 sky130_fd_sc_hd__xnor2_2 _15579_ (.A(_12633_),
    .B(_12634_),
    .Y(_12636_));
 sky130_fd_sc_hd__xnor2_2 _15580_ (.A(_12611_),
    .B(_12636_),
    .Y(_12637_));
 sky130_fd_sc_hd__nand2b_2 _15581_ (.A_N(_12610_),
    .B(_12637_),
    .Y(_12638_));
 sky130_fd_sc_hd__and2b_2 _15582_ (.A_N(_12637_),
    .B(_12610_),
    .X(_12639_));
 sky130_fd_sc_hd__xnor2_2 _15583_ (.A(_12610_),
    .B(_12637_),
    .Y(_12640_));
 sky130_fd_sc_hd__o21ai_2 _15584_ (.A1(_12605_),
    .A2(_12608_),
    .B1(_12640_),
    .Y(_12641_));
 sky130_fd_sc_hd__o31a_2 _15585_ (.A1(_12605_),
    .A2(_12608_),
    .A3(_12640_),
    .B1(\systolic_inst.ce_local ),
    .X(_12642_));
 sky130_fd_sc_hd__a22o_2 _15586_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[9] ),
    .B1(_12641_),
    .B2(_12642_),
    .X(_01099_));
 sky130_fd_sc_hd__o21ba_2 _15587_ (.A1(_12616_),
    .A2(_12617_),
    .B1_N(_12618_),
    .X(_12643_));
 sky130_fd_sc_hd__nor2_2 _15588_ (.A(_12577_),
    .B(_12643_),
    .Y(_12644_));
 sky130_fd_sc_hd__and2_2 _15589_ (.A(_12577_),
    .B(_12643_),
    .X(_12645_));
 sky130_fd_sc_hd__or2_2 _15590_ (.A(_12644_),
    .B(_12645_),
    .X(_12646_));
 sky130_fd_sc_hd__a22o_2 _15591_ (.A1(\systolic_inst.B_outs[13][4] ),
    .A2(\systolic_inst.A_outs[13][6] ),
    .B1(\systolic_inst.A_outs[13][7] ),
    .B2(\systolic_inst.B_outs[13][3] ),
    .X(_12647_));
 sky130_fd_sc_hd__and3_2 _15592_ (.A(\systolic_inst.B_outs[13][3] ),
    .B(\systolic_inst.B_outs[13][4] ),
    .C(\systolic_inst.A_outs[13][7] ),
    .X(_12648_));
 sky130_fd_sc_hd__a21bo_2 _15593_ (.A1(\systolic_inst.A_outs[13][6] ),
    .A2(_12648_),
    .B1_N(_12647_),
    .X(_12649_));
 sky130_fd_sc_hd__xor2_2 _15594_ (.A(_12616_),
    .B(_12649_),
    .X(_12650_));
 sky130_fd_sc_hd__nand2_2 _15595_ (.A(\systolic_inst.B_outs[13][5] ),
    .B(\systolic_inst.A_outs[13][5] ),
    .Y(_12651_));
 sky130_fd_sc_hd__and4b_2 _15596_ (.A_N(\systolic_inst.A_outs[13][3] ),
    .B(\systolic_inst.A_outs[13][4] ),
    .C(\systolic_inst.B_outs[13][6] ),
    .D(\systolic_inst.B_outs[13][7] ),
    .X(_12652_));
 sky130_fd_sc_hd__o2bb2a_2 _15597_ (.A1_N(\systolic_inst.A_outs[13][4] ),
    .A2_N(\systolic_inst.B_outs[13][6] ),
    .B1(_11272_),
    .B2(\systolic_inst.A_outs[13][3] ),
    .X(_12653_));
 sky130_fd_sc_hd__nor2_2 _15598_ (.A(_12652_),
    .B(_12653_),
    .Y(_12654_));
 sky130_fd_sc_hd__xnor2_2 _15599_ (.A(_12651_),
    .B(_12654_),
    .Y(_12655_));
 sky130_fd_sc_hd__o21ba_2 _15600_ (.A1(_12621_),
    .A2(_12623_),
    .B1_N(_12622_),
    .X(_12656_));
 sky130_fd_sc_hd__nand2b_2 _15601_ (.A_N(_12656_),
    .B(_12655_),
    .Y(_12657_));
 sky130_fd_sc_hd__xnor2_2 _15602_ (.A(_12655_),
    .B(_12656_),
    .Y(_12658_));
 sky130_fd_sc_hd__nand2_2 _15603_ (.A(_12650_),
    .B(_12658_),
    .Y(_12659_));
 sky130_fd_sc_hd__or2_2 _15604_ (.A(_12650_),
    .B(_12658_),
    .X(_12660_));
 sky130_fd_sc_hd__nand2_2 _15605_ (.A(_12659_),
    .B(_12660_),
    .Y(_12661_));
 sky130_fd_sc_hd__a21bo_2 _15606_ (.A1(_12620_),
    .A2(_12628_),
    .B1_N(_12627_),
    .X(_12662_));
 sky130_fd_sc_hd__nand2b_2 _15607_ (.A_N(_12661_),
    .B(_12662_),
    .Y(_12663_));
 sky130_fd_sc_hd__xor2_2 _15608_ (.A(_12661_),
    .B(_12662_),
    .X(_12664_));
 sky130_fd_sc_hd__xor2_2 _15609_ (.A(_12646_),
    .B(_12664_),
    .X(_12665_));
 sky130_fd_sc_hd__o21ba_2 _15610_ (.A1(_12615_),
    .A2(_12632_),
    .B1_N(_12631_),
    .X(_12666_));
 sky130_fd_sc_hd__nand2b_2 _15611_ (.A_N(_12666_),
    .B(_12665_),
    .Y(_12667_));
 sky130_fd_sc_hd__xnor2_2 _15612_ (.A(_12665_),
    .B(_12666_),
    .Y(_12668_));
 sky130_fd_sc_hd__nand2_2 _15613_ (.A(_12613_),
    .B(_12668_),
    .Y(_12669_));
 sky130_fd_sc_hd__xnor2_2 _15614_ (.A(_12613_),
    .B(_12668_),
    .Y(_12670_));
 sky130_fd_sc_hd__a21boi_2 _15615_ (.A1(_12611_),
    .A2(_12636_),
    .B1_N(_12635_),
    .Y(_12671_));
 sky130_fd_sc_hd__or2_2 _15616_ (.A(_12670_),
    .B(_12671_),
    .X(_12672_));
 sky130_fd_sc_hd__nand2_2 _15617_ (.A(_12670_),
    .B(_12671_),
    .Y(_12673_));
 sky130_fd_sc_hd__and2_2 _15618_ (.A(_12672_),
    .B(_12673_),
    .X(_12674_));
 sky130_fd_sc_hd__a21o_2 _15619_ (.A1(_12605_),
    .A2(_12638_),
    .B1(_12639_),
    .X(_12675_));
 sky130_fd_sc_hd__a21o_2 _15620_ (.A1(_12608_),
    .A2(_12640_),
    .B1(_12675_),
    .X(_12676_));
 sky130_fd_sc_hd__or2_2 _15621_ (.A(_12674_),
    .B(_12676_),
    .X(_12677_));
 sky130_fd_sc_hd__nand2_2 _15622_ (.A(_12674_),
    .B(_12676_),
    .Y(_12678_));
 sky130_fd_sc_hd__and2_2 _15623_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[10] ),
    .X(_12679_));
 sky130_fd_sc_hd__a31o_2 _15624_ (.A1(\systolic_inst.ce_local ),
    .A2(_12677_),
    .A3(_12678_),
    .B1(_12679_),
    .X(_01100_));
 sky130_fd_sc_hd__or2_2 _15625_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[11] ),
    .X(_12680_));
 sky130_fd_sc_hd__o2bb2a_2 _15626_ (.A1_N(\systolic_inst.A_outs[13][6] ),
    .A2_N(_12648_),
    .B1(_12649_),
    .B2(_12616_),
    .X(_12681_));
 sky130_fd_sc_hd__or2_2 _15627_ (.A(_12577_),
    .B(_12681_),
    .X(_12682_));
 sky130_fd_sc_hd__nand2_2 _15628_ (.A(_12577_),
    .B(_12681_),
    .Y(_12683_));
 sky130_fd_sc_hd__nand2_2 _15629_ (.A(_12682_),
    .B(_12683_),
    .Y(_12684_));
 sky130_fd_sc_hd__or2_2 _15630_ (.A(\systolic_inst.B_outs[13][3] ),
    .B(\systolic_inst.B_outs[13][4] ),
    .X(_12685_));
 sky130_fd_sc_hd__and3b_2 _15631_ (.A_N(_12648_),
    .B(_12685_),
    .C(\systolic_inst.A_outs[13][7] ),
    .X(_12686_));
 sky130_fd_sc_hd__xnor2_2 _15632_ (.A(_12616_),
    .B(_12686_),
    .Y(_12687_));
 sky130_fd_sc_hd__nand2_2 _15633_ (.A(\systolic_inst.B_outs[13][5] ),
    .B(\systolic_inst.A_outs[13][6] ),
    .Y(_12688_));
 sky130_fd_sc_hd__and4b_2 _15634_ (.A_N(\systolic_inst.A_outs[13][4] ),
    .B(\systolic_inst.A_outs[13][5] ),
    .C(\systolic_inst.B_outs[13][6] ),
    .D(\systolic_inst.B_outs[13][7] ),
    .X(_12689_));
 sky130_fd_sc_hd__o2bb2a_2 _15635_ (.A1_N(\systolic_inst.A_outs[13][5] ),
    .A2_N(\systolic_inst.B_outs[13][6] ),
    .B1(_11272_),
    .B2(\systolic_inst.A_outs[13][4] ),
    .X(_12690_));
 sky130_fd_sc_hd__or2_2 _15636_ (.A(_12689_),
    .B(_12690_),
    .X(_12691_));
 sky130_fd_sc_hd__xor2_2 _15637_ (.A(_12688_),
    .B(_12691_),
    .X(_12692_));
 sky130_fd_sc_hd__o21ba_2 _15638_ (.A1(_12651_),
    .A2(_12653_),
    .B1_N(_12652_),
    .X(_12693_));
 sky130_fd_sc_hd__nand2b_2 _15639_ (.A_N(_12693_),
    .B(_12692_),
    .Y(_12694_));
 sky130_fd_sc_hd__xnor2_2 _15640_ (.A(_12692_),
    .B(_12693_),
    .Y(_12695_));
 sky130_fd_sc_hd__nand2_2 _15641_ (.A(_12687_),
    .B(_12695_),
    .Y(_12696_));
 sky130_fd_sc_hd__xnor2_2 _15642_ (.A(_12687_),
    .B(_12695_),
    .Y(_12697_));
 sky130_fd_sc_hd__a21o_2 _15643_ (.A1(_12657_),
    .A2(_12659_),
    .B1(_12697_),
    .X(_12698_));
 sky130_fd_sc_hd__nand3_2 _15644_ (.A(_12657_),
    .B(_12659_),
    .C(_12697_),
    .Y(_12699_));
 sky130_fd_sc_hd__nand2_2 _15645_ (.A(_12698_),
    .B(_12699_),
    .Y(_12700_));
 sky130_fd_sc_hd__xor2_2 _15646_ (.A(_12684_),
    .B(_12700_),
    .X(_12701_));
 sky130_fd_sc_hd__o21a_2 _15647_ (.A1(_12646_),
    .A2(_12664_),
    .B1(_12663_),
    .X(_12702_));
 sky130_fd_sc_hd__and2b_2 _15648_ (.A_N(_12702_),
    .B(_12701_),
    .X(_12703_));
 sky130_fd_sc_hd__and2b_2 _15649_ (.A_N(_12701_),
    .B(_12702_),
    .X(_12704_));
 sky130_fd_sc_hd__nor2_2 _15650_ (.A(_12703_),
    .B(_12704_),
    .Y(_12705_));
 sky130_fd_sc_hd__xnor2_2 _15651_ (.A(_12644_),
    .B(_12705_),
    .Y(_12706_));
 sky130_fd_sc_hd__and3_2 _15652_ (.A(_12667_),
    .B(_12669_),
    .C(_12706_),
    .X(_12707_));
 sky130_fd_sc_hd__a21o_2 _15653_ (.A1(_12667_),
    .A2(_12669_),
    .B1(_12706_),
    .X(_12708_));
 sky130_fd_sc_hd__and2b_2 _15654_ (.A_N(_12707_),
    .B(_12708_),
    .X(_12709_));
 sky130_fd_sc_hd__a21oi_2 _15655_ (.A1(_12672_),
    .A2(_12678_),
    .B1(_12709_),
    .Y(_12710_));
 sky130_fd_sc_hd__and3_2 _15656_ (.A(_12672_),
    .B(_12678_),
    .C(_12709_),
    .X(_12711_));
 sky130_fd_sc_hd__o31a_2 _15657_ (.A1(_11258_),
    .A2(_12710_),
    .A3(_12711_),
    .B1(_12680_),
    .X(_01101_));
 sky130_fd_sc_hd__a31o_2 _15658_ (.A1(\systolic_inst.B_outs[13][2] ),
    .A2(\systolic_inst.A_outs[13][7] ),
    .A3(_12685_),
    .B1(_12648_),
    .X(_12712_));
 sky130_fd_sc_hd__or2_2 _15659_ (.A(_12576_),
    .B(_12712_),
    .X(_12713_));
 sky130_fd_sc_hd__nand2_2 _15660_ (.A(_12576_),
    .B(_12712_),
    .Y(_12714_));
 sky130_fd_sc_hd__nand2_2 _15661_ (.A(_12713_),
    .B(_12714_),
    .Y(_12715_));
 sky130_fd_sc_hd__inv_2 _15662_ (.A(_12715_),
    .Y(_12716_));
 sky130_fd_sc_hd__o2bb2a_2 _15663_ (.A1_N(\systolic_inst.B_outs[13][6] ),
    .A2_N(\systolic_inst.A_outs[13][6] ),
    .B1(_11272_),
    .B2(\systolic_inst.A_outs[13][5] ),
    .X(_12717_));
 sky130_fd_sc_hd__and4b_2 _15664_ (.A_N(\systolic_inst.A_outs[13][5] ),
    .B(\systolic_inst.B_outs[13][6] ),
    .C(\systolic_inst.A_outs[13][6] ),
    .D(\systolic_inst.B_outs[13][7] ),
    .X(_12718_));
 sky130_fd_sc_hd__nor2_2 _15665_ (.A(_12717_),
    .B(_12718_),
    .Y(_12719_));
 sky130_fd_sc_hd__nand2_2 _15666_ (.A(\systolic_inst.B_outs[13][5] ),
    .B(\systolic_inst.A_outs[13][7] ),
    .Y(_12720_));
 sky130_fd_sc_hd__and3_2 _15667_ (.A(\systolic_inst.B_outs[13][5] ),
    .B(\systolic_inst.A_outs[13][7] ),
    .C(_12719_),
    .X(_12721_));
 sky130_fd_sc_hd__xnor2_2 _15668_ (.A(_12719_),
    .B(_12720_),
    .Y(_12722_));
 sky130_fd_sc_hd__o21ba_2 _15669_ (.A1(_12688_),
    .A2(_12690_),
    .B1_N(_12689_),
    .X(_12723_));
 sky130_fd_sc_hd__nand2b_2 _15670_ (.A_N(_12723_),
    .B(_12722_),
    .Y(_12724_));
 sky130_fd_sc_hd__xnor2_2 _15671_ (.A(_12722_),
    .B(_12723_),
    .Y(_12725_));
 sky130_fd_sc_hd__xnor2_2 _15672_ (.A(_12687_),
    .B(_12725_),
    .Y(_12726_));
 sky130_fd_sc_hd__a21o_2 _15673_ (.A1(_12694_),
    .A2(_12696_),
    .B1(_12726_),
    .X(_12727_));
 sky130_fd_sc_hd__nand3_2 _15674_ (.A(_12694_),
    .B(_12696_),
    .C(_12726_),
    .Y(_12728_));
 sky130_fd_sc_hd__nand2_2 _15675_ (.A(_12727_),
    .B(_12728_),
    .Y(_12729_));
 sky130_fd_sc_hd__xnor2_2 _15676_ (.A(_12716_),
    .B(_12729_),
    .Y(_12730_));
 sky130_fd_sc_hd__o21a_2 _15677_ (.A1(_12684_),
    .A2(_12700_),
    .B1(_12698_),
    .X(_12731_));
 sky130_fd_sc_hd__and2b_2 _15678_ (.A_N(_12731_),
    .B(_12730_),
    .X(_12732_));
 sky130_fd_sc_hd__and2b_2 _15679_ (.A_N(_12730_),
    .B(_12731_),
    .X(_12733_));
 sky130_fd_sc_hd__nor2_2 _15680_ (.A(_12732_),
    .B(_12733_),
    .Y(_12734_));
 sky130_fd_sc_hd__and2b_2 _15681_ (.A_N(_12682_),
    .B(_12734_),
    .X(_12735_));
 sky130_fd_sc_hd__xor2_2 _15682_ (.A(_12682_),
    .B(_12734_),
    .X(_12736_));
 sky130_fd_sc_hd__a21oi_2 _15683_ (.A1(_12644_),
    .A2(_12705_),
    .B1(_12703_),
    .Y(_12737_));
 sky130_fd_sc_hd__or2_2 _15684_ (.A(_12736_),
    .B(_12737_),
    .X(_12738_));
 sky130_fd_sc_hd__inv_2 _15685_ (.A(_12738_),
    .Y(_12739_));
 sky130_fd_sc_hd__nand2_2 _15686_ (.A(_12736_),
    .B(_12737_),
    .Y(_12740_));
 sky130_fd_sc_hd__nand2_2 _15687_ (.A(_12738_),
    .B(_12740_),
    .Y(_12741_));
 sky130_fd_sc_hd__a31o_2 _15688_ (.A1(_12672_),
    .A2(_12678_),
    .A3(_12708_),
    .B1(_12707_),
    .X(_12742_));
 sky130_fd_sc_hd__nand2_2 _15689_ (.A(_12741_),
    .B(_12742_),
    .Y(_12743_));
 sky130_fd_sc_hd__a311oi_2 _15690_ (.A1(_12672_),
    .A2(_12678_),
    .A3(_12708_),
    .B1(_12741_),
    .C1(_12707_),
    .Y(_12744_));
 sky130_fd_sc_hd__nor2_2 _15691_ (.A(_11258_),
    .B(_12744_),
    .Y(_12745_));
 sky130_fd_sc_hd__a22o_2 _15692_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[12] ),
    .B1(_12743_),
    .B2(_12745_),
    .X(_01102_));
 sky130_fd_sc_hd__nand2_2 _15693_ (.A(\systolic_inst.B_outs[13][6] ),
    .B(\systolic_inst.A_outs[13][7] ),
    .Y(_12746_));
 sky130_fd_sc_hd__nor2_2 _15694_ (.A(\systolic_inst.A_outs[13][6] ),
    .B(_11272_),
    .Y(_12747_));
 sky130_fd_sc_hd__xnor2_2 _15695_ (.A(_12746_),
    .B(_12747_),
    .Y(_12748_));
 sky130_fd_sc_hd__nand2b_2 _15696_ (.A_N(_12720_),
    .B(_12748_),
    .Y(_12749_));
 sky130_fd_sc_hd__xnor2_2 _15697_ (.A(_12720_),
    .B(_12748_),
    .Y(_12750_));
 sky130_fd_sc_hd__o21ai_2 _15698_ (.A1(_12718_),
    .A2(_12721_),
    .B1(_12750_),
    .Y(_12751_));
 sky130_fd_sc_hd__or3_2 _15699_ (.A(_12718_),
    .B(_12721_),
    .C(_12750_),
    .X(_12752_));
 sky130_fd_sc_hd__and2_2 _15700_ (.A(_12751_),
    .B(_12752_),
    .X(_12753_));
 sky130_fd_sc_hd__nand2_2 _15701_ (.A(_12687_),
    .B(_12753_),
    .Y(_12754_));
 sky130_fd_sc_hd__or2_2 _15702_ (.A(_12687_),
    .B(_12753_),
    .X(_12755_));
 sky130_fd_sc_hd__nand2_2 _15703_ (.A(_12754_),
    .B(_12755_),
    .Y(_12756_));
 sky130_fd_sc_hd__a21bo_2 _15704_ (.A1(_12687_),
    .A2(_12725_),
    .B1_N(_12724_),
    .X(_12757_));
 sky130_fd_sc_hd__nand2b_2 _15705_ (.A_N(_12756_),
    .B(_12757_),
    .Y(_12758_));
 sky130_fd_sc_hd__xor2_2 _15706_ (.A(_12756_),
    .B(_12757_),
    .X(_12759_));
 sky130_fd_sc_hd__xnor2_2 _15707_ (.A(_12716_),
    .B(_12759_),
    .Y(_12760_));
 sky130_fd_sc_hd__o21a_2 _15708_ (.A1(_12715_),
    .A2(_12729_),
    .B1(_12727_),
    .X(_12761_));
 sky130_fd_sc_hd__and2b_2 _15709_ (.A_N(_12761_),
    .B(_12760_),
    .X(_12762_));
 sky130_fd_sc_hd__and2b_2 _15710_ (.A_N(_12760_),
    .B(_12761_),
    .X(_12763_));
 sky130_fd_sc_hd__nor2_2 _15711_ (.A(_12762_),
    .B(_12763_),
    .Y(_12764_));
 sky130_fd_sc_hd__xnor2_2 _15712_ (.A(_12714_),
    .B(_12764_),
    .Y(_12765_));
 sky130_fd_sc_hd__nor3_2 _15713_ (.A(_12732_),
    .B(_12735_),
    .C(_12765_),
    .Y(_12766_));
 sky130_fd_sc_hd__o21ai_2 _15714_ (.A1(_12732_),
    .A2(_12735_),
    .B1(_12765_),
    .Y(_12767_));
 sky130_fd_sc_hd__and2b_2 _15715_ (.A_N(_12766_),
    .B(_12767_),
    .X(_12768_));
 sky130_fd_sc_hd__or3_2 _15716_ (.A(_12739_),
    .B(_12744_),
    .C(_12768_),
    .X(_12769_));
 sky130_fd_sc_hd__o21ai_2 _15717_ (.A1(_12739_),
    .A2(_12744_),
    .B1(_12768_),
    .Y(_12770_));
 sky130_fd_sc_hd__and3_2 _15718_ (.A(\systolic_inst.ce_local ),
    .B(_12769_),
    .C(_12770_),
    .X(_12771_));
 sky130_fd_sc_hd__a21o_2 _15719_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[13] ),
    .B1(_12771_),
    .X(_01103_));
 sky130_fd_sc_hd__o211ai_2 _15720_ (.A1(_11272_),
    .A2(\systolic_inst.A_outs[13][7] ),
    .B1(_12720_),
    .C1(_12746_),
    .Y(_12772_));
 sky130_fd_sc_hd__o311a_2 _15721_ (.A1(\systolic_inst.A_outs[13][6] ),
    .A2(_11272_),
    .A3(_12746_),
    .B1(_12749_),
    .C1(_12772_),
    .X(_12773_));
 sky130_fd_sc_hd__a31o_2 _15722_ (.A1(\systolic_inst.B_outs[13][5] ),
    .A2(\systolic_inst.B_outs[13][6] ),
    .A3(\systolic_inst.A_outs[13][7] ),
    .B1(_12773_),
    .X(_12774_));
 sky130_fd_sc_hd__nor2_2 _15723_ (.A(_12687_),
    .B(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__and2_2 _15724_ (.A(_12687_),
    .B(_12774_),
    .X(_12776_));
 sky130_fd_sc_hd__or2_2 _15725_ (.A(_12775_),
    .B(_12776_),
    .X(_12777_));
 sky130_fd_sc_hd__a21oi_2 _15726_ (.A1(_12751_),
    .A2(_12754_),
    .B1(_12777_),
    .Y(_12778_));
 sky130_fd_sc_hd__and3_2 _15727_ (.A(_12751_),
    .B(_12754_),
    .C(_12777_),
    .X(_12779_));
 sky130_fd_sc_hd__nor2_2 _15728_ (.A(_12778_),
    .B(_12779_),
    .Y(_12780_));
 sky130_fd_sc_hd__xnor2_2 _15729_ (.A(_12715_),
    .B(_12780_),
    .Y(_12781_));
 sky130_fd_sc_hd__o21a_2 _15730_ (.A1(_12715_),
    .A2(_12759_),
    .B1(_12758_),
    .X(_12782_));
 sky130_fd_sc_hd__and2b_2 _15731_ (.A_N(_12782_),
    .B(_12781_),
    .X(_12783_));
 sky130_fd_sc_hd__and2b_2 _15732_ (.A_N(_12781_),
    .B(_12782_),
    .X(_12784_));
 sky130_fd_sc_hd__nor2_2 _15733_ (.A(_12783_),
    .B(_12784_),
    .Y(_12785_));
 sky130_fd_sc_hd__xnor2_2 _15734_ (.A(_12714_),
    .B(_12785_),
    .Y(_12786_));
 sky130_fd_sc_hd__o21ba_2 _15735_ (.A1(_12714_),
    .A2(_12763_),
    .B1_N(_12762_),
    .X(_12787_));
 sky130_fd_sc_hd__nand2b_2 _15736_ (.A_N(_12787_),
    .B(_12786_),
    .Y(_12788_));
 sky130_fd_sc_hd__xnor2_2 _15737_ (.A(_12786_),
    .B(_12787_),
    .Y(_12789_));
 sky130_fd_sc_hd__o21ai_2 _15738_ (.A1(_12738_),
    .A2(_12766_),
    .B1(_12767_),
    .Y(_12790_));
 sky130_fd_sc_hd__a21o_2 _15739_ (.A1(_12744_),
    .A2(_12768_),
    .B1(_12790_),
    .X(_12791_));
 sky130_fd_sc_hd__nand2_2 _15740_ (.A(_12789_),
    .B(_12791_),
    .Y(_12792_));
 sky130_fd_sc_hd__xor2_2 _15741_ (.A(_12789_),
    .B(_12791_),
    .X(_12793_));
 sky130_fd_sc_hd__mux2_1 _15742_ (.A0(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[14] ),
    .A1(_12793_),
    .S(\systolic_inst.ce_local ),
    .X(_01104_));
 sky130_fd_sc_hd__a31oi_2 _15743_ (.A1(_12576_),
    .A2(_12712_),
    .A3(_12785_),
    .B1(_12783_),
    .Y(_12794_));
 sky130_fd_sc_hd__a21oi_2 _15744_ (.A1(_12716_),
    .A2(_12780_),
    .B1(_12778_),
    .Y(_12795_));
 sky130_fd_sc_hd__xnor2_2 _15745_ (.A(_12713_),
    .B(_12775_),
    .Y(_12796_));
 sky130_fd_sc_hd__xnor2_2 _15746_ (.A(_12795_),
    .B(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__xnor2_2 _15747_ (.A(_12794_),
    .B(_12797_),
    .Y(_12798_));
 sky130_fd_sc_hd__and3_2 _15748_ (.A(\systolic_inst.ce_local ),
    .B(_12788_),
    .C(_12798_),
    .X(_12799_));
 sky130_fd_sc_hd__a22o_2 _15749_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B1(_12792_),
    .B2(_12799_),
    .X(_01105_));
 sky130_fd_sc_hd__a21o_2 _15750_ (.A1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[13][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_12800_));
 sky130_fd_sc_hd__a21oi_2 _15751_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[13][0] ),
    .Y(_12801_));
 sky130_fd_sc_hd__a21oi_2 _15752_ (.A1(\systolic_inst.ce_local ),
    .A2(_12800_),
    .B1(_12801_),
    .Y(_01106_));
 sky130_fd_sc_hd__and2_2 _15753_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[13][1] ),
    .X(_12802_));
 sky130_fd_sc_hd__nand2_2 _15754_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[13][1] ),
    .Y(_12803_));
 sky130_fd_sc_hd__or2_2 _15755_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[13][1] ),
    .X(_12804_));
 sky130_fd_sc_hd__and4_2 _15756_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[13][0] ),
    .C(_12803_),
    .D(_12804_),
    .X(_12805_));
 sky130_fd_sc_hd__inv_2 _15757_ (.A(_12805_),
    .Y(_12806_));
 sky130_fd_sc_hd__a22o_2 _15758_ (.A1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[13][0] ),
    .B1(_12803_),
    .B2(_12804_),
    .X(_12807_));
 sky130_fd_sc_hd__a32o_2 _15759_ (.A1(_11712_),
    .A2(_12806_),
    .A3(_12807_),
    .B1(\systolic_inst.acc_wires[13][1] ),
    .B2(_11258_),
    .X(_01107_));
 sky130_fd_sc_hd__nand2_2 _15760_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[13][2] ),
    .Y(_12808_));
 sky130_fd_sc_hd__or2_2 _15761_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[13][2] ),
    .X(_12809_));
 sky130_fd_sc_hd__a31o_2 _15762_ (.A1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[13][0] ),
    .A3(_12804_),
    .B1(_12802_),
    .X(_12810_));
 sky130_fd_sc_hd__a21o_2 _15763_ (.A1(_12808_),
    .A2(_12809_),
    .B1(_12810_),
    .X(_12811_));
 sky130_fd_sc_hd__and3_2 _15764_ (.A(_12808_),
    .B(_12809_),
    .C(_12810_),
    .X(_12812_));
 sky130_fd_sc_hd__inv_2 _15765_ (.A(_12812_),
    .Y(_12813_));
 sky130_fd_sc_hd__a32o_2 _15766_ (.A1(_11712_),
    .A2(_12811_),
    .A3(_12813_),
    .B1(\systolic_inst.acc_wires[13][2] ),
    .B2(_11258_),
    .X(_01108_));
 sky130_fd_sc_hd__nand2_2 _15767_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[13][3] ),
    .Y(_12814_));
 sky130_fd_sc_hd__or2_2 _15768_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[13][3] ),
    .X(_12815_));
 sky130_fd_sc_hd__a21bo_2 _15769_ (.A1(_12809_),
    .A2(_12810_),
    .B1_N(_12808_),
    .X(_12816_));
 sky130_fd_sc_hd__a21o_2 _15770_ (.A1(_12814_),
    .A2(_12815_),
    .B1(_12816_),
    .X(_12817_));
 sky130_fd_sc_hd__and3_2 _15771_ (.A(_12814_),
    .B(_12815_),
    .C(_12816_),
    .X(_12818_));
 sky130_fd_sc_hd__inv_2 _15772_ (.A(_12818_),
    .Y(_12819_));
 sky130_fd_sc_hd__a32o_2 _15773_ (.A1(_11712_),
    .A2(_12817_),
    .A3(_12819_),
    .B1(\systolic_inst.acc_wires[13][3] ),
    .B2(_11258_),
    .X(_01109_));
 sky130_fd_sc_hd__nand2_2 _15774_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[13][4] ),
    .Y(_12820_));
 sky130_fd_sc_hd__or2_2 _15775_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[13][4] ),
    .X(_12821_));
 sky130_fd_sc_hd__a21bo_2 _15776_ (.A1(_12815_),
    .A2(_12816_),
    .B1_N(_12814_),
    .X(_12822_));
 sky130_fd_sc_hd__a21o_2 _15777_ (.A1(_12820_),
    .A2(_12821_),
    .B1(_12822_),
    .X(_12823_));
 sky130_fd_sc_hd__and3_2 _15778_ (.A(_12820_),
    .B(_12821_),
    .C(_12822_),
    .X(_12824_));
 sky130_fd_sc_hd__inv_2 _15779_ (.A(_12824_),
    .Y(_12825_));
 sky130_fd_sc_hd__a32o_2 _15780_ (.A1(_11712_),
    .A2(_12823_),
    .A3(_12825_),
    .B1(\systolic_inst.acc_wires[13][4] ),
    .B2(_11258_),
    .X(_01110_));
 sky130_fd_sc_hd__nand2_2 _15781_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[13][5] ),
    .Y(_12826_));
 sky130_fd_sc_hd__or2_2 _15782_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[13][5] ),
    .X(_12827_));
 sky130_fd_sc_hd__a21bo_2 _15783_ (.A1(_12821_),
    .A2(_12822_),
    .B1_N(_12820_),
    .X(_12828_));
 sky130_fd_sc_hd__a21o_2 _15784_ (.A1(_12826_),
    .A2(_12827_),
    .B1(_12828_),
    .X(_12829_));
 sky130_fd_sc_hd__and3_2 _15785_ (.A(_12826_),
    .B(_12827_),
    .C(_12828_),
    .X(_12830_));
 sky130_fd_sc_hd__inv_2 _15786_ (.A(_12830_),
    .Y(_12831_));
 sky130_fd_sc_hd__a32o_2 _15787_ (.A1(_11712_),
    .A2(_12829_),
    .A3(_12831_),
    .B1(\systolic_inst.acc_wires[13][5] ),
    .B2(_11258_),
    .X(_01111_));
 sky130_fd_sc_hd__nand2_2 _15788_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[13][6] ),
    .Y(_12832_));
 sky130_fd_sc_hd__or2_2 _15789_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[13][6] ),
    .X(_12833_));
 sky130_fd_sc_hd__a21bo_2 _15790_ (.A1(_12827_),
    .A2(_12828_),
    .B1_N(_12826_),
    .X(_12834_));
 sky130_fd_sc_hd__a21o_2 _15791_ (.A1(_12832_),
    .A2(_12833_),
    .B1(_12834_),
    .X(_12835_));
 sky130_fd_sc_hd__and3_2 _15792_ (.A(_12832_),
    .B(_12833_),
    .C(_12834_),
    .X(_12836_));
 sky130_fd_sc_hd__inv_2 _15793_ (.A(_12836_),
    .Y(_12837_));
 sky130_fd_sc_hd__a32o_2 _15794_ (.A1(_11712_),
    .A2(_12835_),
    .A3(_12837_),
    .B1(\systolic_inst.acc_wires[13][6] ),
    .B2(_11258_),
    .X(_01112_));
 sky130_fd_sc_hd__nand2_2 _15795_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[13][7] ),
    .Y(_12838_));
 sky130_fd_sc_hd__or2_2 _15796_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[13][7] ),
    .X(_12839_));
 sky130_fd_sc_hd__a21bo_2 _15797_ (.A1(_12833_),
    .A2(_12834_),
    .B1_N(_12832_),
    .X(_12840_));
 sky130_fd_sc_hd__a21o_2 _15798_ (.A1(_12838_),
    .A2(_12839_),
    .B1(_12840_),
    .X(_12841_));
 sky130_fd_sc_hd__nand3_2 _15799_ (.A(_12838_),
    .B(_12839_),
    .C(_12840_),
    .Y(_12842_));
 sky130_fd_sc_hd__a32o_2 _15800_ (.A1(_11712_),
    .A2(_12841_),
    .A3(_12842_),
    .B1(\systolic_inst.acc_wires[13][7] ),
    .B2(_11258_),
    .X(_01113_));
 sky130_fd_sc_hd__a21bo_2 _15801_ (.A1(_12839_),
    .A2(_12840_),
    .B1_N(_12838_),
    .X(_12843_));
 sky130_fd_sc_hd__xor2_2 _15802_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[13][8] ),
    .X(_12844_));
 sky130_fd_sc_hd__and2_2 _15803_ (.A(_12843_),
    .B(_12844_),
    .X(_12845_));
 sky130_fd_sc_hd__o21ai_2 _15804_ (.A1(_12843_),
    .A2(_12844_),
    .B1(_11712_),
    .Y(_12846_));
 sky130_fd_sc_hd__a2bb2o_2 _15805_ (.A1_N(_12846_),
    .A2_N(_12845_),
    .B1(\systolic_inst.acc_wires[13][8] ),
    .B2(_11258_),
    .X(_01114_));
 sky130_fd_sc_hd__xor2_2 _15806_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[13][9] ),
    .X(_12847_));
 sky130_fd_sc_hd__a211o_2 _15807_ (.A1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[13][8] ),
    .B1(_12845_),
    .C1(_12847_),
    .X(_12848_));
 sky130_fd_sc_hd__nand2_2 _15808_ (.A(_12844_),
    .B(_12847_),
    .Y(_12849_));
 sky130_fd_sc_hd__nand2_2 _15809_ (.A(_12845_),
    .B(_12847_),
    .Y(_12850_));
 sky130_fd_sc_hd__and3_2 _15810_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[13][8] ),
    .C(_12847_),
    .X(_12851_));
 sky130_fd_sc_hd__nor2_2 _15811_ (.A(_11713_),
    .B(_12851_),
    .Y(_12852_));
 sky130_fd_sc_hd__a32o_2 _15812_ (.A1(_12848_),
    .A2(_12850_),
    .A3(_12852_),
    .B1(\systolic_inst.acc_wires[13][9] ),
    .B2(_11258_),
    .X(_01115_));
 sky130_fd_sc_hd__nand2_2 _15813_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[13][10] ),
    .Y(_12853_));
 sky130_fd_sc_hd__or2_2 _15814_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[13][10] ),
    .X(_12854_));
 sky130_fd_sc_hd__and2_2 _15815_ (.A(_12853_),
    .B(_12854_),
    .X(_12855_));
 sky130_fd_sc_hd__a21oi_2 _15816_ (.A1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[13][9] ),
    .B1(_12851_),
    .Y(_12856_));
 sky130_fd_sc_hd__nand2_2 _15817_ (.A(_12850_),
    .B(_12856_),
    .Y(_12857_));
 sky130_fd_sc_hd__xor2_2 _15818_ (.A(_12855_),
    .B(_12857_),
    .X(_12858_));
 sky130_fd_sc_hd__a22o_2 _15819_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][10] ),
    .B1(_11712_),
    .B2(_12858_),
    .X(_01116_));
 sky130_fd_sc_hd__nor2_2 _15820_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[13][11] ),
    .Y(_12859_));
 sky130_fd_sc_hd__or2_2 _15821_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[13][11] ),
    .X(_12860_));
 sky130_fd_sc_hd__nand2_2 _15822_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[13][11] ),
    .Y(_12861_));
 sky130_fd_sc_hd__nand2_2 _15823_ (.A(_12860_),
    .B(_12861_),
    .Y(_12862_));
 sky130_fd_sc_hd__a21bo_2 _15824_ (.A1(_12855_),
    .A2(_12857_),
    .B1_N(_12853_),
    .X(_12863_));
 sky130_fd_sc_hd__xnor2_2 _15825_ (.A(_12862_),
    .B(_12863_),
    .Y(_12864_));
 sky130_fd_sc_hd__a22o_2 _15826_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][11] ),
    .B1(_11712_),
    .B2(_12864_),
    .X(_01117_));
 sky130_fd_sc_hd__nand3_2 _15827_ (.A(_12855_),
    .B(_12860_),
    .C(_12861_),
    .Y(_12865_));
 sky130_fd_sc_hd__nor2_2 _15828_ (.A(_12849_),
    .B(_12865_),
    .Y(_12866_));
 sky130_fd_sc_hd__o2bb2a_2 _15829_ (.A1_N(_12843_),
    .A2_N(_12866_),
    .B1(_12856_),
    .B2(_12865_),
    .X(_12867_));
 sky130_fd_sc_hd__o21a_2 _15830_ (.A1(_12853_),
    .A2(_12859_),
    .B1(_12861_),
    .X(_12868_));
 sky130_fd_sc_hd__xnor2_2 _15831_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[13][12] ),
    .Y(_12869_));
 sky130_fd_sc_hd__and3_2 _15832_ (.A(_12867_),
    .B(_12868_),
    .C(_12869_),
    .X(_12870_));
 sky130_fd_sc_hd__a21oi_2 _15833_ (.A1(_12867_),
    .A2(_12868_),
    .B1(_12869_),
    .Y(_12871_));
 sky130_fd_sc_hd__nor2_2 _15834_ (.A(_12870_),
    .B(_12871_),
    .Y(_12872_));
 sky130_fd_sc_hd__a22o_2 _15835_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][12] ),
    .B1(_11712_),
    .B2(_12872_),
    .X(_01118_));
 sky130_fd_sc_hd__xor2_2 _15836_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[13][13] ),
    .X(_12873_));
 sky130_fd_sc_hd__a211o_2 _15837_ (.A1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[13][12] ),
    .B1(_12871_),
    .C1(_12873_),
    .X(_12874_));
 sky130_fd_sc_hd__nand2b_2 _15838_ (.A_N(_12869_),
    .B(_12873_),
    .Y(_12875_));
 sky130_fd_sc_hd__a21o_2 _15839_ (.A1(_12867_),
    .A2(_12868_),
    .B1(_12875_),
    .X(_12876_));
 sky130_fd_sc_hd__and3_2 _15840_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[13][12] ),
    .C(_12873_),
    .X(_12877_));
 sky130_fd_sc_hd__nor2_2 _15841_ (.A(_11713_),
    .B(_12877_),
    .Y(_12878_));
 sky130_fd_sc_hd__a32o_2 _15842_ (.A1(_12874_),
    .A2(_12876_),
    .A3(_12878_),
    .B1(\systolic_inst.acc_wires[13][13] ),
    .B2(_11258_),
    .X(_01119_));
 sky130_fd_sc_hd__or2_2 _15843_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[13][14] ),
    .X(_12879_));
 sky130_fd_sc_hd__nand2_2 _15844_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[13][14] ),
    .Y(_12880_));
 sky130_fd_sc_hd__and2_2 _15845_ (.A(_12879_),
    .B(_12880_),
    .X(_12881_));
 sky130_fd_sc_hd__nand2_2 _15846_ (.A(_12879_),
    .B(_12880_),
    .Y(_12882_));
 sky130_fd_sc_hd__a21oi_2 _15847_ (.A1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[13][13] ),
    .B1(_12877_),
    .Y(_12883_));
 sky130_fd_sc_hd__nand2_2 _15848_ (.A(_12876_),
    .B(_12883_),
    .Y(_12884_));
 sky130_fd_sc_hd__nand2_2 _15849_ (.A(_12881_),
    .B(_12884_),
    .Y(_12885_));
 sky130_fd_sc_hd__or2_2 _15850_ (.A(_12881_),
    .B(_12884_),
    .X(_12886_));
 sky130_fd_sc_hd__a32o_2 _15851_ (.A1(_11712_),
    .A2(_12885_),
    .A3(_12886_),
    .B1(\systolic_inst.acc_wires[13][14] ),
    .B2(_11258_),
    .X(_01120_));
 sky130_fd_sc_hd__nor2_2 _15852_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][15] ),
    .Y(_12887_));
 sky130_fd_sc_hd__and2_2 _15853_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][15] ),
    .X(_12888_));
 sky130_fd_sc_hd__or2_2 _15854_ (.A(_12887_),
    .B(_12888_),
    .X(_12889_));
 sky130_fd_sc_hd__a21oi_2 _15855_ (.A1(_12880_),
    .A2(_12885_),
    .B1(_12889_),
    .Y(_12890_));
 sky130_fd_sc_hd__a31o_2 _15856_ (.A1(_12880_),
    .A2(_12885_),
    .A3(_12889_),
    .B1(_11713_),
    .X(_12891_));
 sky130_fd_sc_hd__a2bb2o_2 _15857_ (.A1_N(_12891_),
    .A2_N(_12890_),
    .B1(\systolic_inst.acc_wires[13][15] ),
    .B2(_11258_),
    .X(_01121_));
 sky130_fd_sc_hd__a211o_2 _15858_ (.A1(_12876_),
    .A2(_12883_),
    .B1(_12889_),
    .C1(_12882_),
    .X(_12892_));
 sky130_fd_sc_hd__o21ba_2 _15859_ (.A1(_12880_),
    .A2(_12887_),
    .B1_N(_12888_),
    .X(_12893_));
 sky130_fd_sc_hd__and2_2 _15860_ (.A(_12892_),
    .B(_12893_),
    .X(_12894_));
 sky130_fd_sc_hd__xnor2_2 _15861_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][16] ),
    .Y(_12895_));
 sky130_fd_sc_hd__nand2_2 _15862_ (.A(_12894_),
    .B(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__nor2_2 _15863_ (.A(_12894_),
    .B(_12895_),
    .Y(_12897_));
 sky130_fd_sc_hd__nor2_2 _15864_ (.A(_11713_),
    .B(_12897_),
    .Y(_12898_));
 sky130_fd_sc_hd__a22o_2 _15865_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][16] ),
    .B1(_12896_),
    .B2(_12898_),
    .X(_01122_));
 sky130_fd_sc_hd__xor2_2 _15866_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][17] ),
    .X(_12899_));
 sky130_fd_sc_hd__inv_2 _15867_ (.A(_12899_),
    .Y(_12900_));
 sky130_fd_sc_hd__a21oi_2 _15868_ (.A1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[13][16] ),
    .B1(_12897_),
    .Y(_12901_));
 sky130_fd_sc_hd__xnor2_2 _15869_ (.A(_12899_),
    .B(_12901_),
    .Y(_12902_));
 sky130_fd_sc_hd__a22o_2 _15870_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][17] ),
    .B1(_11712_),
    .B2(_12902_),
    .X(_01123_));
 sky130_fd_sc_hd__or2_2 _15871_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][18] ),
    .X(_12903_));
 sky130_fd_sc_hd__nand2_2 _15872_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][18] ),
    .Y(_12904_));
 sky130_fd_sc_hd__nand2_2 _15873_ (.A(_12903_),
    .B(_12904_),
    .Y(_12905_));
 sky130_fd_sc_hd__o21a_2 _15874_ (.A1(\systolic_inst.acc_wires[13][16] ),
    .A2(\systolic_inst.acc_wires[13][17] ),
    .B1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .X(_12906_));
 sky130_fd_sc_hd__a21oi_2 _15875_ (.A1(_12897_),
    .A2(_12899_),
    .B1(_12906_),
    .Y(_12907_));
 sky130_fd_sc_hd__xor2_2 _15876_ (.A(_12905_),
    .B(_12907_),
    .X(_12908_));
 sky130_fd_sc_hd__a22o_2 _15877_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][18] ),
    .B1(_11712_),
    .B2(_12908_),
    .X(_01124_));
 sky130_fd_sc_hd__xnor2_2 _15878_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][19] ),
    .Y(_12909_));
 sky130_fd_sc_hd__o21ai_2 _15879_ (.A1(_12905_),
    .A2(_12907_),
    .B1(_12904_),
    .Y(_12910_));
 sky130_fd_sc_hd__xnor2_2 _15880_ (.A(_12909_),
    .B(_12910_),
    .Y(_12911_));
 sky130_fd_sc_hd__a22o_2 _15881_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][19] ),
    .B1(_11712_),
    .B2(_12911_),
    .X(_01125_));
 sky130_fd_sc_hd__or2_2 _15882_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][20] ),
    .X(_12912_));
 sky130_fd_sc_hd__nand2_2 _15883_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][20] ),
    .Y(_12913_));
 sky130_fd_sc_hd__and2_2 _15884_ (.A(_12912_),
    .B(_12913_),
    .X(_12914_));
 sky130_fd_sc_hd__or4_2 _15885_ (.A(_12895_),
    .B(_12900_),
    .C(_12905_),
    .D(_12909_),
    .X(_12915_));
 sky130_fd_sc_hd__nor2_2 _15886_ (.A(_12894_),
    .B(_12915_),
    .Y(_12916_));
 sky130_fd_sc_hd__o41a_2 _15887_ (.A1(\systolic_inst.acc_wires[13][16] ),
    .A2(\systolic_inst.acc_wires[13][17] ),
    .A3(\systolic_inst.acc_wires[13][18] ),
    .A4(\systolic_inst.acc_wires[13][19] ),
    .B1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .X(_12917_));
 sky130_fd_sc_hd__or3_2 _15888_ (.A(_12914_),
    .B(_12916_),
    .C(_12917_),
    .X(_12918_));
 sky130_fd_sc_hd__o21ai_2 _15889_ (.A1(_12916_),
    .A2(_12917_),
    .B1(_12914_),
    .Y(_12919_));
 sky130_fd_sc_hd__a32o_2 _15890_ (.A1(_11712_),
    .A2(_12918_),
    .A3(_12919_),
    .B1(\systolic_inst.acc_wires[13][20] ),
    .B2(_11258_),
    .X(_01126_));
 sky130_fd_sc_hd__xnor2_2 _15891_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][21] ),
    .Y(_12920_));
 sky130_fd_sc_hd__inv_2 _15892_ (.A(_12920_),
    .Y(_12921_));
 sky130_fd_sc_hd__a21oi_2 _15893_ (.A1(_12913_),
    .A2(_12919_),
    .B1(_12920_),
    .Y(_12922_));
 sky130_fd_sc_hd__a31o_2 _15894_ (.A1(_12913_),
    .A2(_12919_),
    .A3(_12920_),
    .B1(_11713_),
    .X(_12923_));
 sky130_fd_sc_hd__a2bb2o_2 _15895_ (.A1_N(_12923_),
    .A2_N(_12922_),
    .B1(\systolic_inst.acc_wires[13][21] ),
    .B2(_11258_),
    .X(_01127_));
 sky130_fd_sc_hd__or2_2 _15896_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][22] ),
    .X(_12924_));
 sky130_fd_sc_hd__nand2_2 _15897_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][22] ),
    .Y(_12925_));
 sky130_fd_sc_hd__and2_2 _15898_ (.A(_12924_),
    .B(_12925_),
    .X(_12926_));
 sky130_fd_sc_hd__o21a_2 _15899_ (.A1(\systolic_inst.acc_wires[13][20] ),
    .A2(\systolic_inst.acc_wires[13][21] ),
    .B1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .X(_12927_));
 sky130_fd_sc_hd__nor2_2 _15900_ (.A(_12919_),
    .B(_12920_),
    .Y(_12928_));
 sky130_fd_sc_hd__o21ai_2 _15901_ (.A1(_12927_),
    .A2(_12928_),
    .B1(_12926_),
    .Y(_12929_));
 sky130_fd_sc_hd__or3_2 _15902_ (.A(_12926_),
    .B(_12927_),
    .C(_12928_),
    .X(_12930_));
 sky130_fd_sc_hd__a32o_2 _15903_ (.A1(_11712_),
    .A2(_12929_),
    .A3(_12930_),
    .B1(\systolic_inst.acc_wires[13][22] ),
    .B2(_11258_),
    .X(_01128_));
 sky130_fd_sc_hd__xor2_2 _15904_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][23] ),
    .X(_12931_));
 sky130_fd_sc_hd__inv_2 _15905_ (.A(_12931_),
    .Y(_12932_));
 sky130_fd_sc_hd__nand3_2 _15906_ (.A(_12925_),
    .B(_12929_),
    .C(_12932_),
    .Y(_12933_));
 sky130_fd_sc_hd__a21o_2 _15907_ (.A1(_12925_),
    .A2(_12929_),
    .B1(_12932_),
    .X(_12934_));
 sky130_fd_sc_hd__a32o_2 _15908_ (.A1(_11712_),
    .A2(_12933_),
    .A3(_12934_),
    .B1(\systolic_inst.acc_wires[13][23] ),
    .B2(_11258_),
    .X(_01129_));
 sky130_fd_sc_hd__nand4_2 _15909_ (.A(_12914_),
    .B(_12921_),
    .C(_12926_),
    .D(_12931_),
    .Y(_12935_));
 sky130_fd_sc_hd__a211o_2 _15910_ (.A1(_12892_),
    .A2(_12893_),
    .B1(_12915_),
    .C1(_12935_),
    .X(_12936_));
 sky130_fd_sc_hd__o41a_2 _15911_ (.A1(\systolic_inst.acc_wires[13][20] ),
    .A2(\systolic_inst.acc_wires[13][21] ),
    .A3(\systolic_inst.acc_wires[13][22] ),
    .A4(\systolic_inst.acc_wires[13][23] ),
    .B1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .X(_12937_));
 sky130_fd_sc_hd__nor2_2 _15912_ (.A(_12917_),
    .B(_12937_),
    .Y(_12938_));
 sky130_fd_sc_hd__nor2_2 _15913_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][24] ),
    .Y(_12939_));
 sky130_fd_sc_hd__and2_2 _15914_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][24] ),
    .X(_12940_));
 sky130_fd_sc_hd__or2_2 _15915_ (.A(_12939_),
    .B(_12940_),
    .X(_12941_));
 sky130_fd_sc_hd__a21oi_2 _15916_ (.A1(_12936_),
    .A2(_12938_),
    .B1(_12941_),
    .Y(_12942_));
 sky130_fd_sc_hd__a31o_2 _15917_ (.A1(_12936_),
    .A2(_12938_),
    .A3(_12941_),
    .B1(_11713_),
    .X(_12943_));
 sky130_fd_sc_hd__a2bb2o_2 _15918_ (.A1_N(_12943_),
    .A2_N(_12942_),
    .B1(\systolic_inst.acc_wires[13][24] ),
    .B2(_11258_),
    .X(_01130_));
 sky130_fd_sc_hd__xor2_2 _15919_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][25] ),
    .X(_12944_));
 sky130_fd_sc_hd__or3_2 _15920_ (.A(_12940_),
    .B(_12942_),
    .C(_12944_),
    .X(_12945_));
 sky130_fd_sc_hd__o21ai_2 _15921_ (.A1(_12940_),
    .A2(_12942_),
    .B1(_12944_),
    .Y(_12946_));
 sky130_fd_sc_hd__a32o_2 _15922_ (.A1(_11712_),
    .A2(_12945_),
    .A3(_12946_),
    .B1(\systolic_inst.acc_wires[13][25] ),
    .B2(_11258_),
    .X(_01131_));
 sky130_fd_sc_hd__or2_2 _15923_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][26] ),
    .X(_12947_));
 sky130_fd_sc_hd__nand2_2 _15924_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][26] ),
    .Y(_12948_));
 sky130_fd_sc_hd__nand2_2 _15925_ (.A(_12947_),
    .B(_12948_),
    .Y(_12949_));
 sky130_fd_sc_hd__o21a_2 _15926_ (.A1(\systolic_inst.acc_wires[13][24] ),
    .A2(\systolic_inst.acc_wires[13][25] ),
    .B1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .X(_12950_));
 sky130_fd_sc_hd__a21o_2 _15927_ (.A1(_12942_),
    .A2(_12944_),
    .B1(_12950_),
    .X(_12951_));
 sky130_fd_sc_hd__xnor2_2 _15928_ (.A(_12949_),
    .B(_12951_),
    .Y(_12952_));
 sky130_fd_sc_hd__a22o_2 _15929_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][26] ),
    .B1(_11712_),
    .B2(_12952_),
    .X(_01132_));
 sky130_fd_sc_hd__xnor2_2 _15930_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][27] ),
    .Y(_12953_));
 sky130_fd_sc_hd__a21bo_2 _15931_ (.A1(_12947_),
    .A2(_12951_),
    .B1_N(_12948_),
    .X(_12954_));
 sky130_fd_sc_hd__xnor2_2 _15932_ (.A(_12953_),
    .B(_12954_),
    .Y(_12955_));
 sky130_fd_sc_hd__a22o_2 _15933_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][27] ),
    .B1(_11712_),
    .B2(_12955_),
    .X(_01133_));
 sky130_fd_sc_hd__nor2_2 _15934_ (.A(_12949_),
    .B(_12953_),
    .Y(_12956_));
 sky130_fd_sc_hd__o21a_2 _15935_ (.A1(\systolic_inst.acc_wires[13][26] ),
    .A2(\systolic_inst.acc_wires[13][27] ),
    .B1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .X(_12957_));
 sky130_fd_sc_hd__a311oi_2 _15936_ (.A1(_12942_),
    .A2(_12944_),
    .A3(_12956_),
    .B1(_12957_),
    .C1(_12950_),
    .Y(_12958_));
 sky130_fd_sc_hd__or2_2 _15937_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][28] ),
    .X(_12959_));
 sky130_fd_sc_hd__nand2_2 _15938_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][28] ),
    .Y(_12960_));
 sky130_fd_sc_hd__nand2_2 _15939_ (.A(_12959_),
    .B(_12960_),
    .Y(_12961_));
 sky130_fd_sc_hd__xor2_2 _15940_ (.A(_12958_),
    .B(_12961_),
    .X(_12962_));
 sky130_fd_sc_hd__a22o_2 _15941_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][28] ),
    .B1(_11712_),
    .B2(_12962_),
    .X(_01134_));
 sky130_fd_sc_hd__xor2_2 _15942_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][29] ),
    .X(_12963_));
 sky130_fd_sc_hd__inv_2 _15943_ (.A(_12963_),
    .Y(_12964_));
 sky130_fd_sc_hd__o21a_2 _15944_ (.A1(_12958_),
    .A2(_12961_),
    .B1(_12960_),
    .X(_12965_));
 sky130_fd_sc_hd__xnor2_2 _15945_ (.A(_12963_),
    .B(_12965_),
    .Y(_12966_));
 sky130_fd_sc_hd__a22o_2 _15946_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[13][29] ),
    .B1(_11712_),
    .B2(_12966_),
    .X(_01135_));
 sky130_fd_sc_hd__o21ai_2 _15947_ (.A1(\systolic_inst.acc_wires[13][28] ),
    .A2(\systolic_inst.acc_wires[13][29] ),
    .B1(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .Y(_12967_));
 sky130_fd_sc_hd__o31a_2 _15948_ (.A1(_12958_),
    .A2(_12961_),
    .A3(_12964_),
    .B1(_12967_),
    .X(_12968_));
 sky130_fd_sc_hd__nand2_2 _15949_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][30] ),
    .Y(_12969_));
 sky130_fd_sc_hd__or2_2 _15950_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][30] ),
    .X(_12970_));
 sky130_fd_sc_hd__nand2_2 _15951_ (.A(_12969_),
    .B(_12970_),
    .Y(_12971_));
 sky130_fd_sc_hd__nand2_2 _15952_ (.A(_12968_),
    .B(_12971_),
    .Y(_12972_));
 sky130_fd_sc_hd__or2_2 _15953_ (.A(_12968_),
    .B(_12971_),
    .X(_12973_));
 sky130_fd_sc_hd__a32o_2 _15954_ (.A1(_11712_),
    .A2(_12972_),
    .A3(_12973_),
    .B1(\systolic_inst.acc_wires[13][30] ),
    .B2(_11258_),
    .X(_01136_));
 sky130_fd_sc_hd__xnor2_2 _15955_ (.A(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[13][31] ),
    .Y(_12974_));
 sky130_fd_sc_hd__a21oi_2 _15956_ (.A1(_12969_),
    .A2(_12973_),
    .B1(_12974_),
    .Y(_12975_));
 sky130_fd_sc_hd__a31o_2 _15957_ (.A1(_12969_),
    .A2(_12973_),
    .A3(_12974_),
    .B1(_11713_),
    .X(_12976_));
 sky130_fd_sc_hd__a2bb2o_2 _15958_ (.A1_N(_12976_),
    .A2_N(_12975_),
    .B1(\systolic_inst.acc_wires[13][31] ),
    .B2(_11258_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _15959_ (.A0(\systolic_inst.A_outs[12][0] ),
    .A1(\systolic_inst.A_shift[24][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _15960_ (.A0(\systolic_inst.A_outs[12][1] ),
    .A1(\systolic_inst.A_shift[24][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _15961_ (.A0(\systolic_inst.A_outs[12][2] ),
    .A1(\systolic_inst.A_shift[24][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _15962_ (.A0(\systolic_inst.A_outs[12][3] ),
    .A1(\systolic_inst.A_shift[24][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _15963_ (.A0(\systolic_inst.A_outs[12][4] ),
    .A1(\systolic_inst.A_shift[24][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _15964_ (.A0(\systolic_inst.A_outs[12][5] ),
    .A1(\systolic_inst.A_shift[24][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _15965_ (.A0(\systolic_inst.A_outs[12][6] ),
    .A1(\systolic_inst.A_shift[24][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _15966_ (.A0(\systolic_inst.A_outs[12][7] ),
    .A1(\systolic_inst.A_shift[24][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _15967_ (.A0(\systolic_inst.B_outs[11][0] ),
    .A1(\systolic_inst.B_outs[7][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _15968_ (.A0(\systolic_inst.B_outs[11][1] ),
    .A1(\systolic_inst.B_outs[7][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _15969_ (.A0(\systolic_inst.B_outs[11][2] ),
    .A1(\systolic_inst.B_outs[7][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _15970_ (.A0(\systolic_inst.B_outs[11][3] ),
    .A1(\systolic_inst.B_outs[7][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _15971_ (.A0(\systolic_inst.B_outs[11][4] ),
    .A1(\systolic_inst.B_outs[7][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _15972_ (.A0(\systolic_inst.B_outs[11][5] ),
    .A1(\systolic_inst.B_outs[7][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _15973_ (.A0(\systolic_inst.B_outs[11][6] ),
    .A1(\systolic_inst.B_outs[7][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _15974_ (.A0(\systolic_inst.B_outs[11][7] ),
    .A1(\systolic_inst.B_outs[7][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01153_));
 sky130_fd_sc_hd__and3_2 _15975_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[12][0] ),
    .C(\systolic_inst.A_outs[12][0] ),
    .X(_12977_));
 sky130_fd_sc_hd__a21o_2 _15976_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[0] ),
    .B1(_12977_),
    .X(_01154_));
 sky130_fd_sc_hd__and4_2 _15977_ (.A(\systolic_inst.B_outs[12][0] ),
    .B(\systolic_inst.A_outs[12][0] ),
    .C(\systolic_inst.B_outs[12][1] ),
    .D(\systolic_inst.A_outs[12][1] ),
    .X(_12978_));
 sky130_fd_sc_hd__a22o_2 _15978_ (.A1(\systolic_inst.A_outs[12][0] ),
    .A2(\systolic_inst.B_outs[12][1] ),
    .B1(\systolic_inst.A_outs[12][1] ),
    .B2(\systolic_inst.B_outs[12][0] ),
    .X(_12979_));
 sky130_fd_sc_hd__nand2_2 _15979_ (.A(\systolic_inst.ce_local ),
    .B(_12979_),
    .Y(_12980_));
 sky130_fd_sc_hd__a2bb2o_2 _15980_ (.A1_N(_12980_),
    .A2_N(_12978_),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01155_));
 sky130_fd_sc_hd__nand2_2 _15981_ (.A(\systolic_inst.B_outs[12][1] ),
    .B(\systolic_inst.A_outs[12][1] ),
    .Y(_12981_));
 sky130_fd_sc_hd__nand2_2 _15982_ (.A(\systolic_inst.B_outs[12][0] ),
    .B(\systolic_inst.A_outs[12][2] ),
    .Y(_12982_));
 sky130_fd_sc_hd__and4_2 _15983_ (.A(\systolic_inst.B_outs[12][0] ),
    .B(\systolic_inst.B_outs[12][1] ),
    .C(\systolic_inst.A_outs[12][1] ),
    .D(\systolic_inst.A_outs[12][2] ),
    .X(_12983_));
 sky130_fd_sc_hd__a21o_2 _15984_ (.A1(_12981_),
    .A2(_12982_),
    .B1(_12983_),
    .X(_12984_));
 sky130_fd_sc_hd__inv_2 _15985_ (.A(_12984_),
    .Y(_12985_));
 sky130_fd_sc_hd__xnor2_2 _15986_ (.A(_12978_),
    .B(_12984_),
    .Y(_12986_));
 sky130_fd_sc_hd__nand3_2 _15987_ (.A(\systolic_inst.A_outs[12][0] ),
    .B(\systolic_inst.B_outs[12][2] ),
    .C(_12986_),
    .Y(_12987_));
 sky130_fd_sc_hd__a21o_2 _15988_ (.A1(\systolic_inst.A_outs[12][0] ),
    .A2(\systolic_inst.B_outs[12][2] ),
    .B1(_12986_),
    .X(_12988_));
 sky130_fd_sc_hd__and2_2 _15989_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[2] ),
    .X(_12989_));
 sky130_fd_sc_hd__a31o_2 _15990_ (.A1(\systolic_inst.ce_local ),
    .A2(_12987_),
    .A3(_12988_),
    .B1(_12989_),
    .X(_01156_));
 sky130_fd_sc_hd__a22oi_2 _15991_ (.A1(\systolic_inst.A_outs[12][1] ),
    .A2(\systolic_inst.B_outs[12][2] ),
    .B1(\systolic_inst.B_outs[12][3] ),
    .B2(\systolic_inst.A_outs[12][0] ),
    .Y(_12990_));
 sky130_fd_sc_hd__and4_2 _15992_ (.A(\systolic_inst.A_outs[12][0] ),
    .B(\systolic_inst.A_outs[12][1] ),
    .C(\systolic_inst.B_outs[12][2] ),
    .D(\systolic_inst.B_outs[12][3] ),
    .X(_12991_));
 sky130_fd_sc_hd__or2_2 _15993_ (.A(_12990_),
    .B(_12991_),
    .X(_12992_));
 sky130_fd_sc_hd__nand2_2 _15994_ (.A(\systolic_inst.B_outs[12][1] ),
    .B(\systolic_inst.A_outs[12][3] ),
    .Y(_12993_));
 sky130_fd_sc_hd__or2_2 _15995_ (.A(_12982_),
    .B(_12993_),
    .X(_12994_));
 sky130_fd_sc_hd__a22o_2 _15996_ (.A1(\systolic_inst.B_outs[12][1] ),
    .A2(\systolic_inst.A_outs[12][2] ),
    .B1(\systolic_inst.A_outs[12][3] ),
    .B2(\systolic_inst.B_outs[12][0] ),
    .X(_12995_));
 sky130_fd_sc_hd__nand3_2 _15997_ (.A(_12983_),
    .B(_12994_),
    .C(_12995_),
    .Y(_12996_));
 sky130_fd_sc_hd__a21o_2 _15998_ (.A1(_12994_),
    .A2(_12995_),
    .B1(_12983_),
    .X(_12997_));
 sky130_fd_sc_hd__nand2_2 _15999_ (.A(_12996_),
    .B(_12997_),
    .Y(_12998_));
 sky130_fd_sc_hd__or2_2 _16000_ (.A(_12992_),
    .B(_12998_),
    .X(_12999_));
 sky130_fd_sc_hd__xnor2_2 _16001_ (.A(_12992_),
    .B(_12998_),
    .Y(_13000_));
 sky130_fd_sc_hd__a21bo_2 _16002_ (.A1(_12978_),
    .A2(_12985_),
    .B1_N(_12987_),
    .X(_13001_));
 sky130_fd_sc_hd__and2b_2 _16003_ (.A_N(_13000_),
    .B(_13001_),
    .X(_13002_));
 sky130_fd_sc_hd__xnor2_2 _16004_ (.A(_13000_),
    .B(_13001_),
    .Y(_13003_));
 sky130_fd_sc_hd__mux2_1 _16005_ (.A0(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[3] ),
    .A1(_13003_),
    .S(\systolic_inst.ce_local ),
    .X(_01157_));
 sky130_fd_sc_hd__and2_2 _16006_ (.A(\systolic_inst.B_outs[12][2] ),
    .B(\systolic_inst.A_outs[12][2] ),
    .X(_13004_));
 sky130_fd_sc_hd__nand4_2 _16007_ (.A(\systolic_inst.A_outs[12][0] ),
    .B(\systolic_inst.A_outs[12][1] ),
    .C(\systolic_inst.B_outs[12][3] ),
    .D(\systolic_inst.B_outs[12][4] ),
    .Y(_13005_));
 sky130_fd_sc_hd__a22o_2 _16008_ (.A1(\systolic_inst.A_outs[12][1] ),
    .A2(\systolic_inst.B_outs[12][3] ),
    .B1(\systolic_inst.B_outs[12][4] ),
    .B2(\systolic_inst.A_outs[12][0] ),
    .X(_13006_));
 sky130_fd_sc_hd__nand2_2 _16009_ (.A(_13005_),
    .B(_13006_),
    .Y(_13007_));
 sky130_fd_sc_hd__xnor2_2 _16010_ (.A(_13004_),
    .B(_13007_),
    .Y(_13008_));
 sky130_fd_sc_hd__inv_2 _16011_ (.A(_13008_),
    .Y(_13009_));
 sky130_fd_sc_hd__nand2_2 _16012_ (.A(\systolic_inst.B_outs[12][0] ),
    .B(\systolic_inst.A_outs[12][4] ),
    .Y(_13010_));
 sky130_fd_sc_hd__and4_2 _16013_ (.A(\systolic_inst.B_outs[12][0] ),
    .B(\systolic_inst.B_outs[12][1] ),
    .C(\systolic_inst.A_outs[12][3] ),
    .D(\systolic_inst.A_outs[12][4] ),
    .X(_13011_));
 sky130_fd_sc_hd__a21oi_2 _16014_ (.A1(_12993_),
    .A2(_13010_),
    .B1(_13011_),
    .Y(_13012_));
 sky130_fd_sc_hd__xnor2_2 _16015_ (.A(_12991_),
    .B(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__nor2_2 _16016_ (.A(_12994_),
    .B(_13013_),
    .Y(_13014_));
 sky130_fd_sc_hd__xnor2_2 _16017_ (.A(_12994_),
    .B(_13013_),
    .Y(_13015_));
 sky130_fd_sc_hd__nor2_2 _16018_ (.A(_13009_),
    .B(_13015_),
    .Y(_13016_));
 sky130_fd_sc_hd__and2_2 _16019_ (.A(_13009_),
    .B(_13015_),
    .X(_13017_));
 sky130_fd_sc_hd__or2_2 _16020_ (.A(_13016_),
    .B(_13017_),
    .X(_13018_));
 sky130_fd_sc_hd__a21o_2 _16021_ (.A1(_12996_),
    .A2(_12999_),
    .B1(_13018_),
    .X(_13019_));
 sky130_fd_sc_hd__inv_2 _16022_ (.A(_13019_),
    .Y(_13020_));
 sky130_fd_sc_hd__nand3_2 _16023_ (.A(_12996_),
    .B(_12999_),
    .C(_13018_),
    .Y(_13021_));
 sky130_fd_sc_hd__a21oi_2 _16024_ (.A1(_13019_),
    .A2(_13021_),
    .B1(_13002_),
    .Y(_13022_));
 sky130_fd_sc_hd__and3_2 _16025_ (.A(_13002_),
    .B(_13019_),
    .C(_13021_),
    .X(_13023_));
 sky130_fd_sc_hd__or3_2 _16026_ (.A(_11258_),
    .B(_13022_),
    .C(_13023_),
    .X(_13024_));
 sky130_fd_sc_hd__a21bo_2 _16027_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[4] ),
    .B1_N(_13024_),
    .X(_01158_));
 sky130_fd_sc_hd__and2_2 _16028_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[5] ),
    .X(_13025_));
 sky130_fd_sc_hd__a21oi_2 _16029_ (.A1(_12991_),
    .A2(_13012_),
    .B1(_13014_),
    .Y(_13026_));
 sky130_fd_sc_hd__a21bo_2 _16030_ (.A1(_13004_),
    .A2(_13006_),
    .B1_N(_13005_),
    .X(_13027_));
 sky130_fd_sc_hd__a22oi_2 _16031_ (.A1(\systolic_inst.B_outs[12][1] ),
    .A2(\systolic_inst.A_outs[12][4] ),
    .B1(\systolic_inst.A_outs[12][5] ),
    .B2(\systolic_inst.B_outs[12][0] ),
    .Y(_13028_));
 sky130_fd_sc_hd__and4_2 _16032_ (.A(\systolic_inst.B_outs[12][0] ),
    .B(\systolic_inst.B_outs[12][1] ),
    .C(\systolic_inst.A_outs[12][4] ),
    .D(\systolic_inst.A_outs[12][5] ),
    .X(_13029_));
 sky130_fd_sc_hd__or2_2 _16033_ (.A(_13028_),
    .B(_13029_),
    .X(_13030_));
 sky130_fd_sc_hd__nand2b_2 _16034_ (.A_N(_13030_),
    .B(_13027_),
    .Y(_13031_));
 sky130_fd_sc_hd__xnor2_2 _16035_ (.A(_13027_),
    .B(_13030_),
    .Y(_13032_));
 sky130_fd_sc_hd__nand2_2 _16036_ (.A(_13011_),
    .B(_13032_),
    .Y(_13033_));
 sky130_fd_sc_hd__xnor2_2 _16037_ (.A(_13011_),
    .B(_13032_),
    .Y(_13034_));
 sky130_fd_sc_hd__nand2_2 _16038_ (.A(\systolic_inst.A_outs[12][0] ),
    .B(\systolic_inst.B_outs[12][5] ),
    .Y(_13035_));
 sky130_fd_sc_hd__nand2_2 _16039_ (.A(\systolic_inst.B_outs[12][2] ),
    .B(\systolic_inst.A_outs[12][3] ),
    .Y(_13036_));
 sky130_fd_sc_hd__and4_2 _16040_ (.A(\systolic_inst.A_outs[12][1] ),
    .B(\systolic_inst.A_outs[12][2] ),
    .C(\systolic_inst.B_outs[12][3] ),
    .D(\systolic_inst.B_outs[12][4] ),
    .X(_13037_));
 sky130_fd_sc_hd__a22o_2 _16041_ (.A1(\systolic_inst.A_outs[12][2] ),
    .A2(\systolic_inst.B_outs[12][3] ),
    .B1(\systolic_inst.B_outs[12][4] ),
    .B2(\systolic_inst.A_outs[12][1] ),
    .X(_13038_));
 sky130_fd_sc_hd__and2b_2 _16042_ (.A_N(_13037_),
    .B(_13038_),
    .X(_13039_));
 sky130_fd_sc_hd__xnor2_2 _16043_ (.A(_13036_),
    .B(_13039_),
    .Y(_13040_));
 sky130_fd_sc_hd__nand2b_2 _16044_ (.A_N(_13035_),
    .B(_13040_),
    .Y(_13041_));
 sky130_fd_sc_hd__xor2_2 _16045_ (.A(_13035_),
    .B(_13040_),
    .X(_13042_));
 sky130_fd_sc_hd__nor2_2 _16046_ (.A(_13034_),
    .B(_13042_),
    .Y(_13043_));
 sky130_fd_sc_hd__inv_2 _16047_ (.A(_13043_),
    .Y(_13044_));
 sky130_fd_sc_hd__and2_2 _16048_ (.A(_13034_),
    .B(_13042_),
    .X(_13045_));
 sky130_fd_sc_hd__nor2_2 _16049_ (.A(_13043_),
    .B(_13045_),
    .Y(_13046_));
 sky130_fd_sc_hd__nand2_2 _16050_ (.A(_13016_),
    .B(_13046_),
    .Y(_13047_));
 sky130_fd_sc_hd__or2_2 _16051_ (.A(_13016_),
    .B(_13046_),
    .X(_13048_));
 sky130_fd_sc_hd__and2_2 _16052_ (.A(_13047_),
    .B(_13048_),
    .X(_13049_));
 sky130_fd_sc_hd__nand2b_2 _16053_ (.A_N(_13026_),
    .B(_13049_),
    .Y(_13050_));
 sky130_fd_sc_hd__xnor2_2 _16054_ (.A(_13026_),
    .B(_13049_),
    .Y(_13051_));
 sky130_fd_sc_hd__nor2_2 _16055_ (.A(_13020_),
    .B(_13023_),
    .Y(_13052_));
 sky130_fd_sc_hd__or3_2 _16056_ (.A(_13020_),
    .B(_13023_),
    .C(_13051_),
    .X(_13053_));
 sky130_fd_sc_hd__nand2b_2 _16057_ (.A_N(_13052_),
    .B(_13051_),
    .Y(_13054_));
 sky130_fd_sc_hd__a31o_2 _16058_ (.A1(\systolic_inst.ce_local ),
    .A2(_13053_),
    .A3(_13054_),
    .B1(_13025_),
    .X(_01159_));
 sky130_fd_sc_hd__a31o_2 _16059_ (.A1(\systolic_inst.B_outs[12][2] ),
    .A2(\systolic_inst.A_outs[12][3] ),
    .A3(_13038_),
    .B1(_13037_),
    .X(_13055_));
 sky130_fd_sc_hd__a22oi_2 _16060_ (.A1(\systolic_inst.B_outs[12][1] ),
    .A2(\systolic_inst.A_outs[12][5] ),
    .B1(\systolic_inst.A_outs[12][6] ),
    .B2(\systolic_inst.B_outs[12][0] ),
    .Y(_13056_));
 sky130_fd_sc_hd__and4_2 _16061_ (.A(\systolic_inst.B_outs[12][0] ),
    .B(\systolic_inst.B_outs[12][1] ),
    .C(\systolic_inst.A_outs[12][5] ),
    .D(\systolic_inst.A_outs[12][6] ),
    .X(_13057_));
 sky130_fd_sc_hd__nor2_2 _16062_ (.A(_13056_),
    .B(_13057_),
    .Y(_13058_));
 sky130_fd_sc_hd__xor2_2 _16063_ (.A(_13055_),
    .B(_13058_),
    .X(_13059_));
 sky130_fd_sc_hd__and2_2 _16064_ (.A(_13029_),
    .B(_13059_),
    .X(_13060_));
 sky130_fd_sc_hd__nor2_2 _16065_ (.A(_13029_),
    .B(_13059_),
    .Y(_13061_));
 sky130_fd_sc_hd__or2_2 _16066_ (.A(_13060_),
    .B(_13061_),
    .X(_13062_));
 sky130_fd_sc_hd__nand2_2 _16067_ (.A(\systolic_inst.B_outs[12][2] ),
    .B(\systolic_inst.A_outs[12][4] ),
    .Y(_13063_));
 sky130_fd_sc_hd__and4_2 _16068_ (.A(\systolic_inst.A_outs[12][2] ),
    .B(\systolic_inst.B_outs[12][3] ),
    .C(\systolic_inst.A_outs[12][3] ),
    .D(\systolic_inst.B_outs[12][4] ),
    .X(_13064_));
 sky130_fd_sc_hd__a22oi_2 _16069_ (.A1(\systolic_inst.B_outs[12][3] ),
    .A2(\systolic_inst.A_outs[12][3] ),
    .B1(\systolic_inst.B_outs[12][4] ),
    .B2(\systolic_inst.A_outs[12][2] ),
    .Y(_13065_));
 sky130_fd_sc_hd__or2_2 _16070_ (.A(_13064_),
    .B(_13065_),
    .X(_13066_));
 sky130_fd_sc_hd__xnor2_2 _16071_ (.A(_13063_),
    .B(_13066_),
    .Y(_13067_));
 sky130_fd_sc_hd__a22oi_2 _16072_ (.A1(\systolic_inst.A_outs[12][1] ),
    .A2(\systolic_inst.B_outs[12][5] ),
    .B1(\systolic_inst.B_outs[12][6] ),
    .B2(\systolic_inst.A_outs[12][0] ),
    .Y(_13068_));
 sky130_fd_sc_hd__nand2_2 _16073_ (.A(\systolic_inst.A_outs[12][1] ),
    .B(\systolic_inst.B_outs[12][6] ),
    .Y(_13069_));
 sky130_fd_sc_hd__nor2_2 _16074_ (.A(_13035_),
    .B(_13069_),
    .Y(_13070_));
 sky130_fd_sc_hd__nor2_2 _16075_ (.A(_13068_),
    .B(_13070_),
    .Y(_13071_));
 sky130_fd_sc_hd__or3_2 _16076_ (.A(_13067_),
    .B(_13068_),
    .C(_13070_),
    .X(_13072_));
 sky130_fd_sc_hd__xor2_2 _16077_ (.A(_13067_),
    .B(_13071_),
    .X(_13073_));
 sky130_fd_sc_hd__xnor2_2 _16078_ (.A(_13041_),
    .B(_13073_),
    .Y(_13074_));
 sky130_fd_sc_hd__xnor2_2 _16079_ (.A(_13062_),
    .B(_13074_),
    .Y(_13075_));
 sky130_fd_sc_hd__xnor2_2 _16080_ (.A(_13044_),
    .B(_13075_),
    .Y(_13076_));
 sky130_fd_sc_hd__a21oi_2 _16081_ (.A1(_13031_),
    .A2(_13033_),
    .B1(_13076_),
    .Y(_13077_));
 sky130_fd_sc_hd__and3_2 _16082_ (.A(_13031_),
    .B(_13033_),
    .C(_13076_),
    .X(_13078_));
 sky130_fd_sc_hd__a211oi_2 _16083_ (.A1(_13047_),
    .A2(_13050_),
    .B1(_13077_),
    .C1(_13078_),
    .Y(_13079_));
 sky130_fd_sc_hd__o211a_2 _16084_ (.A1(_13077_),
    .A2(_13078_),
    .B1(_13047_),
    .C1(_13050_),
    .X(_13080_));
 sky130_fd_sc_hd__o21ai_2 _16085_ (.A1(_13079_),
    .A2(_13080_),
    .B1(_13054_),
    .Y(_13081_));
 sky130_fd_sc_hd__nor3_2 _16086_ (.A(_13054_),
    .B(_13079_),
    .C(_13080_),
    .Y(_13082_));
 sky130_fd_sc_hd__nor2_2 _16087_ (.A(_11258_),
    .B(_13082_),
    .Y(_13083_));
 sky130_fd_sc_hd__a22o_2 _16088_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[6] ),
    .B1(_13081_),
    .B2(_13083_),
    .X(_01160_));
 sky130_fd_sc_hd__o21ba_2 _16089_ (.A1(_13044_),
    .A2(_13075_),
    .B1_N(_13077_),
    .X(_13084_));
 sky130_fd_sc_hd__a21oi_2 _16090_ (.A1(_13055_),
    .A2(_13058_),
    .B1(_13060_),
    .Y(_13085_));
 sky130_fd_sc_hd__o21ba_2 _16091_ (.A1(_13063_),
    .A2(_13065_),
    .B1_N(_13064_),
    .X(_13086_));
 sky130_fd_sc_hd__a22o_2 _16092_ (.A1(\systolic_inst.B_outs[12][1] ),
    .A2(\systolic_inst.A_outs[12][6] ),
    .B1(\systolic_inst.A_outs[12][7] ),
    .B2(\systolic_inst.B_outs[12][0] ),
    .X(_13087_));
 sky130_fd_sc_hd__nand4_2 _16093_ (.A(\systolic_inst.B_outs[12][0] ),
    .B(\systolic_inst.B_outs[12][1] ),
    .C(\systolic_inst.A_outs[12][6] ),
    .D(\systolic_inst.A_outs[12][7] ),
    .Y(_13088_));
 sky130_fd_sc_hd__nand2_2 _16094_ (.A(_13087_),
    .B(_13088_),
    .Y(_13089_));
 sky130_fd_sc_hd__xnor2_2 _16095_ (.A(_11260_),
    .B(_13089_),
    .Y(_13090_));
 sky130_fd_sc_hd__nor2_2 _16096_ (.A(_13086_),
    .B(_13090_),
    .Y(_13091_));
 sky130_fd_sc_hd__and2_2 _16097_ (.A(_13086_),
    .B(_13090_),
    .X(_13092_));
 sky130_fd_sc_hd__nor2_2 _16098_ (.A(_13091_),
    .B(_13092_),
    .Y(_13093_));
 sky130_fd_sc_hd__xnor2_2 _16099_ (.A(_13057_),
    .B(_13093_),
    .Y(_13094_));
 sky130_fd_sc_hd__nand2_2 _16100_ (.A(\systolic_inst.B_outs[12][2] ),
    .B(\systolic_inst.A_outs[12][5] ),
    .Y(_13095_));
 sky130_fd_sc_hd__and4_2 _16101_ (.A(\systolic_inst.B_outs[12][3] ),
    .B(\systolic_inst.A_outs[12][3] ),
    .C(\systolic_inst.B_outs[12][4] ),
    .D(\systolic_inst.A_outs[12][4] ),
    .X(_13096_));
 sky130_fd_sc_hd__a22oi_2 _16102_ (.A1(\systolic_inst.A_outs[12][3] ),
    .A2(\systolic_inst.B_outs[12][4] ),
    .B1(\systolic_inst.A_outs[12][4] ),
    .B2(\systolic_inst.B_outs[12][3] ),
    .Y(_13097_));
 sky130_fd_sc_hd__or2_2 _16103_ (.A(_13096_),
    .B(_13097_),
    .X(_13098_));
 sky130_fd_sc_hd__xnor2_2 _16104_ (.A(_13095_),
    .B(_13098_),
    .Y(_13099_));
 sky130_fd_sc_hd__nand2_2 _16105_ (.A(\systolic_inst.A_outs[12][2] ),
    .B(\systolic_inst.B_outs[12][5] ),
    .Y(_13100_));
 sky130_fd_sc_hd__and2b_2 _16106_ (.A_N(\systolic_inst.A_outs[12][0] ),
    .B(\systolic_inst.B_outs[12][7] ),
    .X(_03492_));
 sky130_fd_sc_hd__and3_2 _16107_ (.A(\systolic_inst.A_outs[12][1] ),
    .B(\systolic_inst.B_outs[12][6] ),
    .C(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__xnor2_2 _16108_ (.A(_13069_),
    .B(_03492_),
    .Y(_03494_));
 sky130_fd_sc_hd__xnor2_2 _16109_ (.A(_13100_),
    .B(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__xnor2_2 _16110_ (.A(_13070_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__nor2_2 _16111_ (.A(_13099_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__xnor2_2 _16112_ (.A(_13099_),
    .B(_03496_),
    .Y(_03498_));
 sky130_fd_sc_hd__or2_2 _16113_ (.A(_13072_),
    .B(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__and2_2 _16114_ (.A(_13072_),
    .B(_03498_),
    .X(_03500_));
 sky130_fd_sc_hd__xor2_2 _16115_ (.A(_13072_),
    .B(_03498_),
    .X(_03501_));
 sky130_fd_sc_hd__xnor2_2 _16116_ (.A(_13094_),
    .B(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__o32a_2 _16117_ (.A1(_13060_),
    .A2(_13061_),
    .A3(_13074_),
    .B1(_13073_),
    .B2(_13041_),
    .X(_03503_));
 sky130_fd_sc_hd__nand2b_2 _16118_ (.A_N(_03503_),
    .B(_03502_),
    .Y(_03504_));
 sky130_fd_sc_hd__xnor2_2 _16119_ (.A(_03502_),
    .B(_03503_),
    .Y(_03505_));
 sky130_fd_sc_hd__nand2b_2 _16120_ (.A_N(_13085_),
    .B(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__xnor2_2 _16121_ (.A(_13085_),
    .B(_03505_),
    .Y(_03507_));
 sky130_fd_sc_hd__and2b_2 _16122_ (.A_N(_13084_),
    .B(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__xnor2_2 _16123_ (.A(_13084_),
    .B(_03507_),
    .Y(_03509_));
 sky130_fd_sc_hd__nor3_2 _16124_ (.A(_13079_),
    .B(_13082_),
    .C(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__o21a_2 _16125_ (.A1(_13079_),
    .A2(_13082_),
    .B1(_03509_),
    .X(_03511_));
 sky130_fd_sc_hd__nand2_2 _16126_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[7] ),
    .Y(_03512_));
 sky130_fd_sc_hd__o31ai_2 _16127_ (.A1(_11258_),
    .A2(_03510_),
    .A3(_03511_),
    .B1(_03512_),
    .Y(_01161_));
 sky130_fd_sc_hd__a21o_2 _16128_ (.A1(_13057_),
    .A2(_13093_),
    .B1(_13091_),
    .X(_03513_));
 sky130_fd_sc_hd__a21bo_2 _16129_ (.A1(\systolic_inst.B_outs[12][7] ),
    .A2(_13087_),
    .B1_N(_13088_),
    .X(_03514_));
 sky130_fd_sc_hd__o21bai_2 _16130_ (.A1(_13095_),
    .A2(_13097_),
    .B1_N(_13096_),
    .Y(_03515_));
 sky130_fd_sc_hd__o21a_2 _16131_ (.A1(\systolic_inst.B_outs[12][0] ),
    .A2(\systolic_inst.B_outs[12][1] ),
    .B1(\systolic_inst.A_outs[12][7] ),
    .X(_03516_));
 sky130_fd_sc_hd__o21ai_2 _16132_ (.A1(\systolic_inst.B_outs[12][0] ),
    .A2(\systolic_inst.B_outs[12][1] ),
    .B1(\systolic_inst.A_outs[12][7] ),
    .Y(_03517_));
 sky130_fd_sc_hd__a21o_2 _16133_ (.A1(\systolic_inst.B_outs[12][0] ),
    .A2(\systolic_inst.B_outs[12][1] ),
    .B1(_03517_),
    .X(_03518_));
 sky130_fd_sc_hd__and2b_2 _16134_ (.A_N(_03518_),
    .B(_03515_),
    .X(_03519_));
 sky130_fd_sc_hd__xnor2_2 _16135_ (.A(_03515_),
    .B(_03518_),
    .Y(_03520_));
 sky130_fd_sc_hd__xnor2_2 _16136_ (.A(_03514_),
    .B(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__and4_2 _16137_ (.A(\systolic_inst.B_outs[12][3] ),
    .B(\systolic_inst.B_outs[12][4] ),
    .C(\systolic_inst.A_outs[12][4] ),
    .D(\systolic_inst.A_outs[12][5] ),
    .X(_03522_));
 sky130_fd_sc_hd__a22oi_2 _16138_ (.A1(\systolic_inst.B_outs[12][4] ),
    .A2(\systolic_inst.A_outs[12][4] ),
    .B1(\systolic_inst.A_outs[12][5] ),
    .B2(\systolic_inst.B_outs[12][3] ),
    .Y(_03523_));
 sky130_fd_sc_hd__nor2_2 _16139_ (.A(_03522_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__nand2_2 _16140_ (.A(\systolic_inst.B_outs[12][2] ),
    .B(\systolic_inst.A_outs[12][6] ),
    .Y(_03525_));
 sky130_fd_sc_hd__xnor2_2 _16141_ (.A(_03524_),
    .B(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2_2 _16142_ (.A(\systolic_inst.A_outs[12][3] ),
    .B(\systolic_inst.B_outs[12][5] ),
    .Y(_03527_));
 sky130_fd_sc_hd__and4b_2 _16143_ (.A_N(\systolic_inst.A_outs[12][1] ),
    .B(\systolic_inst.A_outs[12][2] ),
    .C(\systolic_inst.B_outs[12][6] ),
    .D(\systolic_inst.B_outs[12][7] ),
    .X(_03528_));
 sky130_fd_sc_hd__o2bb2a_2 _16144_ (.A1_N(\systolic_inst.A_outs[12][2] ),
    .A2_N(\systolic_inst.B_outs[12][6] ),
    .B1(_11260_),
    .B2(\systolic_inst.A_outs[12][1] ),
    .X(_03529_));
 sky130_fd_sc_hd__nor2_2 _16145_ (.A(_03528_),
    .B(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__xnor2_2 _16146_ (.A(_03527_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__a31oi_2 _16147_ (.A1(\systolic_inst.A_outs[12][2] ),
    .A2(\systolic_inst.B_outs[12][5] ),
    .A3(_03494_),
    .B1(_03493_),
    .Y(_03532_));
 sky130_fd_sc_hd__nand2b_2 _16148_ (.A_N(_03532_),
    .B(_03531_),
    .Y(_03533_));
 sky130_fd_sc_hd__xnor2_2 _16149_ (.A(_03531_),
    .B(_03532_),
    .Y(_03534_));
 sky130_fd_sc_hd__nand2_2 _16150_ (.A(_03526_),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__xnor2_2 _16151_ (.A(_03526_),
    .B(_03534_),
    .Y(_03536_));
 sky130_fd_sc_hd__a21oi_2 _16152_ (.A1(_13070_),
    .A2(_03495_),
    .B1(_03497_),
    .Y(_03537_));
 sky130_fd_sc_hd__xnor2_2 _16153_ (.A(_03536_),
    .B(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__or2_2 _16154_ (.A(_03521_),
    .B(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__xor2_2 _16155_ (.A(_03521_),
    .B(_03538_),
    .X(_03540_));
 sky130_fd_sc_hd__o21a_2 _16156_ (.A1(_13094_),
    .A2(_03500_),
    .B1(_03499_),
    .X(_03541_));
 sky130_fd_sc_hd__nand2b_2 _16157_ (.A_N(_03541_),
    .B(_03540_),
    .Y(_03542_));
 sky130_fd_sc_hd__xor2_2 _16158_ (.A(_03540_),
    .B(_03541_),
    .X(_03543_));
 sky130_fd_sc_hd__nand2b_2 _16159_ (.A_N(_03543_),
    .B(_03513_),
    .Y(_03544_));
 sky130_fd_sc_hd__xor2_2 _16160_ (.A(_03513_),
    .B(_03543_),
    .X(_03545_));
 sky130_fd_sc_hd__and2_2 _16161_ (.A(_03504_),
    .B(_03506_),
    .X(_03546_));
 sky130_fd_sc_hd__nor2_2 _16162_ (.A(_03545_),
    .B(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__inv_2 _16163_ (.A(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__and2_2 _16164_ (.A(_03545_),
    .B(_03546_),
    .X(_03549_));
 sky130_fd_sc_hd__nor2_2 _16165_ (.A(_03547_),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__o21a_2 _16166_ (.A1(_03508_),
    .A2(_03511_),
    .B1(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__o21ai_2 _16167_ (.A1(_03508_),
    .A2(_03511_),
    .B1(_03550_),
    .Y(_03552_));
 sky130_fd_sc_hd__or3_2 _16168_ (.A(_03508_),
    .B(_03511_),
    .C(_03550_),
    .X(_03553_));
 sky130_fd_sc_hd__and2_2 _16169_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[8] ),
    .X(_03554_));
 sky130_fd_sc_hd__a31o_2 _16170_ (.A1(\systolic_inst.ce_local ),
    .A2(_03552_),
    .A3(_03553_),
    .B1(_03554_),
    .X(_01162_));
 sky130_fd_sc_hd__a21o_2 _16171_ (.A1(_03514_),
    .A2(_03520_),
    .B1(_03519_),
    .X(_03555_));
 sky130_fd_sc_hd__o21ba_2 _16172_ (.A1(_03523_),
    .A2(_03525_),
    .B1_N(_03522_),
    .X(_03556_));
 sky130_fd_sc_hd__nor2_2 _16173_ (.A(_03517_),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__and2_2 _16174_ (.A(_03517_),
    .B(_03556_),
    .X(_03558_));
 sky130_fd_sc_hd__or2_2 _16175_ (.A(_03557_),
    .B(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__nand2_2 _16176_ (.A(\systolic_inst.B_outs[12][2] ),
    .B(\systolic_inst.A_outs[12][7] ),
    .Y(_03560_));
 sky130_fd_sc_hd__a22oi_2 _16177_ (.A1(\systolic_inst.B_outs[12][4] ),
    .A2(\systolic_inst.A_outs[12][5] ),
    .B1(\systolic_inst.A_outs[12][6] ),
    .B2(\systolic_inst.B_outs[12][3] ),
    .Y(_03561_));
 sky130_fd_sc_hd__and4_2 _16178_ (.A(\systolic_inst.B_outs[12][3] ),
    .B(\systolic_inst.B_outs[12][4] ),
    .C(\systolic_inst.A_outs[12][5] ),
    .D(\systolic_inst.A_outs[12][6] ),
    .X(_03562_));
 sky130_fd_sc_hd__nor2_2 _16179_ (.A(_03561_),
    .B(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__xnor2_2 _16180_ (.A(_03560_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand2_2 _16181_ (.A(\systolic_inst.A_outs[12][4] ),
    .B(\systolic_inst.B_outs[12][5] ),
    .Y(_03565_));
 sky130_fd_sc_hd__and4b_2 _16182_ (.A_N(\systolic_inst.A_outs[12][2] ),
    .B(\systolic_inst.A_outs[12][3] ),
    .C(\systolic_inst.B_outs[12][6] ),
    .D(\systolic_inst.B_outs[12][7] ),
    .X(_03566_));
 sky130_fd_sc_hd__o2bb2a_2 _16183_ (.A1_N(\systolic_inst.A_outs[12][3] ),
    .A2_N(\systolic_inst.B_outs[12][6] ),
    .B1(_11260_),
    .B2(\systolic_inst.A_outs[12][2] ),
    .X(_03567_));
 sky130_fd_sc_hd__nor2_2 _16184_ (.A(_03566_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__xnor2_2 _16185_ (.A(_03565_),
    .B(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__o21ba_2 _16186_ (.A1(_03527_),
    .A2(_03529_),
    .B1_N(_03528_),
    .X(_03570_));
 sky130_fd_sc_hd__nand2b_2 _16187_ (.A_N(_03570_),
    .B(_03569_),
    .Y(_03571_));
 sky130_fd_sc_hd__xnor2_2 _16188_ (.A(_03569_),
    .B(_03570_),
    .Y(_03572_));
 sky130_fd_sc_hd__xnor2_2 _16189_ (.A(_03564_),
    .B(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__a21o_2 _16190_ (.A1(_03533_),
    .A2(_03535_),
    .B1(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__nand3_2 _16191_ (.A(_03533_),
    .B(_03535_),
    .C(_03573_),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2_2 _16192_ (.A(_03574_),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__xor2_2 _16193_ (.A(_03559_),
    .B(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__o21a_2 _16194_ (.A1(_03536_),
    .A2(_03537_),
    .B1(_03539_),
    .X(_03578_));
 sky130_fd_sc_hd__nand2b_2 _16195_ (.A_N(_03578_),
    .B(_03577_),
    .Y(_03579_));
 sky130_fd_sc_hd__xnor2_2 _16196_ (.A(_03577_),
    .B(_03578_),
    .Y(_03580_));
 sky130_fd_sc_hd__xnor2_2 _16197_ (.A(_03555_),
    .B(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__a21oi_2 _16198_ (.A1(_03542_),
    .A2(_03544_),
    .B1(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__inv_2 _16199_ (.A(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__and3_2 _16200_ (.A(_03542_),
    .B(_03544_),
    .C(_03581_),
    .X(_03584_));
 sky130_fd_sc_hd__nor2_2 _16201_ (.A(_03582_),
    .B(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__o21ai_2 _16202_ (.A1(_03547_),
    .A2(_03551_),
    .B1(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__or3_2 _16203_ (.A(_03547_),
    .B(_03551_),
    .C(_03585_),
    .X(_03587_));
 sky130_fd_sc_hd__and2_2 _16204_ (.A(_11258_),
    .B(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[9] ),
    .X(_03588_));
 sky130_fd_sc_hd__a31o_2 _16205_ (.A1(\systolic_inst.ce_local ),
    .A2(_03586_),
    .A3(_03587_),
    .B1(_03588_),
    .X(_01163_));
 sky130_fd_sc_hd__o21ba_2 _16206_ (.A1(_03560_),
    .A2(_03561_),
    .B1_N(_03562_),
    .X(_03589_));
 sky130_fd_sc_hd__nor2_2 _16207_ (.A(_03517_),
    .B(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__and2_2 _16208_ (.A(_03517_),
    .B(_03589_),
    .X(_03591_));
 sky130_fd_sc_hd__or2_2 _16209_ (.A(_03590_),
    .B(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__a22o_2 _16210_ (.A1(\systolic_inst.B_outs[12][4] ),
    .A2(\systolic_inst.A_outs[12][6] ),
    .B1(\systolic_inst.A_outs[12][7] ),
    .B2(\systolic_inst.B_outs[12][3] ),
    .X(_03593_));
 sky130_fd_sc_hd__and3_2 _16211_ (.A(\systolic_inst.B_outs[12][3] ),
    .B(\systolic_inst.B_outs[12][4] ),
    .C(\systolic_inst.A_outs[12][7] ),
    .X(_03594_));
 sky130_fd_sc_hd__a21bo_2 _16212_ (.A1(\systolic_inst.A_outs[12][6] ),
    .A2(_03594_),
    .B1_N(_03593_),
    .X(_03595_));
 sky130_fd_sc_hd__xor2_2 _16213_ (.A(_03560_),
    .B(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__nand2_2 _16214_ (.A(\systolic_inst.B_outs[12][5] ),
    .B(\systolic_inst.A_outs[12][5] ),
    .Y(_03597_));
 sky130_fd_sc_hd__and4b_2 _16215_ (.A_N(\systolic_inst.A_outs[12][3] ),
    .B(\systolic_inst.A_outs[12][4] ),
    .C(\systolic_inst.B_outs[12][6] ),
    .D(\systolic_inst.B_outs[12][7] ),
    .X(_03598_));
 sky130_fd_sc_hd__o2bb2a_2 _16216_ (.A1_N(\systolic_inst.A_outs[12][4] ),
    .A2_N(\systolic_inst.B_outs[12][6] ),
    .B1(_11260_),
    .B2(\systolic_inst.A_outs[12][3] ),
    .X(_03599_));
 sky130_fd_sc_hd__nor2_2 _16217_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__xnor2_2 _16218_ (.A(_03597_),
    .B(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__o21ba_2 _16219_ (.A1(_03565_),
    .A2(_03567_),
    .B1_N(_03566_),
    .X(_03602_));
 sky130_fd_sc_hd__nand2b_2 _16220_ (.A_N(_03602_),
    .B(_03601_),
    .Y(_03603_));
 sky130_fd_sc_hd__xnor2_2 _16221_ (.A(_03601_),
    .B(_03602_),
    .Y(_03604_));
 sky130_fd_sc_hd__nand2_2 _16222_ (.A(_03596_),
    .B(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__or2_2 _16223_ (.A(_03596_),
    .B(_03604_),
    .X(_03606_));
 sky130_fd_sc_hd__nand2_2 _16224_ (.A(_03605_),
    .B(_03606_),
    .Y(_03607_));
 sky130_fd_sc_hd__a21bo_2 _16225_ (.A1(_03564_),
    .A2(_03572_),
    .B1_N(_03571_),
    .X(_03608_));
 sky130_fd_sc_hd__nand2b_2 _16226_ (.A_N(_03607_),
    .B(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__xor2_2 _16227_ (.A(_03607_),
    .B(_03608_),
    .X(_03610_));
 sky130_fd_sc_hd__xor2_2 _16228_ (.A(_03592_),
    .B(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__o21a_2 _16229_ (.A1(_03559_),
    .A2(_03576_),
    .B1(_03574_),
    .X(_03612_));
 sky130_fd_sc_hd__nand2b_2 _16230_ (.A_N(_03612_),
    .B(_03611_),
    .Y(_03613_));
 sky130_fd_sc_hd__xnor2_2 _16231_ (.A(_03611_),
    .B(_03612_),
    .Y(_03614_));
 sky130_fd_sc_hd__nand2_2 _16232_ (.A(_03557_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__or2_2 _16233_ (.A(_03557_),
    .B(_03614_),
    .X(_03616_));
 sky130_fd_sc_hd__nand2_2 _16234_ (.A(_03615_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__a21boi_2 _16235_ (.A1(_03555_),
    .A2(_03580_),
    .B1_N(_03579_),
    .Y(_03618_));
 sky130_fd_sc_hd__nor2_2 _16236_ (.A(_03617_),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__inv_2 _16237_ (.A(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__xnor2_2 _16238_ (.A(_03617_),
    .B(_03618_),
    .Y(_03621_));
 sky130_fd_sc_hd__a21oi_2 _16239_ (.A1(_03551_),
    .A2(_03585_),
    .B1(_03582_),
    .Y(_03622_));
 sky130_fd_sc_hd__o211ai_2 _16240_ (.A1(_03548_),
    .A2(_03584_),
    .B1(_03621_),
    .C1(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__a311o_2 _16241_ (.A1(_03548_),
    .A2(_03552_),
    .A3(_03583_),
    .B1(_03584_),
    .C1(_03621_),
    .X(_03624_));
 sky130_fd_sc_hd__and3_2 _16242_ (.A(\systolic_inst.ce_local ),
    .B(_03623_),
    .C(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__a21o_2 _16243_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[10] ),
    .B1(_03625_),
    .X(_01164_));
 sky130_fd_sc_hd__o2bb2a_2 _16244_ (.A1_N(\systolic_inst.A_outs[12][6] ),
    .A2_N(_03594_),
    .B1(_03595_),
    .B2(_03560_),
    .X(_03626_));
 sky130_fd_sc_hd__or2_2 _16245_ (.A(_03517_),
    .B(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__nand2_2 _16246_ (.A(_03517_),
    .B(_03626_),
    .Y(_03628_));
 sky130_fd_sc_hd__nand2_2 _16247_ (.A(_03627_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__or2_2 _16248_ (.A(\systolic_inst.B_outs[12][3] ),
    .B(\systolic_inst.B_outs[12][4] ),
    .X(_03630_));
 sky130_fd_sc_hd__and3b_2 _16249_ (.A_N(_03594_),
    .B(_03630_),
    .C(\systolic_inst.A_outs[12][7] ),
    .X(_03631_));
 sky130_fd_sc_hd__xnor2_2 _16250_ (.A(_03560_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__nand2_2 _16251_ (.A(\systolic_inst.B_outs[12][5] ),
    .B(\systolic_inst.A_outs[12][6] ),
    .Y(_03633_));
 sky130_fd_sc_hd__and4b_2 _16252_ (.A_N(\systolic_inst.A_outs[12][4] ),
    .B(\systolic_inst.A_outs[12][5] ),
    .C(\systolic_inst.B_outs[12][6] ),
    .D(\systolic_inst.B_outs[12][7] ),
    .X(_03634_));
 sky130_fd_sc_hd__o2bb2a_2 _16253_ (.A1_N(\systolic_inst.A_outs[12][5] ),
    .A2_N(\systolic_inst.B_outs[12][6] ),
    .B1(_11260_),
    .B2(\systolic_inst.A_outs[12][4] ),
    .X(_03635_));
 sky130_fd_sc_hd__nor2_2 _16254_ (.A(_03634_),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__xnor2_2 _16255_ (.A(_03633_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__o21ba_2 _16256_ (.A1(_03597_),
    .A2(_03599_),
    .B1_N(_03598_),
    .X(_03638_));
 sky130_fd_sc_hd__nand2b_2 _16257_ (.A_N(_03638_),
    .B(_03637_),
    .Y(_03639_));
 sky130_fd_sc_hd__xnor2_2 _16258_ (.A(_03637_),
    .B(_03638_),
    .Y(_03640_));
 sky130_fd_sc_hd__nand2_2 _16259_ (.A(_03632_),
    .B(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__xnor2_2 _16260_ (.A(_03632_),
    .B(_03640_),
    .Y(_03642_));
 sky130_fd_sc_hd__a21o_2 _16261_ (.A1(_03603_),
    .A2(_03605_),
    .B1(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__nand3_2 _16262_ (.A(_03603_),
    .B(_03605_),
    .C(_03642_),
    .Y(_03644_));
 sky130_fd_sc_hd__nand2_2 _16263_ (.A(_03643_),
    .B(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__xor2_2 _16264_ (.A(_03629_),
    .B(_03645_),
    .X(_03646_));
 sky130_fd_sc_hd__o21a_2 _16265_ (.A1(_03592_),
    .A2(_03610_),
    .B1(_03609_),
    .X(_03647_));
 sky130_fd_sc_hd__and2b_2 _16266_ (.A_N(_03647_),
    .B(_03646_),
    .X(_03648_));
 sky130_fd_sc_hd__xnor2_2 _16267_ (.A(_03646_),
    .B(_03647_),
    .Y(_03649_));
 sky130_fd_sc_hd__xnor2_2 _16268_ (.A(_03590_),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__and3_2 _16269_ (.A(_03613_),
    .B(_03615_),
    .C(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__a21oi_2 _16270_ (.A1(_03613_),
    .A2(_03615_),
    .B1(_03650_),
    .Y(_03652_));
 sky130_fd_sc_hd__inv_2 _16271_ (.A(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__nor2_2 _16272_ (.A(_03651_),
    .B(_03652_),
    .Y(_03654_));
 sky130_fd_sc_hd__and2_2 _16273_ (.A(_03620_),
    .B(_03624_),
    .X(_03655_));
 sky130_fd_sc_hd__xnor2_2 _16274_ (.A(_03654_),
    .B(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__mux2_1 _16275_ (.A0(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[11] ),
    .A1(_03656_),
    .S(\systolic_inst.ce_local ),
    .X(_01165_));
 sky130_fd_sc_hd__a31o_2 _16276_ (.A1(\systolic_inst.B_outs[12][2] ),
    .A2(\systolic_inst.A_outs[12][7] ),
    .A3(_03630_),
    .B1(_03594_),
    .X(_03657_));
 sky130_fd_sc_hd__or2_2 _16277_ (.A(_03516_),
    .B(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__nand2_2 _16278_ (.A(_03516_),
    .B(_03657_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand2_2 _16279_ (.A(_03658_),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__o2bb2a_2 _16280_ (.A1_N(\systolic_inst.B_outs[12][6] ),
    .A2_N(\systolic_inst.A_outs[12][6] ),
    .B1(_11260_),
    .B2(\systolic_inst.A_outs[12][5] ),
    .X(_03661_));
 sky130_fd_sc_hd__and4b_2 _16281_ (.A_N(\systolic_inst.A_outs[12][5] ),
    .B(\systolic_inst.B_outs[12][6] ),
    .C(\systolic_inst.A_outs[12][6] ),
    .D(\systolic_inst.B_outs[12][7] ),
    .X(_03662_));
 sky130_fd_sc_hd__nor2_2 _16282_ (.A(_03661_),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__nand2_2 _16283_ (.A(\systolic_inst.B_outs[12][5] ),
    .B(\systolic_inst.A_outs[12][7] ),
    .Y(_03664_));
 sky130_fd_sc_hd__and3_2 _16284_ (.A(\systolic_inst.B_outs[12][5] ),
    .B(\systolic_inst.A_outs[12][7] ),
    .C(_03663_),
    .X(_03665_));
 sky130_fd_sc_hd__xnor2_2 _16285_ (.A(_03663_),
    .B(_03664_),
    .Y(_03666_));
 sky130_fd_sc_hd__o21ba_2 _16286_ (.A1(_03633_),
    .A2(_03635_),
    .B1_N(_03634_),
    .X(_03667_));
 sky130_fd_sc_hd__nand2b_2 _16287_ (.A_N(_03667_),
    .B(_03666_),
    .Y(_03668_));
 sky130_fd_sc_hd__xnor2_2 _16288_ (.A(_03666_),
    .B(_03667_),
    .Y(_03669_));
 sky130_fd_sc_hd__xnor2_2 _16289_ (.A(_03632_),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__a21o_2 _16290_ (.A1(_03639_),
    .A2(_03641_),
    .B1(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__nand3_2 _16291_ (.A(_03639_),
    .B(_03641_),
    .C(_03670_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_2 _16292_ (.A(_03671_),
    .B(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__xor2_2 _16293_ (.A(_03660_),
    .B(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__o21a_2 _16294_ (.A1(_03629_),
    .A2(_03645_),
    .B1(_03643_),
    .X(_03675_));
 sky130_fd_sc_hd__and2b_2 _16295_ (.A_N(_03675_),
    .B(_03674_),
    .X(_03676_));
 sky130_fd_sc_hd__xnor2_2 _16296_ (.A(_03674_),
    .B(_03675_),
    .Y(_03677_));
 sky130_fd_sc_hd__and2b_2 _16297_ (.A_N(_03627_),
    .B(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__xor2_2 _16298_ (.A(_03627_),
    .B(_03677_),
    .X(_03679_));
 sky130_fd_sc_hd__a21oi_2 _16299_ (.A1(_03590_),
    .A2(_03649_),
    .B1(_03648_),
    .Y(_03680_));
 sky130_fd_sc_hd__nor2_2 _16300_ (.A(_03679_),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__and2_2 _16301_ (.A(_03679_),
    .B(_03680_),
    .X(_03682_));
 sky130_fd_sc_hd__nor2_2 _16302_ (.A(_03681_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__inv_2 _16303_ (.A(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__a31o_2 _16304_ (.A1(_03620_),
    .A2(_03624_),
    .A3(_03653_),
    .B1(_03651_),
    .X(_03685_));
 sky130_fd_sc_hd__a311oi_2 _16305_ (.A1(_03620_),
    .A2(_03624_),
    .A3(_03653_),
    .B1(_03684_),
    .C1(_03651_),
    .Y(_03686_));
 sky130_fd_sc_hd__and2_2 _16306_ (.A(_03684_),
    .B(_03685_),
    .X(_03687_));
 sky130_fd_sc_hd__nor2_2 _16307_ (.A(_03686_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__mux2_1 _16308_ (.A0(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[12] ),
    .A1(_03688_),
    .S(\systolic_inst.ce_local ),
    .X(_01166_));
 sky130_fd_sc_hd__nand2_2 _16309_ (.A(\systolic_inst.B_outs[12][6] ),
    .B(\systolic_inst.A_outs[12][7] ),
    .Y(_03689_));
 sky130_fd_sc_hd__nor2_2 _16310_ (.A(\systolic_inst.A_outs[12][6] ),
    .B(_11260_),
    .Y(_03690_));
 sky130_fd_sc_hd__xnor2_2 _16311_ (.A(_03689_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__nand2b_2 _16312_ (.A_N(_03664_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__xnor2_2 _16313_ (.A(_03664_),
    .B(_03691_),
    .Y(_03693_));
 sky130_fd_sc_hd__o21ai_2 _16314_ (.A1(_03662_),
    .A2(_03665_),
    .B1(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__or3_2 _16315_ (.A(_03662_),
    .B(_03665_),
    .C(_03693_),
    .X(_03695_));
 sky130_fd_sc_hd__and2_2 _16316_ (.A(_03694_),
    .B(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__nand2_2 _16317_ (.A(_03632_),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__or2_2 _16318_ (.A(_03632_),
    .B(_03696_),
    .X(_03698_));
 sky130_fd_sc_hd__nand2_2 _16319_ (.A(_03697_),
    .B(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__a21bo_2 _16320_ (.A1(_03632_),
    .A2(_03669_),
    .B1_N(_03668_),
    .X(_03700_));
 sky130_fd_sc_hd__nand2b_2 _16321_ (.A_N(_03699_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__xor2_2 _16322_ (.A(_03699_),
    .B(_03700_),
    .X(_03702_));
 sky130_fd_sc_hd__xor2_2 _16323_ (.A(_03660_),
    .B(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__o21a_2 _16324_ (.A1(_03660_),
    .A2(_03673_),
    .B1(_03671_),
    .X(_03704_));
 sky130_fd_sc_hd__and2b_2 _16325_ (.A_N(_03704_),
    .B(_03703_),
    .X(_03705_));
 sky130_fd_sc_hd__and2b_2 _16326_ (.A_N(_03703_),
    .B(_03704_),
    .X(_03706_));
 sky130_fd_sc_hd__nor2_2 _16327_ (.A(_03705_),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__xnor2_2 _16328_ (.A(_03659_),
    .B(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__o21a_2 _16329_ (.A1(_03676_),
    .A2(_03678_),
    .B1(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__or3_2 _16330_ (.A(_03676_),
    .B(_03678_),
    .C(_03708_),
    .X(_03710_));
 sky130_fd_sc_hd__and2b_2 _16331_ (.A_N(_03709_),
    .B(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__nor2_2 _16332_ (.A(_03681_),
    .B(_03686_),
    .Y(_03712_));
 sky130_fd_sc_hd__xnor2_2 _16333_ (.A(_03711_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__mux2_1 _16334_ (.A0(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[13] ),
    .A1(_03713_),
    .S(\systolic_inst.ce_local ),
    .X(_01167_));
 sky130_fd_sc_hd__o211ai_2 _16335_ (.A1(_11260_),
    .A2(\systolic_inst.A_outs[12][7] ),
    .B1(_03664_),
    .C1(_03689_),
    .Y(_03714_));
 sky130_fd_sc_hd__o311a_2 _16336_ (.A1(\systolic_inst.A_outs[12][6] ),
    .A2(_11260_),
    .A3(_03689_),
    .B1(_03692_),
    .C1(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__a31o_2 _16337_ (.A1(\systolic_inst.B_outs[12][5] ),
    .A2(\systolic_inst.B_outs[12][6] ),
    .A3(\systolic_inst.A_outs[12][7] ),
    .B1(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__or2_2 _16338_ (.A(_03632_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__nand2_2 _16339_ (.A(_03632_),
    .B(_03716_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_2 _16340_ (.A(_03717_),
    .B(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__a21oi_2 _16341_ (.A1(_03694_),
    .A2(_03697_),
    .B1(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__and3_2 _16342_ (.A(_03694_),
    .B(_03697_),
    .C(_03719_),
    .X(_03721_));
 sky130_fd_sc_hd__nor2_2 _16343_ (.A(_03720_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__xnor2_2 _16344_ (.A(_03660_),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__o21a_2 _16345_ (.A1(_03660_),
    .A2(_03702_),
    .B1(_03701_),
    .X(_03724_));
 sky130_fd_sc_hd__and2b_2 _16346_ (.A_N(_03724_),
    .B(_03723_),
    .X(_03725_));
 sky130_fd_sc_hd__and2b_2 _16347_ (.A_N(_03723_),
    .B(_03724_),
    .X(_03726_));
 sky130_fd_sc_hd__nor2_2 _16348_ (.A(_03725_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__xnor2_2 _16349_ (.A(_03659_),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__o21ba_2 _16350_ (.A1(_03659_),
    .A2(_03706_),
    .B1_N(_03705_),
    .X(_03729_));
 sky130_fd_sc_hd__and2b_2 _16351_ (.A_N(_03729_),
    .B(_03728_),
    .X(_03730_));
 sky130_fd_sc_hd__xnor2_2 _16352_ (.A(_03728_),
    .B(_03729_),
    .Y(_03731_));
 sky130_fd_sc_hd__o31a_2 _16353_ (.A1(_03681_),
    .A2(_03686_),
    .A3(_03709_),
    .B1(_03710_),
    .X(_03732_));
 sky130_fd_sc_hd__or2_2 _16354_ (.A(_03731_),
    .B(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__o311a_2 _16355_ (.A1(_03681_),
    .A2(_03686_),
    .A3(_03709_),
    .B1(_03710_),
    .C1(_03731_),
    .X(_03734_));
 sky130_fd_sc_hd__nor2_2 _16356_ (.A(_11258_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__a22o_2 _16357_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[14] ),
    .B1(_03733_),
    .B2(_03735_),
    .X(_01168_));
 sky130_fd_sc_hd__a31o_2 _16358_ (.A1(_03516_),
    .A2(_03657_),
    .A3(_03727_),
    .B1(_03725_),
    .X(_03736_));
 sky130_fd_sc_hd__a31o_2 _16359_ (.A1(_03658_),
    .A2(_03659_),
    .A3(_03722_),
    .B1(_03720_),
    .X(_03737_));
 sky130_fd_sc_hd__xnor2_2 _16360_ (.A(_03658_),
    .B(_03717_),
    .Y(_03738_));
 sky130_fd_sc_hd__xnor2_2 _16361_ (.A(_03737_),
    .B(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__xnor2_2 _16362_ (.A(_03736_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__or3_2 _16363_ (.A(_11258_),
    .B(_03730_),
    .C(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__a2bb2o_2 _16364_ (.A1_N(_03741_),
    .A2_N(_03734_),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B2(_11258_),
    .X(_01169_));
 sky130_fd_sc_hd__a21o_2 _16365_ (.A1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[12][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_03742_));
 sky130_fd_sc_hd__a21oi_2 _16366_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[12][0] ),
    .Y(_03743_));
 sky130_fd_sc_hd__a21oi_2 _16367_ (.A1(\systolic_inst.ce_local ),
    .A2(_03742_),
    .B1(_03743_),
    .Y(_01170_));
 sky130_fd_sc_hd__nand2_2 _16368_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[12][1] ),
    .Y(_03744_));
 sky130_fd_sc_hd__inv_2 _16369_ (.A(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__or2_2 _16370_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[12][1] ),
    .X(_03746_));
 sky130_fd_sc_hd__and4_2 _16371_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[12][0] ),
    .C(_03744_),
    .D(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__inv_2 _16372_ (.A(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__a22o_2 _16373_ (.A1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[12][0] ),
    .B1(_03744_),
    .B2(_03746_),
    .X(_03749_));
 sky130_fd_sc_hd__a32o_2 _16374_ (.A1(_11712_),
    .A2(_03748_),
    .A3(_03749_),
    .B1(\systolic_inst.acc_wires[12][1] ),
    .B2(_11258_),
    .X(_01171_));
 sky130_fd_sc_hd__nand2_2 _16375_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[12][2] ),
    .Y(_03750_));
 sky130_fd_sc_hd__inv_2 _16376_ (.A(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__or2_2 _16377_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[12][2] ),
    .X(_03752_));
 sky130_fd_sc_hd__a211o_2 _16378_ (.A1(_03750_),
    .A2(_03752_),
    .B1(_03745_),
    .C1(_03747_),
    .X(_03753_));
 sky130_fd_sc_hd__o211a_2 _16379_ (.A1(_03745_),
    .A2(_03747_),
    .B1(_03750_),
    .C1(_03752_),
    .X(_03754_));
 sky130_fd_sc_hd__inv_2 _16380_ (.A(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__a32o_2 _16381_ (.A1(_11712_),
    .A2(_03753_),
    .A3(_03755_),
    .B1(\systolic_inst.acc_wires[12][2] ),
    .B2(_11258_),
    .X(_01172_));
 sky130_fd_sc_hd__nand2_2 _16382_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[12][3] ),
    .Y(_03756_));
 sky130_fd_sc_hd__inv_2 _16383_ (.A(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__or2_2 _16384_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[12][3] ),
    .X(_03758_));
 sky130_fd_sc_hd__a211o_2 _16385_ (.A1(_03756_),
    .A2(_03758_),
    .B1(_03751_),
    .C1(_03754_),
    .X(_03759_));
 sky130_fd_sc_hd__o211a_2 _16386_ (.A1(_03751_),
    .A2(_03754_),
    .B1(_03756_),
    .C1(_03758_),
    .X(_03760_));
 sky130_fd_sc_hd__inv_2 _16387_ (.A(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__a32o_2 _16388_ (.A1(_11712_),
    .A2(_03759_),
    .A3(_03761_),
    .B1(\systolic_inst.acc_wires[12][3] ),
    .B2(_11258_),
    .X(_01173_));
 sky130_fd_sc_hd__nand2_2 _16389_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[12][4] ),
    .Y(_03762_));
 sky130_fd_sc_hd__inv_2 _16390_ (.A(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__or2_2 _16391_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[12][4] ),
    .X(_03764_));
 sky130_fd_sc_hd__a211o_2 _16392_ (.A1(_03762_),
    .A2(_03764_),
    .B1(_03757_),
    .C1(_03760_),
    .X(_03765_));
 sky130_fd_sc_hd__o211a_2 _16393_ (.A1(_03757_),
    .A2(_03760_),
    .B1(_03762_),
    .C1(_03764_),
    .X(_03766_));
 sky130_fd_sc_hd__inv_2 _16394_ (.A(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__a32o_2 _16395_ (.A1(_11712_),
    .A2(_03765_),
    .A3(_03767_),
    .B1(\systolic_inst.acc_wires[12][4] ),
    .B2(_11258_),
    .X(_01174_));
 sky130_fd_sc_hd__nand2_2 _16396_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[12][5] ),
    .Y(_03768_));
 sky130_fd_sc_hd__inv_2 _16397_ (.A(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__or2_2 _16398_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[12][5] ),
    .X(_03770_));
 sky130_fd_sc_hd__a211o_2 _16399_ (.A1(_03768_),
    .A2(_03770_),
    .B1(_03763_),
    .C1(_03766_),
    .X(_03771_));
 sky130_fd_sc_hd__o211a_2 _16400_ (.A1(_03763_),
    .A2(_03766_),
    .B1(_03768_),
    .C1(_03770_),
    .X(_03772_));
 sky130_fd_sc_hd__inv_2 _16401_ (.A(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__a32o_2 _16402_ (.A1(_11712_),
    .A2(_03771_),
    .A3(_03773_),
    .B1(\systolic_inst.acc_wires[12][5] ),
    .B2(_11258_),
    .X(_01175_));
 sky130_fd_sc_hd__nand2_2 _16403_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[12][6] ),
    .Y(_03774_));
 sky130_fd_sc_hd__inv_2 _16404_ (.A(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__or2_2 _16405_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[12][6] ),
    .X(_03776_));
 sky130_fd_sc_hd__a211o_2 _16406_ (.A1(_03774_),
    .A2(_03776_),
    .B1(_03769_),
    .C1(_03772_),
    .X(_03777_));
 sky130_fd_sc_hd__o211a_2 _16407_ (.A1(_03769_),
    .A2(_03772_),
    .B1(_03774_),
    .C1(_03776_),
    .X(_03778_));
 sky130_fd_sc_hd__inv_2 _16408_ (.A(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__a32o_2 _16409_ (.A1(_11712_),
    .A2(_03777_),
    .A3(_03779_),
    .B1(\systolic_inst.acc_wires[12][6] ),
    .B2(_11258_),
    .X(_01176_));
 sky130_fd_sc_hd__nand2_2 _16410_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[12][7] ),
    .Y(_03780_));
 sky130_fd_sc_hd__or2_2 _16411_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[12][7] ),
    .X(_03781_));
 sky130_fd_sc_hd__a211o_2 _16412_ (.A1(_03780_),
    .A2(_03781_),
    .B1(_03775_),
    .C1(_03778_),
    .X(_03782_));
 sky130_fd_sc_hd__o211ai_2 _16413_ (.A1(_03775_),
    .A2(_03778_),
    .B1(_03780_),
    .C1(_03781_),
    .Y(_03783_));
 sky130_fd_sc_hd__a32o_2 _16414_ (.A1(_11712_),
    .A2(_03782_),
    .A3(_03783_),
    .B1(\systolic_inst.acc_wires[12][7] ),
    .B2(_11258_),
    .X(_01177_));
 sky130_fd_sc_hd__nand2_2 _16415_ (.A(_03780_),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__xor2_2 _16416_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[12][8] ),
    .X(_03785_));
 sky130_fd_sc_hd__and2_2 _16417_ (.A(_03784_),
    .B(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__o21ai_2 _16418_ (.A1(_03784_),
    .A2(_03785_),
    .B1(_11712_),
    .Y(_03787_));
 sky130_fd_sc_hd__a2bb2o_2 _16419_ (.A1_N(_03787_),
    .A2_N(_03786_),
    .B1(\systolic_inst.acc_wires[12][8] ),
    .B2(_11258_),
    .X(_01178_));
 sky130_fd_sc_hd__nor2_2 _16420_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[12][9] ),
    .Y(_03788_));
 sky130_fd_sc_hd__and2_2 _16421_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[12][9] ),
    .X(_03789_));
 sky130_fd_sc_hd__nor2_2 _16422_ (.A(_03788_),
    .B(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__a211o_2 _16423_ (.A1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[12][8] ),
    .B1(_03786_),
    .C1(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__and3_2 _16424_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[12][8] ),
    .C(_03790_),
    .X(_03792_));
 sky130_fd_sc_hd__a21oi_2 _16425_ (.A1(_03786_),
    .A2(_03790_),
    .B1(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__a32o_2 _16426_ (.A1(_11712_),
    .A2(_03791_),
    .A3(_03793_),
    .B1(\systolic_inst.acc_wires[12][9] ),
    .B2(_11258_),
    .X(_01179_));
 sky130_fd_sc_hd__and2_2 _16427_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[12][10] ),
    .X(_03794_));
 sky130_fd_sc_hd__nor2_2 _16428_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[12][10] ),
    .Y(_03795_));
 sky130_fd_sc_hd__nor2_2 _16429_ (.A(_03794_),
    .B(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__or2_2 _16430_ (.A(_03789_),
    .B(_03792_),
    .X(_03797_));
 sky130_fd_sc_hd__a31o_2 _16431_ (.A1(_03784_),
    .A2(_03785_),
    .A3(_03790_),
    .B1(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__or2_2 _16432_ (.A(_03796_),
    .B(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__nand2_2 _16433_ (.A(_03796_),
    .B(_03798_),
    .Y(_03800_));
 sky130_fd_sc_hd__a32o_2 _16434_ (.A1(_11712_),
    .A2(_03799_),
    .A3(_03800_),
    .B1(\systolic_inst.acc_wires[12][10] ),
    .B2(_11258_),
    .X(_01180_));
 sky130_fd_sc_hd__or2_2 _16435_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[12][11] ),
    .X(_03801_));
 sky130_fd_sc_hd__nand2_2 _16436_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[12][11] ),
    .Y(_03802_));
 sky130_fd_sc_hd__a21o_2 _16437_ (.A1(_03796_),
    .A2(_03798_),
    .B1(_03794_),
    .X(_03803_));
 sky130_fd_sc_hd__a21oi_2 _16438_ (.A1(_03801_),
    .A2(_03802_),
    .B1(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__a31o_2 _16439_ (.A1(_03801_),
    .A2(_03802_),
    .A3(_03803_),
    .B1(_11713_),
    .X(_03805_));
 sky130_fd_sc_hd__a2bb2o_2 _16440_ (.A1_N(_03805_),
    .A2_N(_03804_),
    .B1(\systolic_inst.acc_wires[12][11] ),
    .B2(_11258_),
    .X(_01181_));
 sky130_fd_sc_hd__and3_2 _16441_ (.A(_03796_),
    .B(_03801_),
    .C(_03802_),
    .X(_03806_));
 sky130_fd_sc_hd__and2_2 _16442_ (.A(_03797_),
    .B(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__nand3_2 _16443_ (.A(_03785_),
    .B(_03790_),
    .C(_03806_),
    .Y(_03808_));
 sky130_fd_sc_hd__a21oi_2 _16444_ (.A1(_03780_),
    .A2(_03783_),
    .B1(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__a21bo_2 _16445_ (.A1(_03794_),
    .A2(_03801_),
    .B1_N(_03802_),
    .X(_03810_));
 sky130_fd_sc_hd__or3_2 _16446_ (.A(_03807_),
    .B(_03809_),
    .C(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__nor2_2 _16447_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[12][12] ),
    .Y(_03812_));
 sky130_fd_sc_hd__nand2_2 _16448_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[12][12] ),
    .Y(_03813_));
 sky130_fd_sc_hd__inv_2 _16449_ (.A(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__nor2_2 _16450_ (.A(_03812_),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__or2_2 _16451_ (.A(_03811_),
    .B(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__and2_2 _16452_ (.A(_03811_),
    .B(_03815_),
    .X(_03817_));
 sky130_fd_sc_hd__inv_2 _16453_ (.A(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__a32o_2 _16454_ (.A1(_11712_),
    .A2(_03816_),
    .A3(_03818_),
    .B1(\systolic_inst.acc_wires[12][12] ),
    .B2(_11258_),
    .X(_01182_));
 sky130_fd_sc_hd__or2_2 _16455_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[12][13] ),
    .X(_03819_));
 sky130_fd_sc_hd__nand2_2 _16456_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[12][13] ),
    .Y(_03820_));
 sky130_fd_sc_hd__and2_2 _16457_ (.A(_03819_),
    .B(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__o21ai_2 _16458_ (.A1(_03814_),
    .A2(_03817_),
    .B1(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__o31a_2 _16459_ (.A1(_03814_),
    .A2(_03817_),
    .A3(_03821_),
    .B1(_11712_),
    .X(_03823_));
 sky130_fd_sc_hd__a22o_2 _16460_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[12][13] ),
    .B1(_03822_),
    .B2(_03823_),
    .X(_01183_));
 sky130_fd_sc_hd__or2_2 _16461_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[12][14] ),
    .X(_03824_));
 sky130_fd_sc_hd__nand2_2 _16462_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[12][14] ),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2_2 _16463_ (.A(_03824_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand3_2 _16464_ (.A(_03820_),
    .B(_03822_),
    .C(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__a21o_2 _16465_ (.A1(_03820_),
    .A2(_03822_),
    .B1(_03826_),
    .X(_03828_));
 sky130_fd_sc_hd__a32o_2 _16466_ (.A1(_11712_),
    .A2(_03827_),
    .A3(_03828_),
    .B1(\systolic_inst.acc_wires[12][14] ),
    .B2(_11258_),
    .X(_01184_));
 sky130_fd_sc_hd__nor2_2 _16467_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][15] ),
    .Y(_03829_));
 sky130_fd_sc_hd__nand2_2 _16468_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][15] ),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2b_2 _16469_ (.A_N(_03829_),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__a21oi_2 _16470_ (.A1(_03825_),
    .A2(_03828_),
    .B1(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__a31o_2 _16471_ (.A1(_03825_),
    .A2(_03828_),
    .A3(_03831_),
    .B1(_11713_),
    .X(_03833_));
 sky130_fd_sc_hd__a2bb2o_2 _16472_ (.A1_N(_03833_),
    .A2_N(_03832_),
    .B1(\systolic_inst.acc_wires[12][15] ),
    .B2(_11258_),
    .X(_01185_));
 sky130_fd_sc_hd__nor2_2 _16473_ (.A(_03826_),
    .B(_03831_),
    .Y(_03834_));
 sky130_fd_sc_hd__inv_2 _16474_ (.A(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__and2_2 _16475_ (.A(_03821_),
    .B(_03834_),
    .X(_03836_));
 sky130_fd_sc_hd__o311a_2 _16476_ (.A1(_03807_),
    .A2(_03809_),
    .A3(_03810_),
    .B1(_03815_),
    .C1(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__a21boi_2 _16477_ (.A1(_03814_),
    .A2(_03819_),
    .B1_N(_03820_),
    .Y(_03838_));
 sky130_fd_sc_hd__o221a_2 _16478_ (.A1(_03825_),
    .A2(_03829_),
    .B1(_03835_),
    .B2(_03838_),
    .C1(_03830_),
    .X(_03839_));
 sky130_fd_sc_hd__inv_2 _16479_ (.A(_03839_),
    .Y(_03840_));
 sky130_fd_sc_hd__or2_2 _16480_ (.A(_03837_),
    .B(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__nor2_2 _16481_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][16] ),
    .Y(_03842_));
 sky130_fd_sc_hd__and2_2 _16482_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][16] ),
    .X(_03843_));
 sky130_fd_sc_hd__nor2_2 _16483_ (.A(_03842_),
    .B(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__and2_2 _16484_ (.A(_03841_),
    .B(_03844_),
    .X(_03845_));
 sky130_fd_sc_hd__o21ai_2 _16485_ (.A1(_03841_),
    .A2(_03844_),
    .B1(_11712_),
    .Y(_03846_));
 sky130_fd_sc_hd__a2bb2o_2 _16486_ (.A1_N(_03846_),
    .A2_N(_03845_),
    .B1(\systolic_inst.acc_wires[12][16] ),
    .B2(_11258_),
    .X(_01186_));
 sky130_fd_sc_hd__xor2_2 _16487_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][17] ),
    .X(_03847_));
 sky130_fd_sc_hd__or3_2 _16488_ (.A(_03843_),
    .B(_03845_),
    .C(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__o21ai_2 _16489_ (.A1(_03843_),
    .A2(_03845_),
    .B1(_03847_),
    .Y(_03849_));
 sky130_fd_sc_hd__a32o_2 _16490_ (.A1(_11712_),
    .A2(_03848_),
    .A3(_03849_),
    .B1(\systolic_inst.acc_wires[12][17] ),
    .B2(_11258_),
    .X(_01187_));
 sky130_fd_sc_hd__or2_2 _16491_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][18] ),
    .X(_03850_));
 sky130_fd_sc_hd__nand2_2 _16492_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][18] ),
    .Y(_03851_));
 sky130_fd_sc_hd__nand2_2 _16493_ (.A(_03850_),
    .B(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__o21ai_2 _16494_ (.A1(\systolic_inst.acc_wires[12][16] ),
    .A2(\systolic_inst.acc_wires[12][17] ),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_2 _16495_ (.A(_03845_),
    .B(_03847_),
    .Y(_03854_));
 sky130_fd_sc_hd__a21o_2 _16496_ (.A1(_03853_),
    .A2(_03854_),
    .B1(_03852_),
    .X(_03855_));
 sky130_fd_sc_hd__nand3_2 _16497_ (.A(_03852_),
    .B(_03853_),
    .C(_03854_),
    .Y(_03856_));
 sky130_fd_sc_hd__a32o_2 _16498_ (.A1(_11712_),
    .A2(_03855_),
    .A3(_03856_),
    .B1(\systolic_inst.acc_wires[12][18] ),
    .B2(_11258_),
    .X(_01188_));
 sky130_fd_sc_hd__xnor2_2 _16499_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][19] ),
    .Y(_03857_));
 sky130_fd_sc_hd__a21oi_2 _16500_ (.A1(_03851_),
    .A2(_03855_),
    .B1(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__a31o_2 _16501_ (.A1(_03851_),
    .A2(_03855_),
    .A3(_03857_),
    .B1(_11713_),
    .X(_03859_));
 sky130_fd_sc_hd__a2bb2o_2 _16502_ (.A1_N(_03859_),
    .A2_N(_03858_),
    .B1(\systolic_inst.acc_wires[12][19] ),
    .B2(_11258_),
    .X(_01189_));
 sky130_fd_sc_hd__xor2_2 _16503_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][20] ),
    .X(_03860_));
 sky130_fd_sc_hd__nor2_2 _16504_ (.A(_03852_),
    .B(_03857_),
    .Y(_03861_));
 sky130_fd_sc_hd__and3_2 _16505_ (.A(_03844_),
    .B(_03847_),
    .C(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__o21a_2 _16506_ (.A1(_03837_),
    .A2(_03840_),
    .B1(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__o41a_2 _16507_ (.A1(\systolic_inst.acc_wires[12][16] ),
    .A2(\systolic_inst.acc_wires[12][17] ),
    .A3(\systolic_inst.acc_wires[12][18] ),
    .A4(\systolic_inst.acc_wires[12][19] ),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .X(_03864_));
 sky130_fd_sc_hd__or3_2 _16508_ (.A(_03860_),
    .B(_03863_),
    .C(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__o21ai_2 _16509_ (.A1(_03863_),
    .A2(_03864_),
    .B1(_03860_),
    .Y(_03866_));
 sky130_fd_sc_hd__a32o_2 _16510_ (.A1(_11712_),
    .A2(_03865_),
    .A3(_03866_),
    .B1(\systolic_inst.acc_wires[12][20] ),
    .B2(_11258_),
    .X(_01190_));
 sky130_fd_sc_hd__xor2_2 _16511_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][21] ),
    .X(_03867_));
 sky130_fd_sc_hd__a21bo_2 _16512_ (.A1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[12][20] ),
    .B1_N(_03866_),
    .X(_03868_));
 sky130_fd_sc_hd__xor2_2 _16513_ (.A(_03867_),
    .B(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__a22o_2 _16514_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[12][21] ),
    .B1(_11712_),
    .B2(_03869_),
    .X(_01191_));
 sky130_fd_sc_hd__or2_2 _16515_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][22] ),
    .X(_03870_));
 sky130_fd_sc_hd__nand2_2 _16516_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][22] ),
    .Y(_03871_));
 sky130_fd_sc_hd__and2_2 _16517_ (.A(_03870_),
    .B(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__o21a_2 _16518_ (.A1(\systolic_inst.acc_wires[12][20] ),
    .A2(\systolic_inst.acc_wires[12][21] ),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .X(_03873_));
 sky130_fd_sc_hd__and2b_2 _16519_ (.A_N(_03866_),
    .B(_03867_),
    .X(_03874_));
 sky130_fd_sc_hd__o21ai_2 _16520_ (.A1(_03873_),
    .A2(_03874_),
    .B1(_03872_),
    .Y(_03875_));
 sky130_fd_sc_hd__or3_2 _16521_ (.A(_03872_),
    .B(_03873_),
    .C(_03874_),
    .X(_03876_));
 sky130_fd_sc_hd__a32o_2 _16522_ (.A1(_11712_),
    .A2(_03875_),
    .A3(_03876_),
    .B1(\systolic_inst.acc_wires[12][22] ),
    .B2(_11258_),
    .X(_01192_));
 sky130_fd_sc_hd__xnor2_2 _16523_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][23] ),
    .Y(_03877_));
 sky130_fd_sc_hd__inv_2 _16524_ (.A(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__a21oi_2 _16525_ (.A1(_03871_),
    .A2(_03875_),
    .B1(_03877_),
    .Y(_03879_));
 sky130_fd_sc_hd__a31o_2 _16526_ (.A1(_03871_),
    .A2(_03875_),
    .A3(_03877_),
    .B1(_11713_),
    .X(_03880_));
 sky130_fd_sc_hd__a2bb2o_2 _16527_ (.A1_N(_03880_),
    .A2_N(_03879_),
    .B1(\systolic_inst.acc_wires[12][23] ),
    .B2(_11258_),
    .X(_01193_));
 sky130_fd_sc_hd__and4_2 _16528_ (.A(_03860_),
    .B(_03867_),
    .C(_03872_),
    .D(_03878_),
    .X(_03881_));
 sky130_fd_sc_hd__o21a_2 _16529_ (.A1(\systolic_inst.acc_wires[12][22] ),
    .A2(\systolic_inst.acc_wires[12][23] ),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .X(_03882_));
 sky130_fd_sc_hd__or3_2 _16530_ (.A(_03864_),
    .B(_03873_),
    .C(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__a21oi_2 _16531_ (.A1(_03863_),
    .A2(_03881_),
    .B1(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__xnor2_2 _16532_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][24] ),
    .Y(_03885_));
 sky130_fd_sc_hd__nor2_2 _16533_ (.A(_03884_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__a21o_2 _16534_ (.A1(_03884_),
    .A2(_03885_),
    .B1(_11713_),
    .X(_03887_));
 sky130_fd_sc_hd__a2bb2o_2 _16535_ (.A1_N(_03887_),
    .A2_N(_03886_),
    .B1(\systolic_inst.acc_wires[12][24] ),
    .B2(_11258_),
    .X(_01194_));
 sky130_fd_sc_hd__xor2_2 _16536_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][25] ),
    .X(_03888_));
 sky130_fd_sc_hd__a21oi_2 _16537_ (.A1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[12][24] ),
    .B1(_03886_),
    .Y(_03889_));
 sky130_fd_sc_hd__xnor2_2 _16538_ (.A(_03888_),
    .B(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__a22o_2 _16539_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[12][25] ),
    .B1(_11712_),
    .B2(_03890_),
    .X(_01195_));
 sky130_fd_sc_hd__or2_2 _16540_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][26] ),
    .X(_03891_));
 sky130_fd_sc_hd__nand2_2 _16541_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][26] ),
    .Y(_03892_));
 sky130_fd_sc_hd__and2_2 _16542_ (.A(_03891_),
    .B(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__inv_2 _16543_ (.A(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__o21a_2 _16544_ (.A1(\systolic_inst.acc_wires[12][24] ),
    .A2(\systolic_inst.acc_wires[12][25] ),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .X(_03895_));
 sky130_fd_sc_hd__a21oi_2 _16545_ (.A1(_03886_),
    .A2(_03888_),
    .B1(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__xnor2_2 _16546_ (.A(_03893_),
    .B(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__a22o_2 _16547_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[12][26] ),
    .B1(_11712_),
    .B2(_03897_),
    .X(_01196_));
 sky130_fd_sc_hd__xnor2_2 _16548_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][27] ),
    .Y(_03898_));
 sky130_fd_sc_hd__o21a_2 _16549_ (.A1(_03894_),
    .A2(_03896_),
    .B1(_03892_),
    .X(_03899_));
 sky130_fd_sc_hd__xnor2_2 _16550_ (.A(_03898_),
    .B(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__a2bb2o_2 _16551_ (.A1_N(_11713_),
    .A2_N(_03900_),
    .B1(_11258_),
    .B2(\systolic_inst.acc_wires[12][27] ),
    .X(_01197_));
 sky130_fd_sc_hd__nand2_2 _16552_ (.A(_03888_),
    .B(_03893_),
    .Y(_03901_));
 sky130_fd_sc_hd__or4_2 _16553_ (.A(_03884_),
    .B(_03885_),
    .C(_03898_),
    .D(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__o21a_2 _16554_ (.A1(\systolic_inst.acc_wires[12][26] ),
    .A2(\systolic_inst.acc_wires[12][27] ),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .X(_03903_));
 sky130_fd_sc_hd__nor2_2 _16555_ (.A(_03895_),
    .B(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__xnor2_2 _16556_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][28] ),
    .Y(_03905_));
 sky130_fd_sc_hd__a21oi_2 _16557_ (.A1(_03902_),
    .A2(_03904_),
    .B1(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__a31o_2 _16558_ (.A1(_03902_),
    .A2(_03904_),
    .A3(_03905_),
    .B1(_11713_),
    .X(_03907_));
 sky130_fd_sc_hd__a2bb2o_2 _16559_ (.A1_N(_03907_),
    .A2_N(_03906_),
    .B1(\systolic_inst.acc_wires[12][28] ),
    .B2(_11258_),
    .X(_01198_));
 sky130_fd_sc_hd__xor2_2 _16560_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][29] ),
    .X(_03908_));
 sky130_fd_sc_hd__a21oi_2 _16561_ (.A1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[12][28] ),
    .B1(_03906_),
    .Y(_03909_));
 sky130_fd_sc_hd__xnor2_2 _16562_ (.A(_03908_),
    .B(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__a22o_2 _16563_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[12][29] ),
    .B1(_11712_),
    .B2(_03910_),
    .X(_01199_));
 sky130_fd_sc_hd__o21a_2 _16564_ (.A1(\systolic_inst.acc_wires[12][28] ),
    .A2(\systolic_inst.acc_wires[12][29] ),
    .B1(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .X(_03911_));
 sky130_fd_sc_hd__a21o_2 _16565_ (.A1(_03906_),
    .A2(_03908_),
    .B1(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__nand2_2 _16566_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][30] ),
    .Y(_03913_));
 sky130_fd_sc_hd__or2_2 _16567_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][30] ),
    .X(_03914_));
 sky130_fd_sc_hd__nand2_2 _16568_ (.A(_03913_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__xnor2_2 _16569_ (.A(_03912_),
    .B(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__a22o_2 _16570_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[12][30] ),
    .B1(_11712_),
    .B2(_03916_),
    .X(_01200_));
 sky130_fd_sc_hd__a21bo_2 _16571_ (.A1(_03912_),
    .A2(_03914_),
    .B1_N(_03913_),
    .X(_03917_));
 sky130_fd_sc_hd__xnor2_2 _16572_ (.A(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[12][31] ),
    .Y(_03918_));
 sky130_fd_sc_hd__xnor2_2 _16573_ (.A(_03917_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__a22o_2 _16574_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[12][31] ),
    .B1(_11712_),
    .B2(_03919_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _16575_ (.A0(\systolic_inst.A_outs[11][0] ),
    .A1(\systolic_inst.A_outs[10][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _16576_ (.A0(\systolic_inst.A_outs[11][1] ),
    .A1(\systolic_inst.A_outs[10][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _16577_ (.A0(\systolic_inst.A_outs[11][2] ),
    .A1(\systolic_inst.A_outs[10][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _16578_ (.A0(\systolic_inst.A_outs[11][3] ),
    .A1(\systolic_inst.A_outs[10][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _16579_ (.A0(\systolic_inst.A_outs[11][4] ),
    .A1(\systolic_inst.A_outs[10][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _16580_ (.A0(\systolic_inst.A_outs[11][5] ),
    .A1(\systolic_inst.A_outs[10][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _16581_ (.A0(\systolic_inst.A_outs[11][6] ),
    .A1(\systolic_inst.A_outs[10][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _16582_ (.A0(\systolic_inst.A_outs[11][7] ),
    .A1(\systolic_inst.A_outs[10][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _16583_ (.A0(\systolic_inst.B_outs[10][0] ),
    .A1(\systolic_inst.B_outs[6][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _16584_ (.A0(\systolic_inst.B_outs[10][1] ),
    .A1(\systolic_inst.B_outs[6][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _16585_ (.A0(\systolic_inst.B_outs[10][2] ),
    .A1(\systolic_inst.B_outs[6][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _16586_ (.A0(\systolic_inst.B_outs[10][3] ),
    .A1(\systolic_inst.B_outs[6][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _16587_ (.A0(\systolic_inst.B_outs[10][4] ),
    .A1(\systolic_inst.B_outs[6][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _16588_ (.A0(\systolic_inst.B_outs[10][5] ),
    .A1(\systolic_inst.B_outs[6][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _16589_ (.A0(\systolic_inst.B_outs[10][6] ),
    .A1(\systolic_inst.B_outs[6][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _16590_ (.A0(\systolic_inst.B_outs[10][7] ),
    .A1(\systolic_inst.B_outs[6][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01217_));
 sky130_fd_sc_hd__and3_2 _16591_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[11][0] ),
    .C(\systolic_inst.A_outs[11][0] ),
    .X(_03920_));
 sky130_fd_sc_hd__a21o_2 _16592_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[0] ),
    .B1(_03920_),
    .X(_01218_));
 sky130_fd_sc_hd__and4_2 _16593_ (.A(\systolic_inst.B_outs[11][0] ),
    .B(\systolic_inst.A_outs[11][0] ),
    .C(\systolic_inst.B_outs[11][1] ),
    .D(\systolic_inst.A_outs[11][1] ),
    .X(_03921_));
 sky130_fd_sc_hd__a22o_2 _16594_ (.A1(\systolic_inst.A_outs[11][0] ),
    .A2(\systolic_inst.B_outs[11][1] ),
    .B1(\systolic_inst.A_outs[11][1] ),
    .B2(\systolic_inst.B_outs[11][0] ),
    .X(_03922_));
 sky130_fd_sc_hd__nand2_2 _16595_ (.A(\systolic_inst.ce_local ),
    .B(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__a2bb2o_2 _16596_ (.A1_N(_03923_),
    .A2_N(_03921_),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01219_));
 sky130_fd_sc_hd__and2_2 _16597_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[2] ),
    .X(_03924_));
 sky130_fd_sc_hd__a22oi_2 _16598_ (.A1(\systolic_inst.B_outs[11][1] ),
    .A2(\systolic_inst.A_outs[11][1] ),
    .B1(\systolic_inst.A_outs[11][2] ),
    .B2(\systolic_inst.B_outs[11][0] ),
    .Y(_03925_));
 sky130_fd_sc_hd__and4_2 _16599_ (.A(\systolic_inst.B_outs[11][0] ),
    .B(\systolic_inst.B_outs[11][1] ),
    .C(\systolic_inst.A_outs[11][1] ),
    .D(\systolic_inst.A_outs[11][2] ),
    .X(_03926_));
 sky130_fd_sc_hd__or2_2 _16600_ (.A(_03925_),
    .B(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__or3b_2 _16601_ (.A(_03925_),
    .B(_03926_),
    .C_N(_03921_),
    .X(_03928_));
 sky130_fd_sc_hd__xnor2_2 _16602_ (.A(_03921_),
    .B(_03927_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand3_2 _16603_ (.A(\systolic_inst.A_outs[11][0] ),
    .B(\systolic_inst.B_outs[11][2] ),
    .C(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__a21o_2 _16604_ (.A1(\systolic_inst.A_outs[11][0] ),
    .A2(\systolic_inst.B_outs[11][2] ),
    .B1(_03929_),
    .X(_03931_));
 sky130_fd_sc_hd__a31o_2 _16605_ (.A1(\systolic_inst.ce_local ),
    .A2(_03930_),
    .A3(_03931_),
    .B1(_03924_),
    .X(_01220_));
 sky130_fd_sc_hd__a22oi_2 _16606_ (.A1(\systolic_inst.A_outs[11][1] ),
    .A2(\systolic_inst.B_outs[11][2] ),
    .B1(\systolic_inst.B_outs[11][3] ),
    .B2(\systolic_inst.A_outs[11][0] ),
    .Y(_03932_));
 sky130_fd_sc_hd__and4_2 _16607_ (.A(\systolic_inst.A_outs[11][0] ),
    .B(\systolic_inst.A_outs[11][1] ),
    .C(\systolic_inst.B_outs[11][2] ),
    .D(\systolic_inst.B_outs[11][3] ),
    .X(_03933_));
 sky130_fd_sc_hd__nor2_2 _16608_ (.A(_03932_),
    .B(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand4_2 _16609_ (.A(\systolic_inst.B_outs[11][0] ),
    .B(\systolic_inst.B_outs[11][1] ),
    .C(\systolic_inst.A_outs[11][2] ),
    .D(\systolic_inst.A_outs[11][3] ),
    .Y(_03935_));
 sky130_fd_sc_hd__a22o_2 _16610_ (.A1(\systolic_inst.B_outs[11][1] ),
    .A2(\systolic_inst.A_outs[11][2] ),
    .B1(\systolic_inst.A_outs[11][3] ),
    .B2(\systolic_inst.B_outs[11][0] ),
    .X(_03936_));
 sky130_fd_sc_hd__nand3_2 _16611_ (.A(_03926_),
    .B(_03935_),
    .C(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__a21o_2 _16612_ (.A1(_03935_),
    .A2(_03936_),
    .B1(_03926_),
    .X(_03938_));
 sky130_fd_sc_hd__and2_2 _16613_ (.A(_03937_),
    .B(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__nand2_2 _16614_ (.A(_03934_),
    .B(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__xnor2_2 _16615_ (.A(_03934_),
    .B(_03939_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21oi_2 _16616_ (.A1(_03928_),
    .A2(_03930_),
    .B1(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__a31o_2 _16617_ (.A1(_03928_),
    .A2(_03930_),
    .A3(_03941_),
    .B1(_11258_),
    .X(_03943_));
 sky130_fd_sc_hd__a2bb2o_2 _16618_ (.A1_N(_03943_),
    .A2_N(_03942_),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[3] ),
    .B2(_11258_),
    .X(_01221_));
 sky130_fd_sc_hd__and2_2 _16619_ (.A(\systolic_inst.B_outs[11][2] ),
    .B(\systolic_inst.A_outs[11][2] ),
    .X(_03944_));
 sky130_fd_sc_hd__nand4_2 _16620_ (.A(\systolic_inst.A_outs[11][0] ),
    .B(\systolic_inst.A_outs[11][1] ),
    .C(\systolic_inst.B_outs[11][3] ),
    .D(\systolic_inst.B_outs[11][4] ),
    .Y(_03945_));
 sky130_fd_sc_hd__a22o_2 _16621_ (.A1(\systolic_inst.A_outs[11][1] ),
    .A2(\systolic_inst.B_outs[11][3] ),
    .B1(\systolic_inst.B_outs[11][4] ),
    .B2(\systolic_inst.A_outs[11][0] ),
    .X(_03946_));
 sky130_fd_sc_hd__nand2_2 _16622_ (.A(_03945_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__xnor2_2 _16623_ (.A(_03944_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__a22o_2 _16624_ (.A1(\systolic_inst.B_outs[11][1] ),
    .A2(\systolic_inst.A_outs[11][3] ),
    .B1(\systolic_inst.A_outs[11][4] ),
    .B2(\systolic_inst.B_outs[11][0] ),
    .X(_03949_));
 sky130_fd_sc_hd__and3_2 _16625_ (.A(\systolic_inst.B_outs[11][0] ),
    .B(\systolic_inst.B_outs[11][1] ),
    .C(\systolic_inst.A_outs[11][3] ),
    .X(_03950_));
 sky130_fd_sc_hd__nand2_2 _16626_ (.A(\systolic_inst.A_outs[11][4] ),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__and3_2 _16627_ (.A(_03933_),
    .B(_03949_),
    .C(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__a21oi_2 _16628_ (.A1(_03949_),
    .A2(_03951_),
    .B1(_03933_),
    .Y(_03953_));
 sky130_fd_sc_hd__o21ai_2 _16629_ (.A1(_03952_),
    .A2(_03953_),
    .B1(_03935_),
    .Y(_03954_));
 sky130_fd_sc_hd__or3_2 _16630_ (.A(_03935_),
    .B(_03952_),
    .C(_03953_),
    .X(_03955_));
 sky130_fd_sc_hd__and3_2 _16631_ (.A(_03948_),
    .B(_03954_),
    .C(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__a21oi_2 _16632_ (.A1(_03954_),
    .A2(_03955_),
    .B1(_03948_),
    .Y(_03957_));
 sky130_fd_sc_hd__a211o_2 _16633_ (.A1(_03937_),
    .A2(_03940_),
    .B1(_03956_),
    .C1(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__o211ai_2 _16634_ (.A1(_03956_),
    .A2(_03957_),
    .B1(_03937_),
    .C1(_03940_),
    .Y(_03959_));
 sky130_fd_sc_hd__a21oi_2 _16635_ (.A1(_03958_),
    .A2(_03959_),
    .B1(_03942_),
    .Y(_03960_));
 sky130_fd_sc_hd__and3_2 _16636_ (.A(_03942_),
    .B(_03958_),
    .C(_03959_),
    .X(_03961_));
 sky130_fd_sc_hd__or3_2 _16637_ (.A(_11258_),
    .B(_03960_),
    .C(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__a21bo_2 _16638_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[4] ),
    .B1_N(_03962_),
    .X(_01222_));
 sky130_fd_sc_hd__and2b_2 _16639_ (.A_N(_03952_),
    .B(_03955_),
    .X(_03963_));
 sky130_fd_sc_hd__a21bo_2 _16640_ (.A1(_03944_),
    .A2(_03946_),
    .B1_N(_03945_),
    .X(_03964_));
 sky130_fd_sc_hd__a22oi_2 _16641_ (.A1(\systolic_inst.B_outs[11][1] ),
    .A2(\systolic_inst.A_outs[11][4] ),
    .B1(\systolic_inst.A_outs[11][5] ),
    .B2(\systolic_inst.B_outs[11][0] ),
    .Y(_03965_));
 sky130_fd_sc_hd__and4_2 _16642_ (.A(\systolic_inst.B_outs[11][0] ),
    .B(\systolic_inst.B_outs[11][1] ),
    .C(\systolic_inst.A_outs[11][4] ),
    .D(\systolic_inst.A_outs[11][5] ),
    .X(_03966_));
 sky130_fd_sc_hd__nor2_2 _16643_ (.A(_03965_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__xor2_2 _16644_ (.A(_03964_),
    .B(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__xor2_2 _16645_ (.A(_03951_),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__and4_2 _16646_ (.A(\systolic_inst.A_outs[11][1] ),
    .B(\systolic_inst.A_outs[11][2] ),
    .C(\systolic_inst.B_outs[11][3] ),
    .D(\systolic_inst.B_outs[11][4] ),
    .X(_03970_));
 sky130_fd_sc_hd__a22oi_2 _16647_ (.A1(\systolic_inst.A_outs[11][2] ),
    .A2(\systolic_inst.B_outs[11][3] ),
    .B1(\systolic_inst.B_outs[11][4] ),
    .B2(\systolic_inst.A_outs[11][1] ),
    .Y(_03971_));
 sky130_fd_sc_hd__a22o_2 _16648_ (.A1(\systolic_inst.A_outs[11][2] ),
    .A2(\systolic_inst.B_outs[11][3] ),
    .B1(\systolic_inst.B_outs[11][4] ),
    .B2(\systolic_inst.A_outs[11][1] ),
    .X(_03972_));
 sky130_fd_sc_hd__and4b_2 _16649_ (.A_N(_03970_),
    .B(_03972_),
    .C(\systolic_inst.B_outs[11][2] ),
    .D(\systolic_inst.A_outs[11][3] ),
    .X(_03973_));
 sky130_fd_sc_hd__o2bb2a_2 _16650_ (.A1_N(\systolic_inst.B_outs[11][2] ),
    .A2_N(\systolic_inst.A_outs[11][3] ),
    .B1(_03970_),
    .B2(_03971_),
    .X(_03974_));
 sky130_fd_sc_hd__and4bb_2 _16651_ (.A_N(_03973_),
    .B_N(_03974_),
    .C(\systolic_inst.A_outs[11][0] ),
    .D(\systolic_inst.B_outs[11][5] ),
    .X(_03975_));
 sky130_fd_sc_hd__o2bb2a_2 _16652_ (.A1_N(\systolic_inst.A_outs[11][0] ),
    .A2_N(\systolic_inst.B_outs[11][5] ),
    .B1(_03973_),
    .B2(_03974_),
    .X(_03976_));
 sky130_fd_sc_hd__or2_2 _16653_ (.A(_03975_),
    .B(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__nor2_2 _16654_ (.A(_03969_),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__xor2_2 _16655_ (.A(_03969_),
    .B(_03977_),
    .X(_03979_));
 sky130_fd_sc_hd__nand2_2 _16656_ (.A(_03956_),
    .B(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__xor2_2 _16657_ (.A(_03956_),
    .B(_03979_),
    .X(_03981_));
 sky130_fd_sc_hd__nand2b_2 _16658_ (.A_N(_03963_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__xnor2_2 _16659_ (.A(_03963_),
    .B(_03981_),
    .Y(_03983_));
 sky130_fd_sc_hd__a21bo_2 _16660_ (.A1(_03942_),
    .A2(_03959_),
    .B1_N(_03958_),
    .X(_03984_));
 sky130_fd_sc_hd__nand2_2 _16661_ (.A(_03983_),
    .B(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__o21a_2 _16662_ (.A1(_03983_),
    .A2(_03984_),
    .B1(\systolic_inst.ce_local ),
    .X(_03986_));
 sky130_fd_sc_hd__a22o_2 _16663_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[5] ),
    .B1(_03985_),
    .B2(_03986_),
    .X(_01223_));
 sky130_fd_sc_hd__a32o_2 _16664_ (.A1(\systolic_inst.A_outs[11][4] ),
    .A2(_03950_),
    .A3(_03968_),
    .B1(_03967_),
    .B2(_03964_),
    .X(_03987_));
 sky130_fd_sc_hd__a31o_2 _16665_ (.A1(\systolic_inst.B_outs[11][2] ),
    .A2(\systolic_inst.A_outs[11][3] ),
    .A3(_03972_),
    .B1(_03970_),
    .X(_03988_));
 sky130_fd_sc_hd__a22oi_2 _16666_ (.A1(\systolic_inst.B_outs[11][1] ),
    .A2(\systolic_inst.A_outs[11][5] ),
    .B1(\systolic_inst.A_outs[11][6] ),
    .B2(\systolic_inst.B_outs[11][0] ),
    .Y(_03989_));
 sky130_fd_sc_hd__and4_2 _16667_ (.A(\systolic_inst.B_outs[11][0] ),
    .B(\systolic_inst.B_outs[11][1] ),
    .C(\systolic_inst.A_outs[11][5] ),
    .D(\systolic_inst.A_outs[11][6] ),
    .X(_03990_));
 sky130_fd_sc_hd__or2_2 _16668_ (.A(_03989_),
    .B(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__and2b_2 _16669_ (.A_N(_03991_),
    .B(_03988_),
    .X(_03992_));
 sky130_fd_sc_hd__xnor2_2 _16670_ (.A(_03988_),
    .B(_03991_),
    .Y(_03993_));
 sky130_fd_sc_hd__xor2_2 _16671_ (.A(_03966_),
    .B(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__nand4_2 _16672_ (.A(\systolic_inst.A_outs[11][2] ),
    .B(\systolic_inst.B_outs[11][3] ),
    .C(\systolic_inst.A_outs[11][3] ),
    .D(\systolic_inst.B_outs[11][4] ),
    .Y(_03995_));
 sky130_fd_sc_hd__a22o_2 _16673_ (.A1(\systolic_inst.B_outs[11][3] ),
    .A2(\systolic_inst.A_outs[11][3] ),
    .B1(\systolic_inst.B_outs[11][4] ),
    .B2(\systolic_inst.A_outs[11][2] ),
    .X(_03996_));
 sky130_fd_sc_hd__nand4_2 _16674_ (.A(\systolic_inst.B_outs[11][2] ),
    .B(\systolic_inst.A_outs[11][4] ),
    .C(_03995_),
    .D(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__a22o_2 _16675_ (.A1(\systolic_inst.B_outs[11][2] ),
    .A2(\systolic_inst.A_outs[11][4] ),
    .B1(_03995_),
    .B2(_03996_),
    .X(_03998_));
 sky130_fd_sc_hd__a22oi_2 _16676_ (.A1(\systolic_inst.A_outs[11][1] ),
    .A2(\systolic_inst.B_outs[11][5] ),
    .B1(\systolic_inst.B_outs[11][6] ),
    .B2(\systolic_inst.A_outs[11][0] ),
    .Y(_03999_));
 sky130_fd_sc_hd__nand2_2 _16677_ (.A(\systolic_inst.A_outs[11][1] ),
    .B(\systolic_inst.B_outs[11][6] ),
    .Y(_04000_));
 sky130_fd_sc_hd__and4_2 _16678_ (.A(\systolic_inst.A_outs[11][0] ),
    .B(\systolic_inst.A_outs[11][1] ),
    .C(\systolic_inst.B_outs[11][5] ),
    .D(\systolic_inst.B_outs[11][6] ),
    .X(_04001_));
 sky130_fd_sc_hd__nor2_2 _16679_ (.A(_03999_),
    .B(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__nand3_2 _16680_ (.A(_03997_),
    .B(_03998_),
    .C(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__a21o_2 _16681_ (.A1(_03997_),
    .A2(_03998_),
    .B1(_04002_),
    .X(_04004_));
 sky130_fd_sc_hd__and3_2 _16682_ (.A(_03975_),
    .B(_04003_),
    .C(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__a21oi_2 _16683_ (.A1(_04003_),
    .A2(_04004_),
    .B1(_03975_),
    .Y(_04006_));
 sky130_fd_sc_hd__or3b_2 _16684_ (.A(_04005_),
    .B(_04006_),
    .C_N(_03994_),
    .X(_04007_));
 sky130_fd_sc_hd__o21bai_2 _16685_ (.A1(_04005_),
    .A2(_04006_),
    .B1_N(_03994_),
    .Y(_04008_));
 sky130_fd_sc_hd__nand3_2 _16686_ (.A(_03978_),
    .B(_04007_),
    .C(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__a21o_2 _16687_ (.A1(_04007_),
    .A2(_04008_),
    .B1(_03978_),
    .X(_04010_));
 sky130_fd_sc_hd__and3_2 _16688_ (.A(_03987_),
    .B(_04009_),
    .C(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__a21oi_2 _16689_ (.A1(_04009_),
    .A2(_04010_),
    .B1(_03987_),
    .Y(_04012_));
 sky130_fd_sc_hd__a211oi_2 _16690_ (.A1(_03980_),
    .A2(_03982_),
    .B1(_04011_),
    .C1(_04012_),
    .Y(_04013_));
 sky130_fd_sc_hd__o211a_2 _16691_ (.A1(_04011_),
    .A2(_04012_),
    .B1(_03980_),
    .C1(_03982_),
    .X(_04014_));
 sky130_fd_sc_hd__nor2_2 _16692_ (.A(_04013_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__xnor2_2 _16693_ (.A(_03985_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__mux2_1 _16694_ (.A0(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[6] ),
    .A1(_04016_),
    .S(\systolic_inst.ce_local ),
    .X(_01224_));
 sky130_fd_sc_hd__a21boi_2 _16695_ (.A1(_03987_),
    .A2(_04010_),
    .B1_N(_04009_),
    .Y(_04017_));
 sky130_fd_sc_hd__a21oi_2 _16696_ (.A1(_03966_),
    .A2(_03993_),
    .B1(_03992_),
    .Y(_04018_));
 sky130_fd_sc_hd__nand2_2 _16697_ (.A(_03995_),
    .B(_03997_),
    .Y(_04019_));
 sky130_fd_sc_hd__a22o_2 _16698_ (.A1(\systolic_inst.B_outs[11][1] ),
    .A2(\systolic_inst.A_outs[11][6] ),
    .B1(\systolic_inst.A_outs[11][7] ),
    .B2(\systolic_inst.B_outs[11][0] ),
    .X(_04020_));
 sky130_fd_sc_hd__nand4_2 _16699_ (.A(\systolic_inst.B_outs[11][0] ),
    .B(\systolic_inst.B_outs[11][1] ),
    .C(\systolic_inst.A_outs[11][6] ),
    .D(\systolic_inst.A_outs[11][7] ),
    .Y(_04021_));
 sky130_fd_sc_hd__nand2_2 _16700_ (.A(_04020_),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__xnor2_2 _16701_ (.A(_11262_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand2b_2 _16702_ (.A_N(_04023_),
    .B(_04019_),
    .Y(_04024_));
 sky130_fd_sc_hd__xnor2_2 _16703_ (.A(_04019_),
    .B(_04023_),
    .Y(_04025_));
 sky130_fd_sc_hd__xnor2_2 _16704_ (.A(_03990_),
    .B(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__nand2_2 _16705_ (.A(\systolic_inst.B_outs[11][2] ),
    .B(\systolic_inst.A_outs[11][5] ),
    .Y(_04027_));
 sky130_fd_sc_hd__and4_2 _16706_ (.A(\systolic_inst.B_outs[11][3] ),
    .B(\systolic_inst.A_outs[11][3] ),
    .C(\systolic_inst.B_outs[11][4] ),
    .D(\systolic_inst.A_outs[11][4] ),
    .X(_04028_));
 sky130_fd_sc_hd__a22oi_2 _16707_ (.A1(\systolic_inst.A_outs[11][3] ),
    .A2(\systolic_inst.B_outs[11][4] ),
    .B1(\systolic_inst.A_outs[11][4] ),
    .B2(\systolic_inst.B_outs[11][3] ),
    .Y(_04029_));
 sky130_fd_sc_hd__or2_2 _16708_ (.A(_04028_),
    .B(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__xnor2_2 _16709_ (.A(_04027_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__nand2_2 _16710_ (.A(\systolic_inst.A_outs[11][2] ),
    .B(\systolic_inst.B_outs[11][5] ),
    .Y(_04032_));
 sky130_fd_sc_hd__and2b_2 _16711_ (.A_N(\systolic_inst.A_outs[11][0] ),
    .B(\systolic_inst.B_outs[11][7] ),
    .X(_04033_));
 sky130_fd_sc_hd__and3_2 _16712_ (.A(\systolic_inst.A_outs[11][1] ),
    .B(\systolic_inst.B_outs[11][6] ),
    .C(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__xnor2_2 _16713_ (.A(_04000_),
    .B(_04033_),
    .Y(_04035_));
 sky130_fd_sc_hd__xnor2_2 _16714_ (.A(_04032_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__xnor2_2 _16715_ (.A(_04001_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__nor2_2 _16716_ (.A(_04031_),
    .B(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__xnor2_2 _16717_ (.A(_04031_),
    .B(_04037_),
    .Y(_04039_));
 sky130_fd_sc_hd__or2_2 _16718_ (.A(_04003_),
    .B(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__and2_2 _16719_ (.A(_04003_),
    .B(_04039_),
    .X(_04041_));
 sky130_fd_sc_hd__xor2_2 _16720_ (.A(_04003_),
    .B(_04039_),
    .X(_04042_));
 sky130_fd_sc_hd__xnor2_2 _16721_ (.A(_04026_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__and2b_2 _16722_ (.A_N(_04005_),
    .B(_04007_),
    .X(_04044_));
 sky130_fd_sc_hd__nand2b_2 _16723_ (.A_N(_04044_),
    .B(_04043_),
    .Y(_04045_));
 sky130_fd_sc_hd__xnor2_2 _16724_ (.A(_04043_),
    .B(_04044_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2b_2 _16725_ (.A_N(_04018_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__xnor2_2 _16726_ (.A(_04018_),
    .B(_04046_),
    .Y(_04048_));
 sky130_fd_sc_hd__and2b_2 _16727_ (.A_N(_04017_),
    .B(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__xnor2_2 _16728_ (.A(_04017_),
    .B(_04048_),
    .Y(_04050_));
 sky130_fd_sc_hd__a31o_2 _16729_ (.A1(_03983_),
    .A2(_03984_),
    .A3(_04015_),
    .B1(_04013_),
    .X(_04051_));
 sky130_fd_sc_hd__xor2_2 _16730_ (.A(_04050_),
    .B(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__mux2_1 _16731_ (.A0(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[7] ),
    .A1(_04052_),
    .S(\systolic_inst.ce_local ),
    .X(_01225_));
 sky130_fd_sc_hd__a21bo_2 _16732_ (.A1(_03990_),
    .A2(_04025_),
    .B1_N(_04024_),
    .X(_04053_));
 sky130_fd_sc_hd__a21bo_2 _16733_ (.A1(\systolic_inst.B_outs[11][7] ),
    .A2(_04020_),
    .B1_N(_04021_),
    .X(_04054_));
 sky130_fd_sc_hd__o21bai_2 _16734_ (.A1(_04027_),
    .A2(_04029_),
    .B1_N(_04028_),
    .Y(_04055_));
 sky130_fd_sc_hd__o21a_2 _16735_ (.A1(\systolic_inst.B_outs[11][0] ),
    .A2(\systolic_inst.B_outs[11][1] ),
    .B1(\systolic_inst.A_outs[11][7] ),
    .X(_04056_));
 sky130_fd_sc_hd__o21ai_2 _16736_ (.A1(\systolic_inst.B_outs[11][0] ),
    .A2(\systolic_inst.B_outs[11][1] ),
    .B1(\systolic_inst.A_outs[11][7] ),
    .Y(_04057_));
 sky130_fd_sc_hd__a21o_2 _16737_ (.A1(\systolic_inst.B_outs[11][0] ),
    .A2(\systolic_inst.B_outs[11][1] ),
    .B1(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__and2b_2 _16738_ (.A_N(_04058_),
    .B(_04055_),
    .X(_04059_));
 sky130_fd_sc_hd__xnor2_2 _16739_ (.A(_04055_),
    .B(_04058_),
    .Y(_04060_));
 sky130_fd_sc_hd__xnor2_2 _16740_ (.A(_04054_),
    .B(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__and4_2 _16741_ (.A(\systolic_inst.B_outs[11][3] ),
    .B(\systolic_inst.B_outs[11][4] ),
    .C(\systolic_inst.A_outs[11][4] ),
    .D(\systolic_inst.A_outs[11][5] ),
    .X(_04062_));
 sky130_fd_sc_hd__a22oi_2 _16742_ (.A1(\systolic_inst.B_outs[11][4] ),
    .A2(\systolic_inst.A_outs[11][4] ),
    .B1(\systolic_inst.A_outs[11][5] ),
    .B2(\systolic_inst.B_outs[11][3] ),
    .Y(_04063_));
 sky130_fd_sc_hd__nor2_2 _16743_ (.A(_04062_),
    .B(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__nand2_2 _16744_ (.A(\systolic_inst.B_outs[11][2] ),
    .B(\systolic_inst.A_outs[11][6] ),
    .Y(_04065_));
 sky130_fd_sc_hd__xnor2_2 _16745_ (.A(_04064_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__nand2_2 _16746_ (.A(\systolic_inst.A_outs[11][3] ),
    .B(\systolic_inst.B_outs[11][5] ),
    .Y(_04067_));
 sky130_fd_sc_hd__and4b_2 _16747_ (.A_N(\systolic_inst.A_outs[11][1] ),
    .B(\systolic_inst.A_outs[11][2] ),
    .C(\systolic_inst.B_outs[11][6] ),
    .D(\systolic_inst.B_outs[11][7] ),
    .X(_04068_));
 sky130_fd_sc_hd__a2bb2o_2 _16748_ (.A1_N(\systolic_inst.A_outs[11][1] ),
    .A2_N(_11262_),
    .B1(\systolic_inst.B_outs[11][6] ),
    .B2(\systolic_inst.A_outs[11][2] ),
    .X(_04069_));
 sky130_fd_sc_hd__and2b_2 _16749_ (.A_N(_04068_),
    .B(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__xnor2_2 _16750_ (.A(_04067_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__a31o_2 _16751_ (.A1(\systolic_inst.A_outs[11][2] ),
    .A2(\systolic_inst.B_outs[11][5] ),
    .A3(_04035_),
    .B1(_04034_),
    .X(_04072_));
 sky130_fd_sc_hd__and2_2 _16752_ (.A(_04071_),
    .B(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__xor2_2 _16753_ (.A(_04071_),
    .B(_04072_),
    .X(_04074_));
 sky130_fd_sc_hd__xor2_2 _16754_ (.A(_04066_),
    .B(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__a21oi_2 _16755_ (.A1(_04001_),
    .A2(_04036_),
    .B1(_04038_),
    .Y(_04076_));
 sky130_fd_sc_hd__and2b_2 _16756_ (.A_N(_04076_),
    .B(_04075_),
    .X(_04077_));
 sky130_fd_sc_hd__xor2_2 _16757_ (.A(_04075_),
    .B(_04076_),
    .X(_04078_));
 sky130_fd_sc_hd__xor2_2 _16758_ (.A(_04061_),
    .B(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__o21a_2 _16759_ (.A1(_04026_),
    .A2(_04041_),
    .B1(_04040_),
    .X(_04080_));
 sky130_fd_sc_hd__nand2b_2 _16760_ (.A_N(_04080_),
    .B(_04079_),
    .Y(_04081_));
 sky130_fd_sc_hd__xor2_2 _16761_ (.A(_04079_),
    .B(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__nand2b_2 _16762_ (.A_N(_04082_),
    .B(_04053_),
    .Y(_04083_));
 sky130_fd_sc_hd__xor2_2 _16763_ (.A(_04053_),
    .B(_04082_),
    .X(_04084_));
 sky130_fd_sc_hd__and2_2 _16764_ (.A(_04045_),
    .B(_04047_),
    .X(_04085_));
 sky130_fd_sc_hd__or2_2 _16765_ (.A(_04084_),
    .B(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__xor2_2 _16766_ (.A(_04084_),
    .B(_04085_),
    .X(_04087_));
 sky130_fd_sc_hd__a21o_2 _16767_ (.A1(_04050_),
    .A2(_04051_),
    .B1(_04049_),
    .X(_04088_));
 sky130_fd_sc_hd__nand2_2 _16768_ (.A(_04087_),
    .B(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__or2_2 _16769_ (.A(_04087_),
    .B(_04088_),
    .X(_04090_));
 sky130_fd_sc_hd__and2_2 _16770_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[8] ),
    .X(_04091_));
 sky130_fd_sc_hd__a31o_2 _16771_ (.A1(\systolic_inst.ce_local ),
    .A2(_04089_),
    .A3(_04090_),
    .B1(_04091_),
    .X(_01226_));
 sky130_fd_sc_hd__a21o_2 _16772_ (.A1(_04054_),
    .A2(_04060_),
    .B1(_04059_),
    .X(_04092_));
 sky130_fd_sc_hd__o21ba_2 _16773_ (.A1(_04063_),
    .A2(_04065_),
    .B1_N(_04062_),
    .X(_04093_));
 sky130_fd_sc_hd__nor2_2 _16774_ (.A(_04057_),
    .B(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__and2_2 _16775_ (.A(_04057_),
    .B(_04093_),
    .X(_04095_));
 sky130_fd_sc_hd__or2_2 _16776_ (.A(_04094_),
    .B(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__nand2_2 _16777_ (.A(\systolic_inst.B_outs[11][2] ),
    .B(\systolic_inst.A_outs[11][7] ),
    .Y(_04097_));
 sky130_fd_sc_hd__a22oi_2 _16778_ (.A1(\systolic_inst.B_outs[11][4] ),
    .A2(\systolic_inst.A_outs[11][5] ),
    .B1(\systolic_inst.A_outs[11][6] ),
    .B2(\systolic_inst.B_outs[11][3] ),
    .Y(_04098_));
 sky130_fd_sc_hd__and4_2 _16779_ (.A(\systolic_inst.B_outs[11][3] ),
    .B(\systolic_inst.B_outs[11][4] ),
    .C(\systolic_inst.A_outs[11][5] ),
    .D(\systolic_inst.A_outs[11][6] ),
    .X(_04099_));
 sky130_fd_sc_hd__nor2_2 _16780_ (.A(_04098_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__xnor2_2 _16781_ (.A(_04097_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_2 _16782_ (.A(\systolic_inst.A_outs[11][4] ),
    .B(\systolic_inst.B_outs[11][5] ),
    .Y(_04102_));
 sky130_fd_sc_hd__and4b_2 _16783_ (.A_N(\systolic_inst.A_outs[11][2] ),
    .B(\systolic_inst.A_outs[11][3] ),
    .C(\systolic_inst.B_outs[11][6] ),
    .D(\systolic_inst.B_outs[11][7] ),
    .X(_04103_));
 sky130_fd_sc_hd__o2bb2a_2 _16784_ (.A1_N(\systolic_inst.A_outs[11][3] ),
    .A2_N(\systolic_inst.B_outs[11][6] ),
    .B1(_11262_),
    .B2(\systolic_inst.A_outs[11][2] ),
    .X(_04104_));
 sky130_fd_sc_hd__nor2_2 _16785_ (.A(_04103_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__xnor2_2 _16786_ (.A(_04102_),
    .B(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__a31oi_2 _16787_ (.A1(\systolic_inst.A_outs[11][3] ),
    .A2(\systolic_inst.B_outs[11][5] ),
    .A3(_04069_),
    .B1(_04068_),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2b_2 _16788_ (.A_N(_04107_),
    .B(_04106_),
    .Y(_04108_));
 sky130_fd_sc_hd__xnor2_2 _16789_ (.A(_04106_),
    .B(_04107_),
    .Y(_04109_));
 sky130_fd_sc_hd__nand2_2 _16790_ (.A(_04101_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__or2_2 _16791_ (.A(_04101_),
    .B(_04109_),
    .X(_04111_));
 sky130_fd_sc_hd__nand2_2 _16792_ (.A(_04110_),
    .B(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__a21o_2 _16793_ (.A1(_04066_),
    .A2(_04074_),
    .B1(_04073_),
    .X(_04113_));
 sky130_fd_sc_hd__and2b_2 _16794_ (.A_N(_04112_),
    .B(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__xor2_2 _16795_ (.A(_04112_),
    .B(_04113_),
    .X(_04115_));
 sky130_fd_sc_hd__xor2_2 _16796_ (.A(_04096_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__o21ba_2 _16797_ (.A1(_04061_),
    .A2(_04078_),
    .B1_N(_04077_),
    .X(_04117_));
 sky130_fd_sc_hd__nand2b_2 _16798_ (.A_N(_04117_),
    .B(_04116_),
    .Y(_04118_));
 sky130_fd_sc_hd__xnor2_2 _16799_ (.A(_04116_),
    .B(_04117_),
    .Y(_04119_));
 sky130_fd_sc_hd__xnor2_2 _16800_ (.A(_04092_),
    .B(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__a21o_2 _16801_ (.A1(_04081_),
    .A2(_04083_),
    .B1(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__and3_2 _16802_ (.A(_04081_),
    .B(_04083_),
    .C(_04120_),
    .X(_04122_));
 sky130_fd_sc_hd__inv_2 _16803_ (.A(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__nand2_2 _16804_ (.A(_04121_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__a21o_2 _16805_ (.A1(_04086_),
    .A2(_04089_),
    .B1(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__a31oi_2 _16806_ (.A1(_04086_),
    .A2(_04089_),
    .A3(_04124_),
    .B1(_11258_),
    .Y(_04126_));
 sky130_fd_sc_hd__a22o_2 _16807_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[9] ),
    .B1(_04125_),
    .B2(_04126_),
    .X(_01227_));
 sky130_fd_sc_hd__o21ba_2 _16808_ (.A1(_04097_),
    .A2(_04098_),
    .B1_N(_04099_),
    .X(_04127_));
 sky130_fd_sc_hd__nor2_2 _16809_ (.A(_04057_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__and2_2 _16810_ (.A(_04057_),
    .B(_04127_),
    .X(_04129_));
 sky130_fd_sc_hd__or2_2 _16811_ (.A(_04128_),
    .B(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__a22o_2 _16812_ (.A1(\systolic_inst.B_outs[11][4] ),
    .A2(\systolic_inst.A_outs[11][6] ),
    .B1(\systolic_inst.A_outs[11][7] ),
    .B2(\systolic_inst.B_outs[11][3] ),
    .X(_04131_));
 sky130_fd_sc_hd__and3_2 _16813_ (.A(\systolic_inst.B_outs[11][3] ),
    .B(\systolic_inst.B_outs[11][4] ),
    .C(\systolic_inst.A_outs[11][7] ),
    .X(_04132_));
 sky130_fd_sc_hd__a21bo_2 _16814_ (.A1(\systolic_inst.A_outs[11][6] ),
    .A2(_04132_),
    .B1_N(_04131_),
    .X(_04133_));
 sky130_fd_sc_hd__xor2_2 _16815_ (.A(_04097_),
    .B(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__nand2_2 _16816_ (.A(\systolic_inst.B_outs[11][5] ),
    .B(\systolic_inst.A_outs[11][5] ),
    .Y(_04135_));
 sky130_fd_sc_hd__and4b_2 _16817_ (.A_N(\systolic_inst.A_outs[11][3] ),
    .B(\systolic_inst.A_outs[11][4] ),
    .C(\systolic_inst.B_outs[11][6] ),
    .D(\systolic_inst.B_outs[11][7] ),
    .X(_04136_));
 sky130_fd_sc_hd__o2bb2a_2 _16818_ (.A1_N(\systolic_inst.A_outs[11][4] ),
    .A2_N(\systolic_inst.B_outs[11][6] ),
    .B1(_11262_),
    .B2(\systolic_inst.A_outs[11][3] ),
    .X(_04137_));
 sky130_fd_sc_hd__nor2_2 _16819_ (.A(_04136_),
    .B(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__xnor2_2 _16820_ (.A(_04135_),
    .B(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__o21ba_2 _16821_ (.A1(_04102_),
    .A2(_04104_),
    .B1_N(_04103_),
    .X(_04140_));
 sky130_fd_sc_hd__nand2b_2 _16822_ (.A_N(_04140_),
    .B(_04139_),
    .Y(_04141_));
 sky130_fd_sc_hd__xnor2_2 _16823_ (.A(_04139_),
    .B(_04140_),
    .Y(_04142_));
 sky130_fd_sc_hd__nand2_2 _16824_ (.A(_04134_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__xnor2_2 _16825_ (.A(_04134_),
    .B(_04142_),
    .Y(_04144_));
 sky130_fd_sc_hd__a21o_2 _16826_ (.A1(_04108_),
    .A2(_04110_),
    .B1(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__nand3_2 _16827_ (.A(_04108_),
    .B(_04110_),
    .C(_04144_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_2 _16828_ (.A(_04145_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__xor2_2 _16829_ (.A(_04130_),
    .B(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__o21ba_2 _16830_ (.A1(_04096_),
    .A2(_04115_),
    .B1_N(_04114_),
    .X(_04149_));
 sky130_fd_sc_hd__nand2b_2 _16831_ (.A_N(_04149_),
    .B(_04148_),
    .Y(_04150_));
 sky130_fd_sc_hd__xnor2_2 _16832_ (.A(_04148_),
    .B(_04149_),
    .Y(_04151_));
 sky130_fd_sc_hd__nand2_2 _16833_ (.A(_04094_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__xnor2_2 _16834_ (.A(_04094_),
    .B(_04151_),
    .Y(_04153_));
 sky130_fd_sc_hd__a21boi_2 _16835_ (.A1(_04092_),
    .A2(_04119_),
    .B1_N(_04118_),
    .Y(_04154_));
 sky130_fd_sc_hd__nor2_2 _16836_ (.A(_04153_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__and2_2 _16837_ (.A(_04153_),
    .B(_04154_),
    .X(_04156_));
 sky130_fd_sc_hd__or2_2 _16838_ (.A(_04155_),
    .B(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__or3b_2 _16839_ (.A(_04122_),
    .B(_04089_),
    .C_N(_04121_),
    .X(_04158_));
 sky130_fd_sc_hd__a21o_2 _16840_ (.A1(_04086_),
    .A2(_04121_),
    .B1(_04122_),
    .X(_04159_));
 sky130_fd_sc_hd__and3_2 _16841_ (.A(_04157_),
    .B(_04158_),
    .C(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__a21oi_2 _16842_ (.A1(_04158_),
    .A2(_04159_),
    .B1(_04157_),
    .Y(_04161_));
 sky130_fd_sc_hd__or3_2 _16843_ (.A(_11258_),
    .B(_04160_),
    .C(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__a21bo_2 _16844_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[10] ),
    .B1_N(_04162_),
    .X(_01228_));
 sky130_fd_sc_hd__o2bb2a_2 _16845_ (.A1_N(\systolic_inst.A_outs[11][6] ),
    .A2_N(_04132_),
    .B1(_04133_),
    .B2(_04097_),
    .X(_04163_));
 sky130_fd_sc_hd__or2_2 _16846_ (.A(_04057_),
    .B(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__nand2_2 _16847_ (.A(_04057_),
    .B(_04163_),
    .Y(_04165_));
 sky130_fd_sc_hd__nand2_2 _16848_ (.A(_04164_),
    .B(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__or2_2 _16849_ (.A(\systolic_inst.B_outs[11][3] ),
    .B(\systolic_inst.B_outs[11][4] ),
    .X(_04167_));
 sky130_fd_sc_hd__and3b_2 _16850_ (.A_N(_04132_),
    .B(_04167_),
    .C(\systolic_inst.A_outs[11][7] ),
    .X(_04168_));
 sky130_fd_sc_hd__xnor2_2 _16851_ (.A(_04097_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__nand2_2 _16852_ (.A(\systolic_inst.B_outs[11][5] ),
    .B(\systolic_inst.A_outs[11][6] ),
    .Y(_04170_));
 sky130_fd_sc_hd__and4b_2 _16853_ (.A_N(\systolic_inst.A_outs[11][4] ),
    .B(\systolic_inst.A_outs[11][5] ),
    .C(\systolic_inst.B_outs[11][6] ),
    .D(\systolic_inst.B_outs[11][7] ),
    .X(_04171_));
 sky130_fd_sc_hd__o2bb2a_2 _16854_ (.A1_N(\systolic_inst.A_outs[11][5] ),
    .A2_N(\systolic_inst.B_outs[11][6] ),
    .B1(_11262_),
    .B2(\systolic_inst.A_outs[11][4] ),
    .X(_04172_));
 sky130_fd_sc_hd__or2_2 _16855_ (.A(_04171_),
    .B(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__xor2_2 _16856_ (.A(_04170_),
    .B(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__o21ba_2 _16857_ (.A1(_04135_),
    .A2(_04137_),
    .B1_N(_04136_),
    .X(_04175_));
 sky130_fd_sc_hd__nand2b_2 _16858_ (.A_N(_04175_),
    .B(_04174_),
    .Y(_04176_));
 sky130_fd_sc_hd__xnor2_2 _16859_ (.A(_04174_),
    .B(_04175_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_2 _16860_ (.A(_04169_),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__xnor2_2 _16861_ (.A(_04169_),
    .B(_04177_),
    .Y(_04179_));
 sky130_fd_sc_hd__a21o_2 _16862_ (.A1(_04141_),
    .A2(_04143_),
    .B1(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__nand3_2 _16863_ (.A(_04141_),
    .B(_04143_),
    .C(_04179_),
    .Y(_04181_));
 sky130_fd_sc_hd__nand2_2 _16864_ (.A(_04180_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__xor2_2 _16865_ (.A(_04166_),
    .B(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__o21a_2 _16866_ (.A1(_04130_),
    .A2(_04147_),
    .B1(_04145_),
    .X(_04184_));
 sky130_fd_sc_hd__and2b_2 _16867_ (.A_N(_04184_),
    .B(_04183_),
    .X(_04185_));
 sky130_fd_sc_hd__and2b_2 _16868_ (.A_N(_04183_),
    .B(_04184_),
    .X(_04186_));
 sky130_fd_sc_hd__nor2_2 _16869_ (.A(_04185_),
    .B(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__xnor2_2 _16870_ (.A(_04128_),
    .B(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand3_2 _16871_ (.A(_04150_),
    .B(_04152_),
    .C(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__inv_2 _16872_ (.A(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__a21oi_2 _16873_ (.A1(_04150_),
    .A2(_04152_),
    .B1(_04188_),
    .Y(_04191_));
 sky130_fd_sc_hd__nor2_2 _16874_ (.A(_04190_),
    .B(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__or3_2 _16875_ (.A(_04155_),
    .B(_04161_),
    .C(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__o21ai_2 _16876_ (.A1(_04155_),
    .A2(_04161_),
    .B1(_04192_),
    .Y(_04194_));
 sky130_fd_sc_hd__and2_2 _16877_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[11] ),
    .X(_04195_));
 sky130_fd_sc_hd__a31o_2 _16878_ (.A1(\systolic_inst.ce_local ),
    .A2(_04193_),
    .A3(_04194_),
    .B1(_04195_),
    .X(_01229_));
 sky130_fd_sc_hd__a31o_2 _16879_ (.A1(\systolic_inst.B_outs[11][2] ),
    .A2(\systolic_inst.A_outs[11][7] ),
    .A3(_04167_),
    .B1(_04132_),
    .X(_04196_));
 sky130_fd_sc_hd__or2_2 _16880_ (.A(_04056_),
    .B(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__nand2_2 _16881_ (.A(_04056_),
    .B(_04196_),
    .Y(_04198_));
 sky130_fd_sc_hd__nand2_2 _16882_ (.A(_04197_),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__inv_2 _16883_ (.A(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__o2bb2a_2 _16884_ (.A1_N(\systolic_inst.B_outs[11][6] ),
    .A2_N(\systolic_inst.A_outs[11][6] ),
    .B1(_11262_),
    .B2(\systolic_inst.A_outs[11][5] ),
    .X(_04201_));
 sky130_fd_sc_hd__and4b_2 _16885_ (.A_N(\systolic_inst.A_outs[11][5] ),
    .B(\systolic_inst.B_outs[11][6] ),
    .C(\systolic_inst.A_outs[11][6] ),
    .D(\systolic_inst.B_outs[11][7] ),
    .X(_04202_));
 sky130_fd_sc_hd__nor2_2 _16886_ (.A(_04201_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__nand2_2 _16887_ (.A(\systolic_inst.B_outs[11][5] ),
    .B(\systolic_inst.A_outs[11][7] ),
    .Y(_04204_));
 sky130_fd_sc_hd__xnor2_2 _16888_ (.A(_04203_),
    .B(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__o21ba_2 _16889_ (.A1(_04170_),
    .A2(_04172_),
    .B1_N(_04171_),
    .X(_04206_));
 sky130_fd_sc_hd__nand2b_2 _16890_ (.A_N(_04206_),
    .B(_04205_),
    .Y(_04207_));
 sky130_fd_sc_hd__xnor2_2 _16891_ (.A(_04205_),
    .B(_04206_),
    .Y(_04208_));
 sky130_fd_sc_hd__xnor2_2 _16892_ (.A(_04169_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__a21o_2 _16893_ (.A1(_04176_),
    .A2(_04178_),
    .B1(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__nand3_2 _16894_ (.A(_04176_),
    .B(_04178_),
    .C(_04209_),
    .Y(_04211_));
 sky130_fd_sc_hd__nand2_2 _16895_ (.A(_04210_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__xnor2_2 _16896_ (.A(_04200_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__o21a_2 _16897_ (.A1(_04166_),
    .A2(_04182_),
    .B1(_04180_),
    .X(_04214_));
 sky130_fd_sc_hd__and2b_2 _16898_ (.A_N(_04214_),
    .B(_04213_),
    .X(_04215_));
 sky130_fd_sc_hd__and2b_2 _16899_ (.A_N(_04213_),
    .B(_04214_),
    .X(_04216_));
 sky130_fd_sc_hd__nor2_2 _16900_ (.A(_04215_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__and2b_2 _16901_ (.A_N(_04164_),
    .B(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__xor2_2 _16902_ (.A(_04164_),
    .B(_04217_),
    .X(_04219_));
 sky130_fd_sc_hd__a21oi_2 _16903_ (.A1(_04128_),
    .A2(_04187_),
    .B1(_04185_),
    .Y(_04220_));
 sky130_fd_sc_hd__or2_2 _16904_ (.A(_04219_),
    .B(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__nand2_2 _16905_ (.A(_04219_),
    .B(_04220_),
    .Y(_04222_));
 sky130_fd_sc_hd__nand2_2 _16906_ (.A(_04221_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__inv_2 _16907_ (.A(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__o31a_2 _16908_ (.A1(_04155_),
    .A2(_04161_),
    .A3(_04191_),
    .B1(_04189_),
    .X(_04225_));
 sky130_fd_sc_hd__xnor2_2 _16909_ (.A(_04223_),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__mux2_1 _16910_ (.A0(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[12] ),
    .A1(_04226_),
    .S(\systolic_inst.ce_local ),
    .X(_01230_));
 sky130_fd_sc_hd__nand2_2 _16911_ (.A(\systolic_inst.B_outs[11][6] ),
    .B(\systolic_inst.A_outs[11][7] ),
    .Y(_04227_));
 sky130_fd_sc_hd__or2_2 _16912_ (.A(\systolic_inst.A_outs[11][6] ),
    .B(_11262_),
    .X(_04228_));
 sky130_fd_sc_hd__and2_2 _16913_ (.A(_04227_),
    .B(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__nor2_2 _16914_ (.A(_04227_),
    .B(_04228_),
    .Y(_04230_));
 sky130_fd_sc_hd__nor2_2 _16915_ (.A(_04229_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__xnor2_2 _16916_ (.A(_04204_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__o21ba_2 _16917_ (.A1(_04201_),
    .A2(_04204_),
    .B1_N(_04202_),
    .X(_04233_));
 sky130_fd_sc_hd__nand2b_2 _16918_ (.A_N(_04233_),
    .B(_04232_),
    .Y(_04234_));
 sky130_fd_sc_hd__xnor2_2 _16919_ (.A(_04232_),
    .B(_04233_),
    .Y(_04235_));
 sky130_fd_sc_hd__nand2_2 _16920_ (.A(_04169_),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__or2_2 _16921_ (.A(_04169_),
    .B(_04235_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_2 _16922_ (.A(_04236_),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__a21bo_2 _16923_ (.A1(_04169_),
    .A2(_04208_),
    .B1_N(_04207_),
    .X(_04239_));
 sky130_fd_sc_hd__nand2b_2 _16924_ (.A_N(_04238_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__xor2_2 _16925_ (.A(_04238_),
    .B(_04239_),
    .X(_04241_));
 sky130_fd_sc_hd__xnor2_2 _16926_ (.A(_04200_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__o21a_2 _16927_ (.A1(_04199_),
    .A2(_04212_),
    .B1(_04210_),
    .X(_04243_));
 sky130_fd_sc_hd__and2b_2 _16928_ (.A_N(_04243_),
    .B(_04242_),
    .X(_04244_));
 sky130_fd_sc_hd__and2b_2 _16929_ (.A_N(_04242_),
    .B(_04243_),
    .X(_04245_));
 sky130_fd_sc_hd__nor2_2 _16930_ (.A(_04244_),
    .B(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__xnor2_2 _16931_ (.A(_04198_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__nor3_2 _16932_ (.A(_04215_),
    .B(_04218_),
    .C(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__o21ai_2 _16933_ (.A1(_04215_),
    .A2(_04218_),
    .B1(_04247_),
    .Y(_04249_));
 sky130_fd_sc_hd__and2b_2 _16934_ (.A_N(_04248_),
    .B(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__a21bo_2 _16935_ (.A1(_04224_),
    .A2(_04225_),
    .B1_N(_04221_),
    .X(_04251_));
 sky130_fd_sc_hd__xor2_2 _16936_ (.A(_04250_),
    .B(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__mux2_1 _16937_ (.A0(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[13] ),
    .A1(_04252_),
    .S(\systolic_inst.ce_local ),
    .X(_01231_));
 sky130_fd_sc_hd__a31o_2 _16938_ (.A1(\systolic_inst.B_outs[11][5] ),
    .A2(\systolic_inst.A_outs[11][7] ),
    .A3(_04231_),
    .B1(_04230_),
    .X(_04253_));
 sky130_fd_sc_hd__nand3_2 _16939_ (.A(\systolic_inst.B_outs[11][5] ),
    .B(\systolic_inst.B_outs[11][6] ),
    .C(\systolic_inst.A_outs[11][7] ),
    .Y(_04254_));
 sky130_fd_sc_hd__o211a_2 _16940_ (.A1(_11262_),
    .A2(\systolic_inst.A_outs[11][7] ),
    .B1(_04204_),
    .C1(_04227_),
    .X(_04255_));
 sky130_fd_sc_hd__a21oi_2 _16941_ (.A1(_04253_),
    .A2(_04254_),
    .B1(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__or2_2 _16942_ (.A(_04169_),
    .B(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__nand2_2 _16943_ (.A(_04169_),
    .B(_04256_),
    .Y(_04258_));
 sky130_fd_sc_hd__nand2_2 _16944_ (.A(_04257_),
    .B(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__a21oi_2 _16945_ (.A1(_04234_),
    .A2(_04236_),
    .B1(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__and3_2 _16946_ (.A(_04234_),
    .B(_04236_),
    .C(_04259_),
    .X(_04261_));
 sky130_fd_sc_hd__nor2_2 _16947_ (.A(_04260_),
    .B(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__xnor2_2 _16948_ (.A(_04199_),
    .B(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__o21a_2 _16949_ (.A1(_04199_),
    .A2(_04241_),
    .B1(_04240_),
    .X(_04264_));
 sky130_fd_sc_hd__and2b_2 _16950_ (.A_N(_04264_),
    .B(_04263_),
    .X(_04265_));
 sky130_fd_sc_hd__and2b_2 _16951_ (.A_N(_04263_),
    .B(_04264_),
    .X(_04266_));
 sky130_fd_sc_hd__nor2_2 _16952_ (.A(_04265_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__xnor2_2 _16953_ (.A(_04198_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__o21ba_2 _16954_ (.A1(_04198_),
    .A2(_04245_),
    .B1_N(_04244_),
    .X(_04269_));
 sky130_fd_sc_hd__nand2b_2 _16955_ (.A_N(_04269_),
    .B(_04268_),
    .Y(_04270_));
 sky130_fd_sc_hd__xnor2_2 _16956_ (.A(_04268_),
    .B(_04269_),
    .Y(_04271_));
 sky130_fd_sc_hd__o21ai_2 _16957_ (.A1(_04221_),
    .A2(_04248_),
    .B1(_04249_),
    .Y(_04272_));
 sky130_fd_sc_hd__a31o_2 _16958_ (.A1(_04224_),
    .A2(_04225_),
    .A3(_04250_),
    .B1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__nand2_2 _16959_ (.A(_04271_),
    .B(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__xor2_2 _16960_ (.A(_04271_),
    .B(_04273_),
    .X(_04275_));
 sky130_fd_sc_hd__mux2_1 _16961_ (.A0(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[14] ),
    .A1(_04275_),
    .S(\systolic_inst.ce_local ),
    .X(_01232_));
 sky130_fd_sc_hd__a31o_2 _16962_ (.A1(_04056_),
    .A2(_04196_),
    .A3(_04267_),
    .B1(_04265_),
    .X(_04276_));
 sky130_fd_sc_hd__a21oi_2 _16963_ (.A1(_04200_),
    .A2(_04262_),
    .B1(_04260_),
    .Y(_04277_));
 sky130_fd_sc_hd__xnor2_2 _16964_ (.A(_04197_),
    .B(_04257_),
    .Y(_04278_));
 sky130_fd_sc_hd__xnor2_2 _16965_ (.A(_04277_),
    .B(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__xnor2_2 _16966_ (.A(_04276_),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__and3_2 _16967_ (.A(\systolic_inst.ce_local ),
    .B(_04270_),
    .C(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__a22o_2 _16968_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B1(_04274_),
    .B2(_04281_),
    .X(_01233_));
 sky130_fd_sc_hd__a21o_2 _16969_ (.A1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[11][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_04282_));
 sky130_fd_sc_hd__a21oi_2 _16970_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[11][0] ),
    .Y(_04283_));
 sky130_fd_sc_hd__a21oi_2 _16971_ (.A1(\systolic_inst.ce_local ),
    .A2(_04282_),
    .B1(_04283_),
    .Y(_01234_));
 sky130_fd_sc_hd__and2_2 _16972_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[11][1] ),
    .X(_04284_));
 sky130_fd_sc_hd__nand2_2 _16973_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[11][1] ),
    .Y(_04285_));
 sky130_fd_sc_hd__or2_2 _16974_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[11][1] ),
    .X(_04286_));
 sky130_fd_sc_hd__and4_2 _16975_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[11][0] ),
    .C(_04285_),
    .D(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__inv_2 _16976_ (.A(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__a22o_2 _16977_ (.A1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[11][0] ),
    .B1(_04285_),
    .B2(_04286_),
    .X(_04289_));
 sky130_fd_sc_hd__a32o_2 _16978_ (.A1(_11712_),
    .A2(_04288_),
    .A3(_04289_),
    .B1(\systolic_inst.acc_wires[11][1] ),
    .B2(_11258_),
    .X(_01235_));
 sky130_fd_sc_hd__nand2_2 _16979_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[11][2] ),
    .Y(_04290_));
 sky130_fd_sc_hd__or2_2 _16980_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[11][2] ),
    .X(_04291_));
 sky130_fd_sc_hd__a31o_2 _16981_ (.A1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[11][0] ),
    .A3(_04286_),
    .B1(_04284_),
    .X(_04292_));
 sky130_fd_sc_hd__a21o_2 _16982_ (.A1(_04290_),
    .A2(_04291_),
    .B1(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__and3_2 _16983_ (.A(_04290_),
    .B(_04291_),
    .C(_04292_),
    .X(_04294_));
 sky130_fd_sc_hd__inv_2 _16984_ (.A(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__a32o_2 _16985_ (.A1(_11712_),
    .A2(_04293_),
    .A3(_04295_),
    .B1(\systolic_inst.acc_wires[11][2] ),
    .B2(_11258_),
    .X(_01236_));
 sky130_fd_sc_hd__nand2_2 _16986_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[11][3] ),
    .Y(_04296_));
 sky130_fd_sc_hd__or2_2 _16987_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[11][3] ),
    .X(_04297_));
 sky130_fd_sc_hd__a21bo_2 _16988_ (.A1(_04291_),
    .A2(_04292_),
    .B1_N(_04290_),
    .X(_04298_));
 sky130_fd_sc_hd__a21o_2 _16989_ (.A1(_04296_),
    .A2(_04297_),
    .B1(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__and3_2 _16990_ (.A(_04296_),
    .B(_04297_),
    .C(_04298_),
    .X(_04300_));
 sky130_fd_sc_hd__inv_2 _16991_ (.A(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__a32o_2 _16992_ (.A1(_11712_),
    .A2(_04299_),
    .A3(_04301_),
    .B1(\systolic_inst.acc_wires[11][3] ),
    .B2(_11258_),
    .X(_01237_));
 sky130_fd_sc_hd__nand2_2 _16993_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[11][4] ),
    .Y(_04302_));
 sky130_fd_sc_hd__or2_2 _16994_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[11][4] ),
    .X(_04303_));
 sky130_fd_sc_hd__a21bo_2 _16995_ (.A1(_04297_),
    .A2(_04298_),
    .B1_N(_04296_),
    .X(_04304_));
 sky130_fd_sc_hd__a21o_2 _16996_ (.A1(_04302_),
    .A2(_04303_),
    .B1(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__and3_2 _16997_ (.A(_04302_),
    .B(_04303_),
    .C(_04304_),
    .X(_04306_));
 sky130_fd_sc_hd__inv_2 _16998_ (.A(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__a32o_2 _16999_ (.A1(_11712_),
    .A2(_04305_),
    .A3(_04307_),
    .B1(\systolic_inst.acc_wires[11][4] ),
    .B2(_11258_),
    .X(_01238_));
 sky130_fd_sc_hd__nand2_2 _17000_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[11][5] ),
    .Y(_04308_));
 sky130_fd_sc_hd__or2_2 _17001_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[11][5] ),
    .X(_04309_));
 sky130_fd_sc_hd__a21bo_2 _17002_ (.A1(_04303_),
    .A2(_04304_),
    .B1_N(_04302_),
    .X(_04310_));
 sky130_fd_sc_hd__a21o_2 _17003_ (.A1(_04308_),
    .A2(_04309_),
    .B1(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__and3_2 _17004_ (.A(_04308_),
    .B(_04309_),
    .C(_04310_),
    .X(_04312_));
 sky130_fd_sc_hd__inv_2 _17005_ (.A(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__a32o_2 _17006_ (.A1(_11712_),
    .A2(_04311_),
    .A3(_04313_),
    .B1(\systolic_inst.acc_wires[11][5] ),
    .B2(_11258_),
    .X(_01239_));
 sky130_fd_sc_hd__nand2_2 _17007_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[11][6] ),
    .Y(_04314_));
 sky130_fd_sc_hd__or2_2 _17008_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[11][6] ),
    .X(_04315_));
 sky130_fd_sc_hd__a21bo_2 _17009_ (.A1(_04309_),
    .A2(_04310_),
    .B1_N(_04308_),
    .X(_04316_));
 sky130_fd_sc_hd__a21o_2 _17010_ (.A1(_04314_),
    .A2(_04315_),
    .B1(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__and3_2 _17011_ (.A(_04314_),
    .B(_04315_),
    .C(_04316_),
    .X(_04318_));
 sky130_fd_sc_hd__inv_2 _17012_ (.A(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__a32o_2 _17013_ (.A1(_11712_),
    .A2(_04317_),
    .A3(_04319_),
    .B1(\systolic_inst.acc_wires[11][6] ),
    .B2(_11258_),
    .X(_01240_));
 sky130_fd_sc_hd__nand2_2 _17014_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[11][7] ),
    .Y(_04320_));
 sky130_fd_sc_hd__or2_2 _17015_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[11][7] ),
    .X(_04321_));
 sky130_fd_sc_hd__a21bo_2 _17016_ (.A1(_04315_),
    .A2(_04316_),
    .B1_N(_04314_),
    .X(_04322_));
 sky130_fd_sc_hd__a21o_2 _17017_ (.A1(_04320_),
    .A2(_04321_),
    .B1(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__nand3_2 _17018_ (.A(_04320_),
    .B(_04321_),
    .C(_04322_),
    .Y(_04324_));
 sky130_fd_sc_hd__a32o_2 _17019_ (.A1(_11712_),
    .A2(_04323_),
    .A3(_04324_),
    .B1(\systolic_inst.acc_wires[11][7] ),
    .B2(_11258_),
    .X(_01241_));
 sky130_fd_sc_hd__a21bo_2 _17020_ (.A1(_04321_),
    .A2(_04322_),
    .B1_N(_04320_),
    .X(_04325_));
 sky130_fd_sc_hd__xor2_2 _17021_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[11][8] ),
    .X(_04326_));
 sky130_fd_sc_hd__and2_2 _17022_ (.A(_04325_),
    .B(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__o21ai_2 _17023_ (.A1(_04325_),
    .A2(_04326_),
    .B1(_11712_),
    .Y(_04328_));
 sky130_fd_sc_hd__a2bb2o_2 _17024_ (.A1_N(_04328_),
    .A2_N(_04327_),
    .B1(\systolic_inst.acc_wires[11][8] ),
    .B2(_11258_),
    .X(_01242_));
 sky130_fd_sc_hd__xor2_2 _17025_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[11][9] ),
    .X(_04329_));
 sky130_fd_sc_hd__a211o_2 _17026_ (.A1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[11][8] ),
    .B1(_04327_),
    .C1(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__nand2_2 _17027_ (.A(_04326_),
    .B(_04329_),
    .Y(_04331_));
 sky130_fd_sc_hd__nand2_2 _17028_ (.A(_04327_),
    .B(_04329_),
    .Y(_04332_));
 sky130_fd_sc_hd__and3_2 _17029_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[11][8] ),
    .C(_04329_),
    .X(_04333_));
 sky130_fd_sc_hd__nor2_2 _17030_ (.A(_11713_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__a32o_2 _17031_ (.A1(_04330_),
    .A2(_04332_),
    .A3(_04334_),
    .B1(\systolic_inst.acc_wires[11][9] ),
    .B2(_11258_),
    .X(_01243_));
 sky130_fd_sc_hd__nand2_2 _17032_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[11][10] ),
    .Y(_04335_));
 sky130_fd_sc_hd__or2_2 _17033_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[11][10] ),
    .X(_04336_));
 sky130_fd_sc_hd__and2_2 _17034_ (.A(_04335_),
    .B(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__a21oi_2 _17035_ (.A1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[11][9] ),
    .B1(_04333_),
    .Y(_04338_));
 sky130_fd_sc_hd__nand2_2 _17036_ (.A(_04332_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__xor2_2 _17037_ (.A(_04337_),
    .B(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__a22o_2 _17038_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][10] ),
    .B1(_11712_),
    .B2(_04340_),
    .X(_01244_));
 sky130_fd_sc_hd__nor2_2 _17039_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[11][11] ),
    .Y(_04341_));
 sky130_fd_sc_hd__or2_2 _17040_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[11][11] ),
    .X(_04342_));
 sky130_fd_sc_hd__nand2_2 _17041_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[11][11] ),
    .Y(_04343_));
 sky130_fd_sc_hd__nand2_2 _17042_ (.A(_04342_),
    .B(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__a21bo_2 _17043_ (.A1(_04337_),
    .A2(_04339_),
    .B1_N(_04335_),
    .X(_04345_));
 sky130_fd_sc_hd__xnor2_2 _17044_ (.A(_04344_),
    .B(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__a22o_2 _17045_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][11] ),
    .B1(_11712_),
    .B2(_04346_),
    .X(_01245_));
 sky130_fd_sc_hd__nand3_2 _17046_ (.A(_04337_),
    .B(_04342_),
    .C(_04343_),
    .Y(_04347_));
 sky130_fd_sc_hd__nor2_2 _17047_ (.A(_04331_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__o2bb2a_2 _17048_ (.A1_N(_04325_),
    .A2_N(_04348_),
    .B1(_04338_),
    .B2(_04347_),
    .X(_04349_));
 sky130_fd_sc_hd__o21a_2 _17049_ (.A1(_04335_),
    .A2(_04341_),
    .B1(_04343_),
    .X(_04350_));
 sky130_fd_sc_hd__xnor2_2 _17050_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[11][12] ),
    .Y(_04351_));
 sky130_fd_sc_hd__and3_2 _17051_ (.A(_04349_),
    .B(_04350_),
    .C(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__a21oi_2 _17052_ (.A1(_04349_),
    .A2(_04350_),
    .B1(_04351_),
    .Y(_04353_));
 sky130_fd_sc_hd__nor2_2 _17053_ (.A(_04352_),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__a22o_2 _17054_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][12] ),
    .B1(_11712_),
    .B2(_04354_),
    .X(_01246_));
 sky130_fd_sc_hd__xor2_2 _17055_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[11][13] ),
    .X(_04355_));
 sky130_fd_sc_hd__a211o_2 _17056_ (.A1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[11][12] ),
    .B1(_04353_),
    .C1(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__nand2b_2 _17057_ (.A_N(_04351_),
    .B(_04355_),
    .Y(_04357_));
 sky130_fd_sc_hd__a21o_2 _17058_ (.A1(_04349_),
    .A2(_04350_),
    .B1(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__and3_2 _17059_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[11][12] ),
    .C(_04355_),
    .X(_04359_));
 sky130_fd_sc_hd__nor2_2 _17060_ (.A(_11713_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__a32o_2 _17061_ (.A1(_04356_),
    .A2(_04358_),
    .A3(_04360_),
    .B1(\systolic_inst.acc_wires[11][13] ),
    .B2(_11258_),
    .X(_01247_));
 sky130_fd_sc_hd__or2_2 _17062_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[11][14] ),
    .X(_04361_));
 sky130_fd_sc_hd__nand2_2 _17063_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[11][14] ),
    .Y(_04362_));
 sky130_fd_sc_hd__and2_2 _17064_ (.A(_04361_),
    .B(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__nand2_2 _17065_ (.A(_04361_),
    .B(_04362_),
    .Y(_04364_));
 sky130_fd_sc_hd__a21oi_2 _17066_ (.A1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[11][13] ),
    .B1(_04359_),
    .Y(_04365_));
 sky130_fd_sc_hd__nand2_2 _17067_ (.A(_04358_),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_2 _17068_ (.A(_04363_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__or2_2 _17069_ (.A(_04363_),
    .B(_04366_),
    .X(_04368_));
 sky130_fd_sc_hd__a32o_2 _17070_ (.A1(_11712_),
    .A2(_04367_),
    .A3(_04368_),
    .B1(\systolic_inst.acc_wires[11][14] ),
    .B2(_11258_),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_2 _17071_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][15] ),
    .Y(_04369_));
 sky130_fd_sc_hd__and2_2 _17072_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][15] ),
    .X(_04370_));
 sky130_fd_sc_hd__or2_2 _17073_ (.A(_04369_),
    .B(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__a21oi_2 _17074_ (.A1(_04362_),
    .A2(_04367_),
    .B1(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__a31o_2 _17075_ (.A1(_04362_),
    .A2(_04367_),
    .A3(_04371_),
    .B1(_11713_),
    .X(_04373_));
 sky130_fd_sc_hd__a2bb2o_2 _17076_ (.A1_N(_04373_),
    .A2_N(_04372_),
    .B1(\systolic_inst.acc_wires[11][15] ),
    .B2(_11258_),
    .X(_01249_));
 sky130_fd_sc_hd__a211o_2 _17077_ (.A1(_04358_),
    .A2(_04365_),
    .B1(_04371_),
    .C1(_04364_),
    .X(_04374_));
 sky130_fd_sc_hd__o21ba_2 _17078_ (.A1(_04362_),
    .A2(_04369_),
    .B1_N(_04370_),
    .X(_04375_));
 sky130_fd_sc_hd__and2_2 _17079_ (.A(_04374_),
    .B(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__xnor2_2 _17080_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][16] ),
    .Y(_04377_));
 sky130_fd_sc_hd__nand2_2 _17081_ (.A(_04376_),
    .B(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__nor2_2 _17082_ (.A(_04376_),
    .B(_04377_),
    .Y(_04379_));
 sky130_fd_sc_hd__nor2_2 _17083_ (.A(_11713_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__a22o_2 _17084_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][16] ),
    .B1(_04378_),
    .B2(_04380_),
    .X(_01250_));
 sky130_fd_sc_hd__xor2_2 _17085_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][17] ),
    .X(_04381_));
 sky130_fd_sc_hd__inv_2 _17086_ (.A(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__a21oi_2 _17087_ (.A1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[11][16] ),
    .B1(_04379_),
    .Y(_04383_));
 sky130_fd_sc_hd__xnor2_2 _17088_ (.A(_04381_),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__a22o_2 _17089_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][17] ),
    .B1(_11712_),
    .B2(_04384_),
    .X(_01251_));
 sky130_fd_sc_hd__or2_2 _17090_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][18] ),
    .X(_04385_));
 sky130_fd_sc_hd__nand2_2 _17091_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][18] ),
    .Y(_04386_));
 sky130_fd_sc_hd__nand2_2 _17092_ (.A(_04385_),
    .B(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__o21a_2 _17093_ (.A1(\systolic_inst.acc_wires[11][16] ),
    .A2(\systolic_inst.acc_wires[11][17] ),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .X(_04388_));
 sky130_fd_sc_hd__a21oi_2 _17094_ (.A1(_04379_),
    .A2(_04381_),
    .B1(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__xor2_2 _17095_ (.A(_04387_),
    .B(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__a22o_2 _17096_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][18] ),
    .B1(_11712_),
    .B2(_04390_),
    .X(_01252_));
 sky130_fd_sc_hd__xnor2_2 _17097_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][19] ),
    .Y(_04391_));
 sky130_fd_sc_hd__o21ai_2 _17098_ (.A1(_04387_),
    .A2(_04389_),
    .B1(_04386_),
    .Y(_04392_));
 sky130_fd_sc_hd__xnor2_2 _17099_ (.A(_04391_),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__a22o_2 _17100_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][19] ),
    .B1(_11712_),
    .B2(_04393_),
    .X(_01253_));
 sky130_fd_sc_hd__or2_2 _17101_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][20] ),
    .X(_04394_));
 sky130_fd_sc_hd__nand2_2 _17102_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][20] ),
    .Y(_04395_));
 sky130_fd_sc_hd__and2_2 _17103_ (.A(_04394_),
    .B(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__or4_2 _17104_ (.A(_04377_),
    .B(_04382_),
    .C(_04387_),
    .D(_04391_),
    .X(_04397_));
 sky130_fd_sc_hd__nor2_2 _17105_ (.A(_04376_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__o41a_2 _17106_ (.A1(\systolic_inst.acc_wires[11][16] ),
    .A2(\systolic_inst.acc_wires[11][17] ),
    .A3(\systolic_inst.acc_wires[11][18] ),
    .A4(\systolic_inst.acc_wires[11][19] ),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .X(_04399_));
 sky130_fd_sc_hd__or3_2 _17107_ (.A(_04396_),
    .B(_04398_),
    .C(_04399_),
    .X(_04400_));
 sky130_fd_sc_hd__o21ai_2 _17108_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04396_),
    .Y(_04401_));
 sky130_fd_sc_hd__a32o_2 _17109_ (.A1(_11712_),
    .A2(_04400_),
    .A3(_04401_),
    .B1(\systolic_inst.acc_wires[11][20] ),
    .B2(_11258_),
    .X(_01254_));
 sky130_fd_sc_hd__xnor2_2 _17110_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][21] ),
    .Y(_04402_));
 sky130_fd_sc_hd__inv_2 _17111_ (.A(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__a21oi_2 _17112_ (.A1(_04395_),
    .A2(_04401_),
    .B1(_04402_),
    .Y(_04404_));
 sky130_fd_sc_hd__a31o_2 _17113_ (.A1(_04395_),
    .A2(_04401_),
    .A3(_04402_),
    .B1(_11713_),
    .X(_04405_));
 sky130_fd_sc_hd__a2bb2o_2 _17114_ (.A1_N(_04405_),
    .A2_N(_04404_),
    .B1(\systolic_inst.acc_wires[11][21] ),
    .B2(_11258_),
    .X(_01255_));
 sky130_fd_sc_hd__or2_2 _17115_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][22] ),
    .X(_04406_));
 sky130_fd_sc_hd__nand2_2 _17116_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][22] ),
    .Y(_04407_));
 sky130_fd_sc_hd__and2_2 _17117_ (.A(_04406_),
    .B(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__o21a_2 _17118_ (.A1(\systolic_inst.acc_wires[11][20] ),
    .A2(\systolic_inst.acc_wires[11][21] ),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .X(_04409_));
 sky130_fd_sc_hd__nor2_2 _17119_ (.A(_04401_),
    .B(_04402_),
    .Y(_04410_));
 sky130_fd_sc_hd__o21ai_2 _17120_ (.A1(_04409_),
    .A2(_04410_),
    .B1(_04408_),
    .Y(_04411_));
 sky130_fd_sc_hd__or3_2 _17121_ (.A(_04408_),
    .B(_04409_),
    .C(_04410_),
    .X(_04412_));
 sky130_fd_sc_hd__a32o_2 _17122_ (.A1(_11712_),
    .A2(_04411_),
    .A3(_04412_),
    .B1(\systolic_inst.acc_wires[11][22] ),
    .B2(_11258_),
    .X(_01256_));
 sky130_fd_sc_hd__xor2_2 _17123_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][23] ),
    .X(_04413_));
 sky130_fd_sc_hd__inv_2 _17124_ (.A(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__nand3_2 _17125_ (.A(_04407_),
    .B(_04411_),
    .C(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__a21o_2 _17126_ (.A1(_04407_),
    .A2(_04411_),
    .B1(_04414_),
    .X(_04416_));
 sky130_fd_sc_hd__a32o_2 _17127_ (.A1(_11712_),
    .A2(_04415_),
    .A3(_04416_),
    .B1(\systolic_inst.acc_wires[11][23] ),
    .B2(_11258_),
    .X(_01257_));
 sky130_fd_sc_hd__nand4_2 _17128_ (.A(_04396_),
    .B(_04403_),
    .C(_04408_),
    .D(_04413_),
    .Y(_04417_));
 sky130_fd_sc_hd__a211o_2 _17129_ (.A1(_04374_),
    .A2(_04375_),
    .B1(_04397_),
    .C1(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__o41a_2 _17130_ (.A1(\systolic_inst.acc_wires[11][20] ),
    .A2(\systolic_inst.acc_wires[11][21] ),
    .A3(\systolic_inst.acc_wires[11][22] ),
    .A4(\systolic_inst.acc_wires[11][23] ),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .X(_04419_));
 sky130_fd_sc_hd__nor2_2 _17131_ (.A(_04399_),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__nor2_2 _17132_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][24] ),
    .Y(_04421_));
 sky130_fd_sc_hd__and2_2 _17133_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][24] ),
    .X(_04422_));
 sky130_fd_sc_hd__or2_2 _17134_ (.A(_04421_),
    .B(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__a21oi_2 _17135_ (.A1(_04418_),
    .A2(_04420_),
    .B1(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__a31o_2 _17136_ (.A1(_04418_),
    .A2(_04420_),
    .A3(_04423_),
    .B1(_11713_),
    .X(_04425_));
 sky130_fd_sc_hd__a2bb2o_2 _17137_ (.A1_N(_04425_),
    .A2_N(_04424_),
    .B1(\systolic_inst.acc_wires[11][24] ),
    .B2(_11258_),
    .X(_01258_));
 sky130_fd_sc_hd__xor2_2 _17138_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][25] ),
    .X(_04426_));
 sky130_fd_sc_hd__or3_2 _17139_ (.A(_04422_),
    .B(_04424_),
    .C(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__o21ai_2 _17140_ (.A1(_04422_),
    .A2(_04424_),
    .B1(_04426_),
    .Y(_04428_));
 sky130_fd_sc_hd__a32o_2 _17141_ (.A1(_11712_),
    .A2(_04427_),
    .A3(_04428_),
    .B1(\systolic_inst.acc_wires[11][25] ),
    .B2(_11258_),
    .X(_01259_));
 sky130_fd_sc_hd__or2_2 _17142_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][26] ),
    .X(_04429_));
 sky130_fd_sc_hd__nand2_2 _17143_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][26] ),
    .Y(_04430_));
 sky130_fd_sc_hd__nand2_2 _17144_ (.A(_04429_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__o21a_2 _17145_ (.A1(\systolic_inst.acc_wires[11][24] ),
    .A2(\systolic_inst.acc_wires[11][25] ),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .X(_04432_));
 sky130_fd_sc_hd__a21o_2 _17146_ (.A1(_04424_),
    .A2(_04426_),
    .B1(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__xnor2_2 _17147_ (.A(_04431_),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__a22o_2 _17148_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][26] ),
    .B1(_11712_),
    .B2(_04434_),
    .X(_01260_));
 sky130_fd_sc_hd__xnor2_2 _17149_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][27] ),
    .Y(_04435_));
 sky130_fd_sc_hd__a21bo_2 _17150_ (.A1(_04429_),
    .A2(_04433_),
    .B1_N(_04430_),
    .X(_04436_));
 sky130_fd_sc_hd__xnor2_2 _17151_ (.A(_04435_),
    .B(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__a22o_2 _17152_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][27] ),
    .B1(_11712_),
    .B2(_04437_),
    .X(_01261_));
 sky130_fd_sc_hd__nor2_2 _17153_ (.A(_04431_),
    .B(_04435_),
    .Y(_04438_));
 sky130_fd_sc_hd__o21a_2 _17154_ (.A1(\systolic_inst.acc_wires[11][26] ),
    .A2(\systolic_inst.acc_wires[11][27] ),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .X(_04439_));
 sky130_fd_sc_hd__a311oi_2 _17155_ (.A1(_04424_),
    .A2(_04426_),
    .A3(_04438_),
    .B1(_04439_),
    .C1(_04432_),
    .Y(_04440_));
 sky130_fd_sc_hd__or2_2 _17156_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][28] ),
    .X(_04441_));
 sky130_fd_sc_hd__nand2_2 _17157_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][28] ),
    .Y(_04442_));
 sky130_fd_sc_hd__nand2_2 _17158_ (.A(_04441_),
    .B(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__xor2_2 _17159_ (.A(_04440_),
    .B(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__a22o_2 _17160_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][28] ),
    .B1(_11712_),
    .B2(_04444_),
    .X(_01262_));
 sky130_fd_sc_hd__xor2_2 _17161_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][29] ),
    .X(_04445_));
 sky130_fd_sc_hd__inv_2 _17162_ (.A(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__o21a_2 _17163_ (.A1(_04440_),
    .A2(_04443_),
    .B1(_04442_),
    .X(_04447_));
 sky130_fd_sc_hd__xnor2_2 _17164_ (.A(_04445_),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__a22o_2 _17165_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[11][29] ),
    .B1(_11712_),
    .B2(_04448_),
    .X(_01263_));
 sky130_fd_sc_hd__o21ai_2 _17166_ (.A1(\systolic_inst.acc_wires[11][28] ),
    .A2(\systolic_inst.acc_wires[11][29] ),
    .B1(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .Y(_04449_));
 sky130_fd_sc_hd__o31a_2 _17167_ (.A1(_04440_),
    .A2(_04443_),
    .A3(_04446_),
    .B1(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__nand2_2 _17168_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][30] ),
    .Y(_04451_));
 sky130_fd_sc_hd__or2_2 _17169_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][30] ),
    .X(_04452_));
 sky130_fd_sc_hd__nand2_2 _17170_ (.A(_04451_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand2_2 _17171_ (.A(_04450_),
    .B(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__or2_2 _17172_ (.A(_04450_),
    .B(_04453_),
    .X(_04455_));
 sky130_fd_sc_hd__a32o_2 _17173_ (.A1(_11712_),
    .A2(_04454_),
    .A3(_04455_),
    .B1(\systolic_inst.acc_wires[11][30] ),
    .B2(_11258_),
    .X(_01264_));
 sky130_fd_sc_hd__xnor2_2 _17174_ (.A(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[11][31] ),
    .Y(_04456_));
 sky130_fd_sc_hd__a21oi_2 _17175_ (.A1(_04451_),
    .A2(_04455_),
    .B1(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__a31o_2 _17176_ (.A1(_04451_),
    .A2(_04455_),
    .A3(_04456_),
    .B1(_11713_),
    .X(_04458_));
 sky130_fd_sc_hd__a2bb2o_2 _17177_ (.A1_N(_04458_),
    .A2_N(_04457_),
    .B1(\systolic_inst.acc_wires[11][31] ),
    .B2(_11258_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _17178_ (.A0(\systolic_inst.A_outs[10][0] ),
    .A1(\systolic_inst.A_outs[9][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _17179_ (.A0(\systolic_inst.A_outs[10][1] ),
    .A1(\systolic_inst.A_outs[9][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _17180_ (.A0(\systolic_inst.A_outs[10][2] ),
    .A1(\systolic_inst.A_outs[9][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _17181_ (.A0(\systolic_inst.A_outs[10][3] ),
    .A1(\systolic_inst.A_outs[9][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _17182_ (.A0(\systolic_inst.A_outs[10][4] ),
    .A1(\systolic_inst.A_outs[9][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _17183_ (.A0(\systolic_inst.A_outs[10][5] ),
    .A1(\systolic_inst.A_outs[9][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _17184_ (.A0(\systolic_inst.A_outs[10][6] ),
    .A1(\systolic_inst.A_outs[9][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _17185_ (.A0(\systolic_inst.A_outs[10][7] ),
    .A1(\systolic_inst.A_outs[9][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _17186_ (.A0(\systolic_inst.B_outs[9][0] ),
    .A1(\systolic_inst.B_outs[5][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _17187_ (.A0(\systolic_inst.B_outs[9][1] ),
    .A1(\systolic_inst.B_outs[5][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _17188_ (.A0(\systolic_inst.B_outs[9][2] ),
    .A1(\systolic_inst.B_outs[5][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _17189_ (.A0(\systolic_inst.B_outs[9][3] ),
    .A1(\systolic_inst.B_outs[5][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _17190_ (.A0(\systolic_inst.B_outs[9][4] ),
    .A1(\systolic_inst.B_outs[5][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _17191_ (.A0(\systolic_inst.B_outs[9][5] ),
    .A1(\systolic_inst.B_outs[5][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _17192_ (.A0(\systolic_inst.B_outs[9][6] ),
    .A1(\systolic_inst.B_outs[5][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _17193_ (.A0(\systolic_inst.B_outs[9][7] ),
    .A1(\systolic_inst.B_outs[5][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01281_));
 sky130_fd_sc_hd__and3_2 _17194_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[10][0] ),
    .C(\systolic_inst.A_outs[10][0] ),
    .X(_04459_));
 sky130_fd_sc_hd__a21o_2 _17195_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[0] ),
    .B1(_04459_),
    .X(_01282_));
 sky130_fd_sc_hd__and4_2 _17196_ (.A(\systolic_inst.B_outs[10][0] ),
    .B(\systolic_inst.A_outs[10][0] ),
    .C(\systolic_inst.B_outs[10][1] ),
    .D(\systolic_inst.A_outs[10][1] ),
    .X(_04460_));
 sky130_fd_sc_hd__inv_2 _17197_ (.A(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__a22o_2 _17198_ (.A1(\systolic_inst.A_outs[10][0] ),
    .A2(\systolic_inst.B_outs[10][1] ),
    .B1(\systolic_inst.A_outs[10][1] ),
    .B2(\systolic_inst.B_outs[10][0] ),
    .X(_04462_));
 sky130_fd_sc_hd__and2_2 _17199_ (.A(\systolic_inst.ce_local ),
    .B(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__a22o_2 _17200_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[1] ),
    .B1(_04461_),
    .B2(_04463_),
    .X(_01283_));
 sky130_fd_sc_hd__nand2_2 _17201_ (.A(\systolic_inst.B_outs[10][1] ),
    .B(\systolic_inst.A_outs[10][1] ),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_2 _17202_ (.A(\systolic_inst.B_outs[10][0] ),
    .B(\systolic_inst.A_outs[10][2] ),
    .Y(_04465_));
 sky130_fd_sc_hd__and4_2 _17203_ (.A(\systolic_inst.B_outs[10][0] ),
    .B(\systolic_inst.B_outs[10][1] ),
    .C(\systolic_inst.A_outs[10][1] ),
    .D(\systolic_inst.A_outs[10][2] ),
    .X(_04466_));
 sky130_fd_sc_hd__a21o_2 _17204_ (.A1(_04464_),
    .A2(_04465_),
    .B1(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__or2_2 _17205_ (.A(_04461_),
    .B(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__xnor2_2 _17206_ (.A(_04460_),
    .B(_04467_),
    .Y(_04469_));
 sky130_fd_sc_hd__and2_2 _17207_ (.A(\systolic_inst.A_outs[10][0] ),
    .B(\systolic_inst.B_outs[10][2] ),
    .X(_04470_));
 sky130_fd_sc_hd__nand2_2 _17208_ (.A(_04469_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__o21a_2 _17209_ (.A1(_04469_),
    .A2(_04470_),
    .B1(\systolic_inst.ce_local ),
    .X(_04472_));
 sky130_fd_sc_hd__a22o_2 _17210_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[2] ),
    .B1(_04471_),
    .B2(_04472_),
    .X(_01284_));
 sky130_fd_sc_hd__a22oi_2 _17211_ (.A1(\systolic_inst.A_outs[10][1] ),
    .A2(\systolic_inst.B_outs[10][2] ),
    .B1(\systolic_inst.B_outs[10][3] ),
    .B2(\systolic_inst.A_outs[10][0] ),
    .Y(_04473_));
 sky130_fd_sc_hd__and3_2 _17212_ (.A(\systolic_inst.A_outs[10][0] ),
    .B(\systolic_inst.A_outs[10][1] ),
    .C(\systolic_inst.B_outs[10][3] ),
    .X(_04474_));
 sky130_fd_sc_hd__and2_2 _17213_ (.A(\systolic_inst.B_outs[10][2] ),
    .B(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__nand2_2 _17214_ (.A(\systolic_inst.B_outs[10][1] ),
    .B(\systolic_inst.A_outs[10][3] ),
    .Y(_04476_));
 sky130_fd_sc_hd__or2_2 _17215_ (.A(_04465_),
    .B(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__a22o_2 _17216_ (.A1(\systolic_inst.B_outs[10][1] ),
    .A2(\systolic_inst.A_outs[10][2] ),
    .B1(\systolic_inst.A_outs[10][3] ),
    .B2(\systolic_inst.B_outs[10][0] ),
    .X(_04478_));
 sky130_fd_sc_hd__and3_2 _17217_ (.A(_04466_),
    .B(_04477_),
    .C(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__a21oi_2 _17218_ (.A1(_04477_),
    .A2(_04478_),
    .B1(_04466_),
    .Y(_04480_));
 sky130_fd_sc_hd__nor4_2 _17219_ (.A(_04473_),
    .B(_04475_),
    .C(_04479_),
    .D(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__o22a_2 _17220_ (.A1(_04473_),
    .A2(_04475_),
    .B1(_04479_),
    .B2(_04480_),
    .X(_04482_));
 sky130_fd_sc_hd__a211o_2 _17221_ (.A1(_04468_),
    .A2(_04471_),
    .B1(_04481_),
    .C1(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__o211a_2 _17222_ (.A1(_04481_),
    .A2(_04482_),
    .B1(_04468_),
    .C1(_04471_),
    .X(_04484_));
 sky130_fd_sc_hd__nor2_2 _17223_ (.A(_11258_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__a22o_2 _17224_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[3] ),
    .B1(_04483_),
    .B2(_04485_),
    .X(_01285_));
 sky130_fd_sc_hd__nand2_2 _17225_ (.A(\systolic_inst.B_outs[10][2] ),
    .B(\systolic_inst.A_outs[10][2] ),
    .Y(_04486_));
 sky130_fd_sc_hd__a22o_2 _17226_ (.A1(\systolic_inst.A_outs[10][1] ),
    .A2(\systolic_inst.B_outs[10][3] ),
    .B1(\systolic_inst.B_outs[10][4] ),
    .B2(\systolic_inst.A_outs[10][0] ),
    .X(_04487_));
 sky130_fd_sc_hd__a21bo_2 _17227_ (.A1(\systolic_inst.B_outs[10][4] ),
    .A2(_04474_),
    .B1_N(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__xnor2_2 _17228_ (.A(_04486_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__nand2_2 _17229_ (.A(\systolic_inst.B_outs[10][0] ),
    .B(\systolic_inst.A_outs[10][4] ),
    .Y(_04490_));
 sky130_fd_sc_hd__and4_2 _17230_ (.A(\systolic_inst.B_outs[10][0] ),
    .B(\systolic_inst.B_outs[10][1] ),
    .C(\systolic_inst.A_outs[10][3] ),
    .D(\systolic_inst.A_outs[10][4] ),
    .X(_04491_));
 sky130_fd_sc_hd__a21oi_2 _17231_ (.A1(_04476_),
    .A2(_04490_),
    .B1(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__xnor2_2 _17232_ (.A(_04475_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__nor2_2 _17233_ (.A(_04477_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__xnor2_2 _17234_ (.A(_04477_),
    .B(_04493_),
    .Y(_04495_));
 sky130_fd_sc_hd__nor2_2 _17235_ (.A(_04489_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__xnor2_2 _17236_ (.A(_04489_),
    .B(_04495_),
    .Y(_04497_));
 sky130_fd_sc_hd__o21bai_2 _17237_ (.A1(_04479_),
    .A2(_04481_),
    .B1_N(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__or3b_2 _17238_ (.A(_04479_),
    .B(_04481_),
    .C_N(_04497_),
    .X(_04499_));
 sky130_fd_sc_hd__nand2_2 _17239_ (.A(_04498_),
    .B(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__nand2_2 _17240_ (.A(_04483_),
    .B(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__nor2_2 _17241_ (.A(_04483_),
    .B(_04500_),
    .Y(_04502_));
 sky130_fd_sc_hd__nor2_2 _17242_ (.A(_11258_),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__a22o_2 _17243_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[4] ),
    .B1(_04501_),
    .B2(_04503_),
    .X(_01286_));
 sky130_fd_sc_hd__a21oi_2 _17244_ (.A1(_04475_),
    .A2(_04492_),
    .B1(_04494_),
    .Y(_04504_));
 sky130_fd_sc_hd__a32o_2 _17245_ (.A1(\systolic_inst.B_outs[10][2] ),
    .A2(\systolic_inst.A_outs[10][2] ),
    .A3(_04487_),
    .B1(_04474_),
    .B2(\systolic_inst.B_outs[10][4] ),
    .X(_04505_));
 sky130_fd_sc_hd__a22oi_2 _17246_ (.A1(\systolic_inst.B_outs[10][1] ),
    .A2(\systolic_inst.A_outs[10][4] ),
    .B1(\systolic_inst.A_outs[10][5] ),
    .B2(\systolic_inst.B_outs[10][0] ),
    .Y(_04506_));
 sky130_fd_sc_hd__and4_2 _17247_ (.A(\systolic_inst.B_outs[10][0] ),
    .B(\systolic_inst.B_outs[10][1] ),
    .C(\systolic_inst.A_outs[10][4] ),
    .D(\systolic_inst.A_outs[10][5] ),
    .X(_04507_));
 sky130_fd_sc_hd__or2_2 _17248_ (.A(_04506_),
    .B(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__nand2b_2 _17249_ (.A_N(_04508_),
    .B(_04505_),
    .Y(_04509_));
 sky130_fd_sc_hd__xnor2_2 _17250_ (.A(_04505_),
    .B(_04508_),
    .Y(_04510_));
 sky130_fd_sc_hd__xnor2_2 _17251_ (.A(_04491_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__nand2_2 _17252_ (.A(\systolic_inst.A_outs[10][0] ),
    .B(\systolic_inst.B_outs[10][5] ),
    .Y(_04512_));
 sky130_fd_sc_hd__and2_2 _17253_ (.A(\systolic_inst.B_outs[10][2] ),
    .B(\systolic_inst.A_outs[10][3] ),
    .X(_04513_));
 sky130_fd_sc_hd__nand4_2 _17254_ (.A(\systolic_inst.A_outs[10][1] ),
    .B(\systolic_inst.A_outs[10][2] ),
    .C(\systolic_inst.B_outs[10][3] ),
    .D(\systolic_inst.B_outs[10][4] ),
    .Y(_04514_));
 sky130_fd_sc_hd__a22o_2 _17255_ (.A1(\systolic_inst.A_outs[10][2] ),
    .A2(\systolic_inst.B_outs[10][3] ),
    .B1(\systolic_inst.B_outs[10][4] ),
    .B2(\systolic_inst.A_outs[10][1] ),
    .X(_04515_));
 sky130_fd_sc_hd__and3_2 _17256_ (.A(_04513_),
    .B(_04514_),
    .C(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__a21o_2 _17257_ (.A1(_04514_),
    .A2(_04515_),
    .B1(_04513_),
    .X(_04517_));
 sky130_fd_sc_hd__and2b_2 _17258_ (.A_N(_04516_),
    .B(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__and4b_2 _17259_ (.A_N(_04516_),
    .B(_04517_),
    .C(\systolic_inst.A_outs[10][0] ),
    .D(\systolic_inst.B_outs[10][5] ),
    .X(_04519_));
 sky130_fd_sc_hd__xor2_2 _17260_ (.A(_04512_),
    .B(_04518_),
    .X(_04520_));
 sky130_fd_sc_hd__nor2_2 _17261_ (.A(_04511_),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__xor2_2 _17262_ (.A(_04511_),
    .B(_04520_),
    .X(_04522_));
 sky130_fd_sc_hd__nand2_2 _17263_ (.A(_04496_),
    .B(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__xor2_2 _17264_ (.A(_04496_),
    .B(_04522_),
    .X(_04524_));
 sky130_fd_sc_hd__nand2b_2 _17265_ (.A_N(_04504_),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__xnor2_2 _17266_ (.A(_04504_),
    .B(_04524_),
    .Y(_04526_));
 sky130_fd_sc_hd__and2b_2 _17267_ (.A_N(_04498_),
    .B(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__xnor2_2 _17268_ (.A(_04498_),
    .B(_04526_),
    .Y(_04528_));
 sky130_fd_sc_hd__xor2_2 _17269_ (.A(_04502_),
    .B(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__mux2_1 _17270_ (.A0(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[5] ),
    .A1(_04529_),
    .S(\systolic_inst.ce_local ),
    .X(_01287_));
 sky130_fd_sc_hd__a21bo_2 _17271_ (.A1(_04491_),
    .A2(_04510_),
    .B1_N(_04509_),
    .X(_04530_));
 sky130_fd_sc_hd__a21bo_2 _17272_ (.A1(_04513_),
    .A2(_04515_),
    .B1_N(_04514_),
    .X(_04531_));
 sky130_fd_sc_hd__a22oi_2 _17273_ (.A1(\systolic_inst.B_outs[10][1] ),
    .A2(\systolic_inst.A_outs[10][5] ),
    .B1(\systolic_inst.A_outs[10][6] ),
    .B2(\systolic_inst.B_outs[10][0] ),
    .Y(_04532_));
 sky130_fd_sc_hd__and4_2 _17274_ (.A(\systolic_inst.B_outs[10][0] ),
    .B(\systolic_inst.B_outs[10][1] ),
    .C(\systolic_inst.A_outs[10][5] ),
    .D(\systolic_inst.A_outs[10][6] ),
    .X(_04533_));
 sky130_fd_sc_hd__or2_2 _17275_ (.A(_04532_),
    .B(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__and2b_2 _17276_ (.A_N(_04534_),
    .B(_04531_),
    .X(_04535_));
 sky130_fd_sc_hd__xnor2_2 _17277_ (.A(_04531_),
    .B(_04534_),
    .Y(_04536_));
 sky130_fd_sc_hd__xor2_2 _17278_ (.A(_04507_),
    .B(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__nand4_2 _17279_ (.A(\systolic_inst.A_outs[10][2] ),
    .B(\systolic_inst.B_outs[10][3] ),
    .C(\systolic_inst.A_outs[10][3] ),
    .D(\systolic_inst.B_outs[10][4] ),
    .Y(_04538_));
 sky130_fd_sc_hd__a22o_2 _17280_ (.A1(\systolic_inst.B_outs[10][3] ),
    .A2(\systolic_inst.A_outs[10][3] ),
    .B1(\systolic_inst.B_outs[10][4] ),
    .B2(\systolic_inst.A_outs[10][2] ),
    .X(_04539_));
 sky130_fd_sc_hd__nand4_2 _17281_ (.A(\systolic_inst.B_outs[10][2] ),
    .B(\systolic_inst.A_outs[10][4] ),
    .C(_04538_),
    .D(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__a22o_2 _17282_ (.A1(\systolic_inst.B_outs[10][2] ),
    .A2(\systolic_inst.A_outs[10][4] ),
    .B1(_04538_),
    .B2(_04539_),
    .X(_04541_));
 sky130_fd_sc_hd__a22oi_2 _17283_ (.A1(\systolic_inst.A_outs[10][1] ),
    .A2(\systolic_inst.B_outs[10][5] ),
    .B1(\systolic_inst.B_outs[10][6] ),
    .B2(\systolic_inst.A_outs[10][0] ),
    .Y(_04542_));
 sky130_fd_sc_hd__nand2_2 _17284_ (.A(\systolic_inst.A_outs[10][1] ),
    .B(\systolic_inst.B_outs[10][6] ),
    .Y(_04543_));
 sky130_fd_sc_hd__and4_2 _17285_ (.A(\systolic_inst.A_outs[10][0] ),
    .B(\systolic_inst.A_outs[10][1] ),
    .C(\systolic_inst.B_outs[10][5] ),
    .D(\systolic_inst.B_outs[10][6] ),
    .X(_04544_));
 sky130_fd_sc_hd__nor2_2 _17286_ (.A(_04542_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand3_2 _17287_ (.A(_04540_),
    .B(_04541_),
    .C(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__a21o_2 _17288_ (.A1(_04540_),
    .A2(_04541_),
    .B1(_04545_),
    .X(_04547_));
 sky130_fd_sc_hd__and3_2 _17289_ (.A(_04519_),
    .B(_04546_),
    .C(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__a21oi_2 _17290_ (.A1(_04546_),
    .A2(_04547_),
    .B1(_04519_),
    .Y(_04549_));
 sky130_fd_sc_hd__or3b_2 _17291_ (.A(_04548_),
    .B(_04549_),
    .C_N(_04537_),
    .X(_04550_));
 sky130_fd_sc_hd__o21bai_2 _17292_ (.A1(_04548_),
    .A2(_04549_),
    .B1_N(_04537_),
    .Y(_04551_));
 sky130_fd_sc_hd__nand3_2 _17293_ (.A(_04521_),
    .B(_04550_),
    .C(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a21o_2 _17294_ (.A1(_04550_),
    .A2(_04551_),
    .B1(_04521_),
    .X(_04553_));
 sky130_fd_sc_hd__and3_2 _17295_ (.A(_04530_),
    .B(_04552_),
    .C(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__a21oi_2 _17296_ (.A1(_04552_),
    .A2(_04553_),
    .B1(_04530_),
    .Y(_04555_));
 sky130_fd_sc_hd__a211o_2 _17297_ (.A1(_04523_),
    .A2(_04525_),
    .B1(_04554_),
    .C1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__o211ai_2 _17298_ (.A1(_04554_),
    .A2(_04555_),
    .B1(_04523_),
    .C1(_04525_),
    .Y(_04557_));
 sky130_fd_sc_hd__nand2_2 _17299_ (.A(_04556_),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__a21oi_2 _17300_ (.A1(_04502_),
    .A2(_04528_),
    .B1(_04527_),
    .Y(_04559_));
 sky130_fd_sc_hd__xnor2_2 _17301_ (.A(_04558_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__nor2_2 _17302_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[6] ),
    .Y(_04561_));
 sky130_fd_sc_hd__a21oi_2 _17303_ (.A1(\systolic_inst.ce_local ),
    .A2(_04560_),
    .B1(_04561_),
    .Y(_01288_));
 sky130_fd_sc_hd__a21boi_2 _17304_ (.A1(_04530_),
    .A2(_04553_),
    .B1_N(_04552_),
    .Y(_04562_));
 sky130_fd_sc_hd__a21oi_2 _17305_ (.A1(_04507_),
    .A2(_04536_),
    .B1(_04535_),
    .Y(_04563_));
 sky130_fd_sc_hd__a22o_2 _17306_ (.A1(\systolic_inst.B_outs[10][1] ),
    .A2(\systolic_inst.A_outs[10][6] ),
    .B1(\systolic_inst.A_outs[10][7] ),
    .B2(\systolic_inst.B_outs[10][0] ),
    .X(_04564_));
 sky130_fd_sc_hd__nand4_2 _17307_ (.A(\systolic_inst.B_outs[10][0] ),
    .B(\systolic_inst.B_outs[10][1] ),
    .C(\systolic_inst.A_outs[10][6] ),
    .D(\systolic_inst.A_outs[10][7] ),
    .Y(_04565_));
 sky130_fd_sc_hd__and3_2 _17308_ (.A(\systolic_inst.B_outs[10][7] ),
    .B(_04564_),
    .C(_04565_),
    .X(_04566_));
 sky130_fd_sc_hd__a21oi_2 _17309_ (.A1(_04564_),
    .A2(_04565_),
    .B1(\systolic_inst.B_outs[10][7] ),
    .Y(_04567_));
 sky130_fd_sc_hd__a211o_2 _17310_ (.A1(_04538_),
    .A2(_04540_),
    .B1(_04566_),
    .C1(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__o211ai_2 _17311_ (.A1(_04566_),
    .A2(_04567_),
    .B1(_04538_),
    .C1(_04540_),
    .Y(_04569_));
 sky130_fd_sc_hd__and2_2 _17312_ (.A(_04568_),
    .B(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__xnor2_2 _17313_ (.A(_04533_),
    .B(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__nand2_2 _17314_ (.A(\systolic_inst.B_outs[10][2] ),
    .B(\systolic_inst.A_outs[10][5] ),
    .Y(_04572_));
 sky130_fd_sc_hd__and4_2 _17315_ (.A(\systolic_inst.B_outs[10][3] ),
    .B(\systolic_inst.A_outs[10][3] ),
    .C(\systolic_inst.B_outs[10][4] ),
    .D(\systolic_inst.A_outs[10][4] ),
    .X(_04573_));
 sky130_fd_sc_hd__a22oi_2 _17316_ (.A1(\systolic_inst.A_outs[10][3] ),
    .A2(\systolic_inst.B_outs[10][4] ),
    .B1(\systolic_inst.A_outs[10][4] ),
    .B2(\systolic_inst.B_outs[10][3] ),
    .Y(_04574_));
 sky130_fd_sc_hd__or2_2 _17317_ (.A(_04573_),
    .B(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__xnor2_2 _17318_ (.A(_04572_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__nand2_2 _17319_ (.A(\systolic_inst.A_outs[10][2] ),
    .B(\systolic_inst.B_outs[10][5] ),
    .Y(_04577_));
 sky130_fd_sc_hd__and2b_2 _17320_ (.A_N(\systolic_inst.A_outs[10][0] ),
    .B(\systolic_inst.B_outs[10][7] ),
    .X(_04578_));
 sky130_fd_sc_hd__and3_2 _17321_ (.A(\systolic_inst.A_outs[10][1] ),
    .B(\systolic_inst.B_outs[10][6] ),
    .C(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__xnor2_2 _17322_ (.A(_04543_),
    .B(_04578_),
    .Y(_04580_));
 sky130_fd_sc_hd__xnor2_2 _17323_ (.A(_04577_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__xnor2_2 _17324_ (.A(_04544_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_2 _17325_ (.A(_04576_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__xnor2_2 _17326_ (.A(_04576_),
    .B(_04582_),
    .Y(_04584_));
 sky130_fd_sc_hd__or2_2 _17327_ (.A(_04546_),
    .B(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__and2_2 _17328_ (.A(_04546_),
    .B(_04584_),
    .X(_04586_));
 sky130_fd_sc_hd__xor2_2 _17329_ (.A(_04546_),
    .B(_04584_),
    .X(_04587_));
 sky130_fd_sc_hd__xnor2_2 _17330_ (.A(_04571_),
    .B(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__and2b_2 _17331_ (.A_N(_04548_),
    .B(_04550_),
    .X(_04589_));
 sky130_fd_sc_hd__and2b_2 _17332_ (.A_N(_04589_),
    .B(_04588_),
    .X(_04590_));
 sky130_fd_sc_hd__xnor2_2 _17333_ (.A(_04588_),
    .B(_04589_),
    .Y(_04591_));
 sky130_fd_sc_hd__and2b_2 _17334_ (.A_N(_04563_),
    .B(_04591_),
    .X(_04592_));
 sky130_fd_sc_hd__xnor2_2 _17335_ (.A(_04563_),
    .B(_04591_),
    .Y(_04593_));
 sky130_fd_sc_hd__and2b_2 _17336_ (.A_N(_04562_),
    .B(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__xnor2_2 _17337_ (.A(_04562_),
    .B(_04593_),
    .Y(_04595_));
 sky130_fd_sc_hd__o21ai_2 _17338_ (.A1(_04558_),
    .A2(_04559_),
    .B1(_04556_),
    .Y(_04596_));
 sky130_fd_sc_hd__xor2_2 _17339_ (.A(_04595_),
    .B(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__mux2_1 _17340_ (.A0(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[7] ),
    .A1(_04597_),
    .S(\systolic_inst.ce_local ),
    .X(_01289_));
 sky130_fd_sc_hd__a21bo_2 _17341_ (.A1(_04533_),
    .A2(_04569_),
    .B1_N(_04568_),
    .X(_04598_));
 sky130_fd_sc_hd__a21bo_2 _17342_ (.A1(\systolic_inst.B_outs[10][7] ),
    .A2(_04564_),
    .B1_N(_04565_),
    .X(_04599_));
 sky130_fd_sc_hd__o21bai_2 _17343_ (.A1(_04572_),
    .A2(_04574_),
    .B1_N(_04573_),
    .Y(_04600_));
 sky130_fd_sc_hd__o21a_2 _17344_ (.A1(\systolic_inst.B_outs[10][0] ),
    .A2(\systolic_inst.B_outs[10][1] ),
    .B1(\systolic_inst.A_outs[10][7] ),
    .X(_04601_));
 sky130_fd_sc_hd__o21ai_2 _17345_ (.A1(\systolic_inst.B_outs[10][0] ),
    .A2(\systolic_inst.B_outs[10][1] ),
    .B1(\systolic_inst.A_outs[10][7] ),
    .Y(_04602_));
 sky130_fd_sc_hd__a21o_2 _17346_ (.A1(\systolic_inst.B_outs[10][0] ),
    .A2(\systolic_inst.B_outs[10][1] ),
    .B1(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__and2b_2 _17347_ (.A_N(_04603_),
    .B(_04600_),
    .X(_04604_));
 sky130_fd_sc_hd__xnor2_2 _17348_ (.A(_04600_),
    .B(_04603_),
    .Y(_04605_));
 sky130_fd_sc_hd__xnor2_2 _17349_ (.A(_04599_),
    .B(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__and4_2 _17350_ (.A(\systolic_inst.B_outs[10][3] ),
    .B(\systolic_inst.B_outs[10][4] ),
    .C(\systolic_inst.A_outs[10][4] ),
    .D(\systolic_inst.A_outs[10][5] ),
    .X(_04607_));
 sky130_fd_sc_hd__a22oi_2 _17351_ (.A1(\systolic_inst.B_outs[10][4] ),
    .A2(\systolic_inst.A_outs[10][4] ),
    .B1(\systolic_inst.A_outs[10][5] ),
    .B2(\systolic_inst.B_outs[10][3] ),
    .Y(_04608_));
 sky130_fd_sc_hd__nor2_2 _17352_ (.A(_04607_),
    .B(_04608_),
    .Y(_04609_));
 sky130_fd_sc_hd__nand2_2 _17353_ (.A(\systolic_inst.B_outs[10][2] ),
    .B(\systolic_inst.A_outs[10][6] ),
    .Y(_04610_));
 sky130_fd_sc_hd__xnor2_2 _17354_ (.A(_04609_),
    .B(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_2 _17355_ (.A(\systolic_inst.A_outs[10][3] ),
    .B(\systolic_inst.B_outs[10][5] ),
    .Y(_04612_));
 sky130_fd_sc_hd__and4b_2 _17356_ (.A_N(\systolic_inst.A_outs[10][1] ),
    .B(\systolic_inst.A_outs[10][2] ),
    .C(\systolic_inst.B_outs[10][6] ),
    .D(\systolic_inst.B_outs[10][7] ),
    .X(_04613_));
 sky130_fd_sc_hd__o2bb2a_2 _17357_ (.A1_N(\systolic_inst.A_outs[10][2] ),
    .A2_N(\systolic_inst.B_outs[10][6] ),
    .B1(_11275_),
    .B2(\systolic_inst.A_outs[10][1] ),
    .X(_04614_));
 sky130_fd_sc_hd__nor2_2 _17358_ (.A(_04613_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__xnor2_2 _17359_ (.A(_04612_),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__a31oi_2 _17360_ (.A1(\systolic_inst.A_outs[10][2] ),
    .A2(\systolic_inst.B_outs[10][5] ),
    .A3(_04580_),
    .B1(_04579_),
    .Y(_04617_));
 sky130_fd_sc_hd__nand2b_2 _17361_ (.A_N(_04617_),
    .B(_04616_),
    .Y(_04618_));
 sky130_fd_sc_hd__xnor2_2 _17362_ (.A(_04616_),
    .B(_04617_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_2 _17363_ (.A(_04611_),
    .B(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__xnor2_2 _17364_ (.A(_04611_),
    .B(_04619_),
    .Y(_04621_));
 sky130_fd_sc_hd__a21oi_2 _17365_ (.A1(_04544_),
    .A2(_04581_),
    .B1(_04583_),
    .Y(_04622_));
 sky130_fd_sc_hd__xnor2_2 _17366_ (.A(_04621_),
    .B(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__or2_2 _17367_ (.A(_04606_),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__xor2_2 _17368_ (.A(_04606_),
    .B(_04623_),
    .X(_04625_));
 sky130_fd_sc_hd__o21a_2 _17369_ (.A1(_04571_),
    .A2(_04586_),
    .B1(_04585_),
    .X(_04626_));
 sky130_fd_sc_hd__nand2b_2 _17370_ (.A_N(_04626_),
    .B(_04625_),
    .Y(_04627_));
 sky130_fd_sc_hd__xor2_2 _17371_ (.A(_04625_),
    .B(_04626_),
    .X(_04628_));
 sky130_fd_sc_hd__nand2b_2 _17372_ (.A_N(_04628_),
    .B(_04598_),
    .Y(_04629_));
 sky130_fd_sc_hd__xor2_2 _17373_ (.A(_04598_),
    .B(_04628_),
    .X(_04630_));
 sky130_fd_sc_hd__nor2_2 _17374_ (.A(_04590_),
    .B(_04592_),
    .Y(_04631_));
 sky130_fd_sc_hd__nor2_2 _17375_ (.A(_04630_),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__xor2_2 _17376_ (.A(_04630_),
    .B(_04631_),
    .X(_04633_));
 sky130_fd_sc_hd__a21oi_2 _17377_ (.A1(_04595_),
    .A2(_04596_),
    .B1(_04594_),
    .Y(_04634_));
 sky130_fd_sc_hd__and2b_2 _17378_ (.A_N(_04634_),
    .B(_04633_),
    .X(_04635_));
 sky130_fd_sc_hd__and2b_2 _17379_ (.A_N(_04633_),
    .B(_04634_),
    .X(_04636_));
 sky130_fd_sc_hd__nor2_2 _17380_ (.A(_04635_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__mux2_1 _17381_ (.A0(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[8] ),
    .A1(_04637_),
    .S(\systolic_inst.ce_local ),
    .X(_01290_));
 sky130_fd_sc_hd__a21o_2 _17382_ (.A1(_04599_),
    .A2(_04605_),
    .B1(_04604_),
    .X(_04638_));
 sky130_fd_sc_hd__o21ba_2 _17383_ (.A1(_04608_),
    .A2(_04610_),
    .B1_N(_04607_),
    .X(_04639_));
 sky130_fd_sc_hd__nor2_2 _17384_ (.A(_04602_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__and2_2 _17385_ (.A(_04602_),
    .B(_04639_),
    .X(_04641_));
 sky130_fd_sc_hd__or2_2 _17386_ (.A(_04640_),
    .B(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__nand2_2 _17387_ (.A(\systolic_inst.B_outs[10][2] ),
    .B(\systolic_inst.A_outs[10][7] ),
    .Y(_04643_));
 sky130_fd_sc_hd__a22oi_2 _17388_ (.A1(\systolic_inst.B_outs[10][4] ),
    .A2(\systolic_inst.A_outs[10][5] ),
    .B1(\systolic_inst.A_outs[10][6] ),
    .B2(\systolic_inst.B_outs[10][3] ),
    .Y(_04644_));
 sky130_fd_sc_hd__and4_2 _17389_ (.A(\systolic_inst.B_outs[10][3] ),
    .B(\systolic_inst.B_outs[10][4] ),
    .C(\systolic_inst.A_outs[10][5] ),
    .D(\systolic_inst.A_outs[10][6] ),
    .X(_04645_));
 sky130_fd_sc_hd__nor2_2 _17390_ (.A(_04644_),
    .B(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__xnor2_2 _17391_ (.A(_04643_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__nand2_2 _17392_ (.A(\systolic_inst.A_outs[10][4] ),
    .B(\systolic_inst.B_outs[10][5] ),
    .Y(_04648_));
 sky130_fd_sc_hd__and4b_2 _17393_ (.A_N(\systolic_inst.A_outs[10][2] ),
    .B(\systolic_inst.A_outs[10][3] ),
    .C(\systolic_inst.B_outs[10][6] ),
    .D(\systolic_inst.B_outs[10][7] ),
    .X(_04649_));
 sky130_fd_sc_hd__o2bb2a_2 _17394_ (.A1_N(\systolic_inst.A_outs[10][3] ),
    .A2_N(\systolic_inst.B_outs[10][6] ),
    .B1(_11275_),
    .B2(\systolic_inst.A_outs[10][2] ),
    .X(_04650_));
 sky130_fd_sc_hd__nor2_2 _17395_ (.A(_04649_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__xnor2_2 _17396_ (.A(_04648_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__o21ba_2 _17397_ (.A1(_04612_),
    .A2(_04614_),
    .B1_N(_04613_),
    .X(_04653_));
 sky130_fd_sc_hd__nand2b_2 _17398_ (.A_N(_04653_),
    .B(_04652_),
    .Y(_04654_));
 sky130_fd_sc_hd__xnor2_2 _17399_ (.A(_04652_),
    .B(_04653_),
    .Y(_04655_));
 sky130_fd_sc_hd__xnor2_2 _17400_ (.A(_04647_),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__a21o_2 _17401_ (.A1(_04618_),
    .A2(_04620_),
    .B1(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__nand3_2 _17402_ (.A(_04618_),
    .B(_04620_),
    .C(_04656_),
    .Y(_04658_));
 sky130_fd_sc_hd__nand2_2 _17403_ (.A(_04657_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__xor2_2 _17404_ (.A(_04642_),
    .B(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__o21a_2 _17405_ (.A1(_04621_),
    .A2(_04622_),
    .B1(_04624_),
    .X(_04661_));
 sky130_fd_sc_hd__nand2b_2 _17406_ (.A_N(_04661_),
    .B(_04660_),
    .Y(_04662_));
 sky130_fd_sc_hd__xnor2_2 _17407_ (.A(_04660_),
    .B(_04661_),
    .Y(_04663_));
 sky130_fd_sc_hd__xnor2_2 _17408_ (.A(_04638_),
    .B(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__a21o_2 _17409_ (.A1(_04627_),
    .A2(_04629_),
    .B1(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__nand3_2 _17410_ (.A(_04627_),
    .B(_04629_),
    .C(_04664_),
    .Y(_04666_));
 sky130_fd_sc_hd__nor2_2 _17411_ (.A(_04632_),
    .B(_04635_),
    .Y(_04667_));
 sky130_fd_sc_hd__a21oi_2 _17412_ (.A1(_04665_),
    .A2(_04666_),
    .B1(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__and3_2 _17413_ (.A(_04665_),
    .B(_04666_),
    .C(_04667_),
    .X(_04669_));
 sky130_fd_sc_hd__or2_2 _17414_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[9] ),
    .X(_04670_));
 sky130_fd_sc_hd__o31a_2 _17415_ (.A1(_11258_),
    .A2(_04668_),
    .A3(_04669_),
    .B1(_04670_),
    .X(_01291_));
 sky130_fd_sc_hd__o21ba_2 _17416_ (.A1(_04643_),
    .A2(_04644_),
    .B1_N(_04645_),
    .X(_04671_));
 sky130_fd_sc_hd__nor2_2 _17417_ (.A(_04602_),
    .B(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__and2_2 _17418_ (.A(_04602_),
    .B(_04671_),
    .X(_04673_));
 sky130_fd_sc_hd__or2_2 _17419_ (.A(_04672_),
    .B(_04673_),
    .X(_04674_));
 sky130_fd_sc_hd__a22o_2 _17420_ (.A1(\systolic_inst.B_outs[10][4] ),
    .A2(\systolic_inst.A_outs[10][6] ),
    .B1(\systolic_inst.A_outs[10][7] ),
    .B2(\systolic_inst.B_outs[10][3] ),
    .X(_04675_));
 sky130_fd_sc_hd__and3_2 _17421_ (.A(\systolic_inst.B_outs[10][3] ),
    .B(\systolic_inst.B_outs[10][4] ),
    .C(\systolic_inst.A_outs[10][7] ),
    .X(_04676_));
 sky130_fd_sc_hd__a21bo_2 _17422_ (.A1(\systolic_inst.A_outs[10][6] ),
    .A2(_04676_),
    .B1_N(_04675_),
    .X(_04677_));
 sky130_fd_sc_hd__xor2_2 _17423_ (.A(_04643_),
    .B(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__nand2_2 _17424_ (.A(\systolic_inst.B_outs[10][5] ),
    .B(\systolic_inst.A_outs[10][5] ),
    .Y(_04679_));
 sky130_fd_sc_hd__and4b_2 _17425_ (.A_N(\systolic_inst.A_outs[10][3] ),
    .B(\systolic_inst.A_outs[10][4] ),
    .C(\systolic_inst.B_outs[10][6] ),
    .D(\systolic_inst.B_outs[10][7] ),
    .X(_04680_));
 sky130_fd_sc_hd__o2bb2a_2 _17426_ (.A1_N(\systolic_inst.A_outs[10][4] ),
    .A2_N(\systolic_inst.B_outs[10][6] ),
    .B1(_11275_),
    .B2(\systolic_inst.A_outs[10][3] ),
    .X(_04681_));
 sky130_fd_sc_hd__nor2_2 _17427_ (.A(_04680_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__xnor2_2 _17428_ (.A(_04679_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__o21ba_2 _17429_ (.A1(_04648_),
    .A2(_04650_),
    .B1_N(_04649_),
    .X(_04684_));
 sky130_fd_sc_hd__nand2b_2 _17430_ (.A_N(_04684_),
    .B(_04683_),
    .Y(_04685_));
 sky130_fd_sc_hd__xnor2_2 _17431_ (.A(_04683_),
    .B(_04684_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand2_2 _17432_ (.A(_04678_),
    .B(_04686_),
    .Y(_04687_));
 sky130_fd_sc_hd__or2_2 _17433_ (.A(_04678_),
    .B(_04686_),
    .X(_04688_));
 sky130_fd_sc_hd__nand2_2 _17434_ (.A(_04687_),
    .B(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__a21bo_2 _17435_ (.A1(_04647_),
    .A2(_04655_),
    .B1_N(_04654_),
    .X(_04690_));
 sky130_fd_sc_hd__nand2b_2 _17436_ (.A_N(_04689_),
    .B(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__xor2_2 _17437_ (.A(_04689_),
    .B(_04690_),
    .X(_04692_));
 sky130_fd_sc_hd__xor2_2 _17438_ (.A(_04674_),
    .B(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__o21a_2 _17439_ (.A1(_04642_),
    .A2(_04659_),
    .B1(_04657_),
    .X(_04694_));
 sky130_fd_sc_hd__nand2b_2 _17440_ (.A_N(_04694_),
    .B(_04693_),
    .Y(_04695_));
 sky130_fd_sc_hd__xnor2_2 _17441_ (.A(_04693_),
    .B(_04694_),
    .Y(_04696_));
 sky130_fd_sc_hd__nand2_2 _17442_ (.A(_04640_),
    .B(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__or2_2 _17443_ (.A(_04640_),
    .B(_04696_),
    .X(_04698_));
 sky130_fd_sc_hd__nand2_2 _17444_ (.A(_04697_),
    .B(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__a21boi_2 _17445_ (.A1(_04638_),
    .A2(_04663_),
    .B1_N(_04662_),
    .Y(_04700_));
 sky130_fd_sc_hd__nor2_2 _17446_ (.A(_04699_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__xnor2_2 _17447_ (.A(_04699_),
    .B(_04700_),
    .Y(_04702_));
 sky130_fd_sc_hd__o21ai_2 _17448_ (.A1(_04632_),
    .A2(_04635_),
    .B1(_04666_),
    .Y(_04703_));
 sky130_fd_sc_hd__and3_2 _17449_ (.A(_04665_),
    .B(_04702_),
    .C(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__a21oi_2 _17450_ (.A1(_04665_),
    .A2(_04703_),
    .B1(_04702_),
    .Y(_04705_));
 sky130_fd_sc_hd__or3_2 _17451_ (.A(_11258_),
    .B(_04704_),
    .C(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__a21bo_2 _17452_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[10] ),
    .B1_N(_04706_),
    .X(_01292_));
 sky130_fd_sc_hd__or2_2 _17453_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[11] ),
    .X(_04707_));
 sky130_fd_sc_hd__o2bb2a_2 _17454_ (.A1_N(\systolic_inst.A_outs[10][6] ),
    .A2_N(_04676_),
    .B1(_04677_),
    .B2(_04643_),
    .X(_04708_));
 sky130_fd_sc_hd__or2_2 _17455_ (.A(_04602_),
    .B(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__nand2_2 _17456_ (.A(_04602_),
    .B(_04708_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_2 _17457_ (.A(_04709_),
    .B(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__or2_2 _17458_ (.A(\systolic_inst.B_outs[10][3] ),
    .B(\systolic_inst.B_outs[10][4] ),
    .X(_04712_));
 sky130_fd_sc_hd__and3b_2 _17459_ (.A_N(_04676_),
    .B(_04712_),
    .C(\systolic_inst.A_outs[10][7] ),
    .X(_04713_));
 sky130_fd_sc_hd__xnor2_2 _17460_ (.A(_04643_),
    .B(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__nand2_2 _17461_ (.A(\systolic_inst.B_outs[10][5] ),
    .B(\systolic_inst.A_outs[10][6] ),
    .Y(_04715_));
 sky130_fd_sc_hd__and4b_2 _17462_ (.A_N(\systolic_inst.A_outs[10][4] ),
    .B(\systolic_inst.A_outs[10][5] ),
    .C(\systolic_inst.B_outs[10][6] ),
    .D(\systolic_inst.B_outs[10][7] ),
    .X(_04716_));
 sky130_fd_sc_hd__o2bb2a_2 _17463_ (.A1_N(\systolic_inst.A_outs[10][5] ),
    .A2_N(\systolic_inst.B_outs[10][6] ),
    .B1(_11275_),
    .B2(\systolic_inst.A_outs[10][4] ),
    .X(_04717_));
 sky130_fd_sc_hd__or2_2 _17464_ (.A(_04716_),
    .B(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__xor2_2 _17465_ (.A(_04715_),
    .B(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__o21ba_2 _17466_ (.A1(_04679_),
    .A2(_04681_),
    .B1_N(_04680_),
    .X(_04720_));
 sky130_fd_sc_hd__nand2b_2 _17467_ (.A_N(_04720_),
    .B(_04719_),
    .Y(_04721_));
 sky130_fd_sc_hd__xnor2_2 _17468_ (.A(_04719_),
    .B(_04720_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_2 _17469_ (.A(_04714_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__xnor2_2 _17470_ (.A(_04714_),
    .B(_04722_),
    .Y(_04724_));
 sky130_fd_sc_hd__a21o_2 _17471_ (.A1(_04685_),
    .A2(_04687_),
    .B1(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__nand3_2 _17472_ (.A(_04685_),
    .B(_04687_),
    .C(_04724_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2_2 _17473_ (.A(_04725_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__xor2_2 _17474_ (.A(_04711_),
    .B(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__o21a_2 _17475_ (.A1(_04674_),
    .A2(_04692_),
    .B1(_04691_),
    .X(_04729_));
 sky130_fd_sc_hd__and2b_2 _17476_ (.A_N(_04729_),
    .B(_04728_),
    .X(_04730_));
 sky130_fd_sc_hd__xnor2_2 _17477_ (.A(_04728_),
    .B(_04729_),
    .Y(_04731_));
 sky130_fd_sc_hd__xnor2_2 _17478_ (.A(_04672_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__and3_2 _17479_ (.A(_04695_),
    .B(_04697_),
    .C(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__inv_2 _17480_ (.A(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__a21oi_2 _17481_ (.A1(_04695_),
    .A2(_04697_),
    .B1(_04732_),
    .Y(_04735_));
 sky130_fd_sc_hd__nor4_2 _17482_ (.A(_04701_),
    .B(_04705_),
    .C(_04733_),
    .D(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__o22a_2 _17483_ (.A1(_04701_),
    .A2(_04705_),
    .B1(_04733_),
    .B2(_04735_),
    .X(_04737_));
 sky130_fd_sc_hd__o31a_2 _17484_ (.A1(_11258_),
    .A2(_04736_),
    .A3(_04737_),
    .B1(_04707_),
    .X(_01293_));
 sky130_fd_sc_hd__a31o_2 _17485_ (.A1(\systolic_inst.B_outs[10][2] ),
    .A2(\systolic_inst.A_outs[10][7] ),
    .A3(_04712_),
    .B1(_04676_),
    .X(_04738_));
 sky130_fd_sc_hd__or2_2 _17486_ (.A(_04601_),
    .B(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__nand2_2 _17487_ (.A(_04601_),
    .B(_04738_),
    .Y(_04740_));
 sky130_fd_sc_hd__nand2_2 _17488_ (.A(_04739_),
    .B(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__inv_2 _17489_ (.A(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__o2bb2a_2 _17490_ (.A1_N(\systolic_inst.B_outs[10][6] ),
    .A2_N(\systolic_inst.A_outs[10][6] ),
    .B1(_11275_),
    .B2(\systolic_inst.A_outs[10][5] ),
    .X(_04743_));
 sky130_fd_sc_hd__and4b_2 _17491_ (.A_N(\systolic_inst.A_outs[10][5] ),
    .B(\systolic_inst.B_outs[10][6] ),
    .C(\systolic_inst.A_outs[10][6] ),
    .D(\systolic_inst.B_outs[10][7] ),
    .X(_04744_));
 sky130_fd_sc_hd__nor2_2 _17492_ (.A(_04743_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2_2 _17493_ (.A(\systolic_inst.B_outs[10][5] ),
    .B(\systolic_inst.A_outs[10][7] ),
    .Y(_04746_));
 sky130_fd_sc_hd__and3_2 _17494_ (.A(\systolic_inst.B_outs[10][5] ),
    .B(\systolic_inst.A_outs[10][7] ),
    .C(_04745_),
    .X(_04747_));
 sky130_fd_sc_hd__xnor2_2 _17495_ (.A(_04745_),
    .B(_04746_),
    .Y(_04748_));
 sky130_fd_sc_hd__o21ba_2 _17496_ (.A1(_04715_),
    .A2(_04717_),
    .B1_N(_04716_),
    .X(_04749_));
 sky130_fd_sc_hd__nand2b_2 _17497_ (.A_N(_04749_),
    .B(_04748_),
    .Y(_04750_));
 sky130_fd_sc_hd__xnor2_2 _17498_ (.A(_04748_),
    .B(_04749_),
    .Y(_04751_));
 sky130_fd_sc_hd__xnor2_2 _17499_ (.A(_04714_),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__a21o_2 _17500_ (.A1(_04721_),
    .A2(_04723_),
    .B1(_04752_),
    .X(_04753_));
 sky130_fd_sc_hd__nand3_2 _17501_ (.A(_04721_),
    .B(_04723_),
    .C(_04752_),
    .Y(_04754_));
 sky130_fd_sc_hd__nand2_2 _17502_ (.A(_04753_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__xnor2_2 _17503_ (.A(_04742_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__o21a_2 _17504_ (.A1(_04711_),
    .A2(_04727_),
    .B1(_04725_),
    .X(_04757_));
 sky130_fd_sc_hd__and2b_2 _17505_ (.A_N(_04757_),
    .B(_04756_),
    .X(_04758_));
 sky130_fd_sc_hd__xnor2_2 _17506_ (.A(_04756_),
    .B(_04757_),
    .Y(_04759_));
 sky130_fd_sc_hd__and2b_2 _17507_ (.A_N(_04709_),
    .B(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__xor2_2 _17508_ (.A(_04709_),
    .B(_04759_),
    .X(_04761_));
 sky130_fd_sc_hd__a21oi_2 _17509_ (.A1(_04672_),
    .A2(_04731_),
    .B1(_04730_),
    .Y(_04762_));
 sky130_fd_sc_hd__nor2_2 _17510_ (.A(_04761_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__and2_2 _17511_ (.A(_04761_),
    .B(_04762_),
    .X(_04764_));
 sky130_fd_sc_hd__or2_2 _17512_ (.A(_04763_),
    .B(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__inv_2 _17513_ (.A(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__o31a_2 _17514_ (.A1(_04701_),
    .A2(_04705_),
    .A3(_04735_),
    .B1(_04734_),
    .X(_04767_));
 sky130_fd_sc_hd__o311a_2 _17515_ (.A1(_04701_),
    .A2(_04705_),
    .A3(_04735_),
    .B1(_04766_),
    .C1(_04734_),
    .X(_04768_));
 sky130_fd_sc_hd__nor2_2 _17516_ (.A(_04766_),
    .B(_04767_),
    .Y(_04769_));
 sky130_fd_sc_hd__nor2_2 _17517_ (.A(_04768_),
    .B(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__mux2_1 _17518_ (.A0(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[12] ),
    .A1(_04770_),
    .S(\systolic_inst.ce_local ),
    .X(_01294_));
 sky130_fd_sc_hd__nand2_2 _17519_ (.A(\systolic_inst.B_outs[10][6] ),
    .B(\systolic_inst.A_outs[10][7] ),
    .Y(_04771_));
 sky130_fd_sc_hd__nor2_2 _17520_ (.A(\systolic_inst.A_outs[10][6] ),
    .B(_11275_),
    .Y(_04772_));
 sky130_fd_sc_hd__xnor2_2 _17521_ (.A(_04771_),
    .B(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__nand2b_2 _17522_ (.A_N(_04746_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__xnor2_2 _17523_ (.A(_04746_),
    .B(_04773_),
    .Y(_04775_));
 sky130_fd_sc_hd__o21ai_2 _17524_ (.A1(_04744_),
    .A2(_04747_),
    .B1(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__or3_2 _17525_ (.A(_04744_),
    .B(_04747_),
    .C(_04775_),
    .X(_04777_));
 sky130_fd_sc_hd__and2_2 _17526_ (.A(_04776_),
    .B(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__nand2_2 _17527_ (.A(_04714_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__or2_2 _17528_ (.A(_04714_),
    .B(_04778_),
    .X(_04780_));
 sky130_fd_sc_hd__nand2_2 _17529_ (.A(_04779_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__a21bo_2 _17530_ (.A1(_04714_),
    .A2(_04751_),
    .B1_N(_04750_),
    .X(_04782_));
 sky130_fd_sc_hd__nand2b_2 _17531_ (.A_N(_04781_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__xor2_2 _17532_ (.A(_04781_),
    .B(_04782_),
    .X(_04784_));
 sky130_fd_sc_hd__xnor2_2 _17533_ (.A(_04742_),
    .B(_04784_),
    .Y(_04785_));
 sky130_fd_sc_hd__o21a_2 _17534_ (.A1(_04741_),
    .A2(_04755_),
    .B1(_04753_),
    .X(_04786_));
 sky130_fd_sc_hd__and2b_2 _17535_ (.A_N(_04786_),
    .B(_04785_),
    .X(_04787_));
 sky130_fd_sc_hd__and2b_2 _17536_ (.A_N(_04785_),
    .B(_04786_),
    .X(_04788_));
 sky130_fd_sc_hd__nor2_2 _17537_ (.A(_04787_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__xnor2_2 _17538_ (.A(_04740_),
    .B(_04789_),
    .Y(_04790_));
 sky130_fd_sc_hd__nor3_2 _17539_ (.A(_04758_),
    .B(_04760_),
    .C(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__o21a_2 _17540_ (.A1(_04758_),
    .A2(_04760_),
    .B1(_04790_),
    .X(_04792_));
 sky130_fd_sc_hd__nor2_2 _17541_ (.A(_04791_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__o21ai_2 _17542_ (.A1(_04763_),
    .A2(_04768_),
    .B1(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__o31a_2 _17543_ (.A1(_04763_),
    .A2(_04768_),
    .A3(_04793_),
    .B1(\systolic_inst.ce_local ),
    .X(_04795_));
 sky130_fd_sc_hd__a22o_2 _17544_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[13] ),
    .B1(_04794_),
    .B2(_04795_),
    .X(_01295_));
 sky130_fd_sc_hd__o211ai_2 _17545_ (.A1(_11275_),
    .A2(\systolic_inst.A_outs[10][7] ),
    .B1(_04746_),
    .C1(_04771_),
    .Y(_04796_));
 sky130_fd_sc_hd__o311a_2 _17546_ (.A1(\systolic_inst.A_outs[10][6] ),
    .A2(_11275_),
    .A3(_04771_),
    .B1(_04774_),
    .C1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__a31o_2 _17547_ (.A1(\systolic_inst.B_outs[10][5] ),
    .A2(\systolic_inst.B_outs[10][6] ),
    .A3(\systolic_inst.A_outs[10][7] ),
    .B1(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__or2_2 _17548_ (.A(_04714_),
    .B(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__nand2_2 _17549_ (.A(_04714_),
    .B(_04798_),
    .Y(_04800_));
 sky130_fd_sc_hd__nand2_2 _17550_ (.A(_04799_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__a21oi_2 _17551_ (.A1(_04776_),
    .A2(_04779_),
    .B1(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__and3_2 _17552_ (.A(_04776_),
    .B(_04779_),
    .C(_04801_),
    .X(_04803_));
 sky130_fd_sc_hd__nor2_2 _17553_ (.A(_04802_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__xnor2_2 _17554_ (.A(_04741_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__o21a_2 _17555_ (.A1(_04741_),
    .A2(_04784_),
    .B1(_04783_),
    .X(_04806_));
 sky130_fd_sc_hd__and2b_2 _17556_ (.A_N(_04806_),
    .B(_04805_),
    .X(_04807_));
 sky130_fd_sc_hd__and2b_2 _17557_ (.A_N(_04805_),
    .B(_04806_),
    .X(_04808_));
 sky130_fd_sc_hd__nor2_2 _17558_ (.A(_04807_),
    .B(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__xnor2_2 _17559_ (.A(_04740_),
    .B(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__o21ba_2 _17560_ (.A1(_04740_),
    .A2(_04788_),
    .B1_N(_04787_),
    .X(_04811_));
 sky130_fd_sc_hd__nand2b_2 _17561_ (.A_N(_04811_),
    .B(_04810_),
    .Y(_04812_));
 sky130_fd_sc_hd__xnor2_2 _17562_ (.A(_04810_),
    .B(_04811_),
    .Y(_04813_));
 sky130_fd_sc_hd__nor2_2 _17563_ (.A(_04763_),
    .B(_04792_),
    .Y(_04814_));
 sky130_fd_sc_hd__a2bb2o_2 _17564_ (.A1_N(_04791_),
    .A2_N(_04814_),
    .B1(_04793_),
    .B2(_04768_),
    .X(_04815_));
 sky130_fd_sc_hd__nand2_2 _17565_ (.A(_04813_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__xor2_2 _17566_ (.A(_04813_),
    .B(_04815_),
    .X(_04817_));
 sky130_fd_sc_hd__mux2_1 _17567_ (.A0(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[14] ),
    .A1(_04817_),
    .S(\systolic_inst.ce_local ),
    .X(_01296_));
 sky130_fd_sc_hd__a31o_2 _17568_ (.A1(_04601_),
    .A2(_04738_),
    .A3(_04809_),
    .B1(_04807_),
    .X(_04818_));
 sky130_fd_sc_hd__a21oi_2 _17569_ (.A1(_04742_),
    .A2(_04804_),
    .B1(_04802_),
    .Y(_04819_));
 sky130_fd_sc_hd__xnor2_2 _17570_ (.A(_04739_),
    .B(_04799_),
    .Y(_04820_));
 sky130_fd_sc_hd__xnor2_2 _17571_ (.A(_04819_),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__xnor2_2 _17572_ (.A(_04818_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__and3_2 _17573_ (.A(\systolic_inst.ce_local ),
    .B(_04812_),
    .C(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__a22o_2 _17574_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B1(_04816_),
    .B2(_04823_),
    .X(_01297_));
 sky130_fd_sc_hd__a21o_2 _17575_ (.A1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[10][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_04824_));
 sky130_fd_sc_hd__a21oi_2 _17576_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[10][0] ),
    .Y(_04825_));
 sky130_fd_sc_hd__a21oi_2 _17577_ (.A1(\systolic_inst.ce_local ),
    .A2(_04824_),
    .B1(_04825_),
    .Y(_01298_));
 sky130_fd_sc_hd__and2_2 _17578_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[10][1] ),
    .X(_04826_));
 sky130_fd_sc_hd__nand2_2 _17579_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[10][1] ),
    .Y(_04827_));
 sky130_fd_sc_hd__or2_2 _17580_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[10][1] ),
    .X(_04828_));
 sky130_fd_sc_hd__and4_2 _17581_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[10][0] ),
    .C(_04827_),
    .D(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__inv_2 _17582_ (.A(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__a22o_2 _17583_ (.A1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[10][0] ),
    .B1(_04827_),
    .B2(_04828_),
    .X(_04831_));
 sky130_fd_sc_hd__a32o_2 _17584_ (.A1(_11712_),
    .A2(_04830_),
    .A3(_04831_),
    .B1(\systolic_inst.acc_wires[10][1] ),
    .B2(_11258_),
    .X(_01299_));
 sky130_fd_sc_hd__nand2_2 _17585_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[10][2] ),
    .Y(_04832_));
 sky130_fd_sc_hd__or2_2 _17586_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[10][2] ),
    .X(_04833_));
 sky130_fd_sc_hd__a31o_2 _17587_ (.A1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[10][0] ),
    .A3(_04828_),
    .B1(_04826_),
    .X(_04834_));
 sky130_fd_sc_hd__a21o_2 _17588_ (.A1(_04832_),
    .A2(_04833_),
    .B1(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__and3_2 _17589_ (.A(_04832_),
    .B(_04833_),
    .C(_04834_),
    .X(_04836_));
 sky130_fd_sc_hd__inv_2 _17590_ (.A(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__a32o_2 _17591_ (.A1(_11712_),
    .A2(_04835_),
    .A3(_04837_),
    .B1(\systolic_inst.acc_wires[10][2] ),
    .B2(_11258_),
    .X(_01300_));
 sky130_fd_sc_hd__nand2_2 _17592_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[10][3] ),
    .Y(_04838_));
 sky130_fd_sc_hd__or2_2 _17593_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[10][3] ),
    .X(_04839_));
 sky130_fd_sc_hd__a21bo_2 _17594_ (.A1(_04833_),
    .A2(_04834_),
    .B1_N(_04832_),
    .X(_04840_));
 sky130_fd_sc_hd__a21o_2 _17595_ (.A1(_04838_),
    .A2(_04839_),
    .B1(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__and3_2 _17596_ (.A(_04838_),
    .B(_04839_),
    .C(_04840_),
    .X(_04842_));
 sky130_fd_sc_hd__inv_2 _17597_ (.A(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__a32o_2 _17598_ (.A1(_11712_),
    .A2(_04841_),
    .A3(_04843_),
    .B1(\systolic_inst.acc_wires[10][3] ),
    .B2(_11258_),
    .X(_01301_));
 sky130_fd_sc_hd__nand2_2 _17599_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[10][4] ),
    .Y(_04844_));
 sky130_fd_sc_hd__or2_2 _17600_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[10][4] ),
    .X(_04845_));
 sky130_fd_sc_hd__a21bo_2 _17601_ (.A1(_04839_),
    .A2(_04840_),
    .B1_N(_04838_),
    .X(_04846_));
 sky130_fd_sc_hd__and3_2 _17602_ (.A(_04844_),
    .B(_04845_),
    .C(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__inv_2 _17603_ (.A(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__a21o_2 _17604_ (.A1(_04844_),
    .A2(_04845_),
    .B1(_04846_),
    .X(_04849_));
 sky130_fd_sc_hd__a32o_2 _17605_ (.A1(_11712_),
    .A2(_04848_),
    .A3(_04849_),
    .B1(\systolic_inst.acc_wires[10][4] ),
    .B2(_11258_),
    .X(_01302_));
 sky130_fd_sc_hd__nand2_2 _17606_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[10][5] ),
    .Y(_04850_));
 sky130_fd_sc_hd__or2_2 _17607_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[10][5] ),
    .X(_04851_));
 sky130_fd_sc_hd__a21bo_2 _17608_ (.A1(_04845_),
    .A2(_04846_),
    .B1_N(_04844_),
    .X(_04852_));
 sky130_fd_sc_hd__a21o_2 _17609_ (.A1(_04850_),
    .A2(_04851_),
    .B1(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__and3_2 _17610_ (.A(_04850_),
    .B(_04851_),
    .C(_04852_),
    .X(_04854_));
 sky130_fd_sc_hd__inv_2 _17611_ (.A(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__a32o_2 _17612_ (.A1(_11712_),
    .A2(_04853_),
    .A3(_04855_),
    .B1(\systolic_inst.acc_wires[10][5] ),
    .B2(_11258_),
    .X(_01303_));
 sky130_fd_sc_hd__nand2_2 _17613_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[10][6] ),
    .Y(_04856_));
 sky130_fd_sc_hd__or2_2 _17614_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[10][6] ),
    .X(_04857_));
 sky130_fd_sc_hd__a21bo_2 _17615_ (.A1(_04851_),
    .A2(_04852_),
    .B1_N(_04850_),
    .X(_04858_));
 sky130_fd_sc_hd__a21o_2 _17616_ (.A1(_04856_),
    .A2(_04857_),
    .B1(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__and3_2 _17617_ (.A(_04856_),
    .B(_04857_),
    .C(_04858_),
    .X(_04860_));
 sky130_fd_sc_hd__inv_2 _17618_ (.A(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__a32o_2 _17619_ (.A1(_11712_),
    .A2(_04859_),
    .A3(_04861_),
    .B1(\systolic_inst.acc_wires[10][6] ),
    .B2(_11258_),
    .X(_01304_));
 sky130_fd_sc_hd__nand2_2 _17620_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[10][7] ),
    .Y(_04862_));
 sky130_fd_sc_hd__or2_2 _17621_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[10][7] ),
    .X(_04863_));
 sky130_fd_sc_hd__a21bo_2 _17622_ (.A1(_04857_),
    .A2(_04858_),
    .B1_N(_04856_),
    .X(_04864_));
 sky130_fd_sc_hd__nand3_2 _17623_ (.A(_04862_),
    .B(_04863_),
    .C(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__a21o_2 _17624_ (.A1(_04862_),
    .A2(_04863_),
    .B1(_04864_),
    .X(_04866_));
 sky130_fd_sc_hd__a32o_2 _17625_ (.A1(_11712_),
    .A2(_04865_),
    .A3(_04866_),
    .B1(\systolic_inst.acc_wires[10][7] ),
    .B2(_11258_),
    .X(_01305_));
 sky130_fd_sc_hd__a21bo_2 _17626_ (.A1(_04863_),
    .A2(_04864_),
    .B1_N(_04862_),
    .X(_04867_));
 sky130_fd_sc_hd__xnor2_2 _17627_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[10][8] ),
    .Y(_04868_));
 sky130_fd_sc_hd__and2b_2 _17628_ (.A_N(_04868_),
    .B(_04867_),
    .X(_04869_));
 sky130_fd_sc_hd__a31o_2 _17629_ (.A1(_04862_),
    .A2(_04865_),
    .A3(_04868_),
    .B1(_11713_),
    .X(_04870_));
 sky130_fd_sc_hd__a2bb2o_2 _17630_ (.A1_N(_04870_),
    .A2_N(_04869_),
    .B1(\systolic_inst.acc_wires[10][8] ),
    .B2(_11258_),
    .X(_01306_));
 sky130_fd_sc_hd__xor2_2 _17631_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[10][9] ),
    .X(_04871_));
 sky130_fd_sc_hd__a211o_2 _17632_ (.A1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[10][8] ),
    .B1(_04869_),
    .C1(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__nand2_2 _17633_ (.A(_04869_),
    .B(_04871_),
    .Y(_04873_));
 sky130_fd_sc_hd__and3_2 _17634_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[10][8] ),
    .C(_04871_),
    .X(_04874_));
 sky130_fd_sc_hd__nor2_2 _17635_ (.A(_11713_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__a32o_2 _17636_ (.A1(_04872_),
    .A2(_04873_),
    .A3(_04875_),
    .B1(\systolic_inst.acc_wires[10][9] ),
    .B2(_11258_),
    .X(_01307_));
 sky130_fd_sc_hd__nand2_2 _17637_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[10][10] ),
    .Y(_04876_));
 sky130_fd_sc_hd__or2_2 _17638_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[10][10] ),
    .X(_04877_));
 sky130_fd_sc_hd__and2_2 _17639_ (.A(_04876_),
    .B(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__a21oi_2 _17640_ (.A1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[10][9] ),
    .B1(_04874_),
    .Y(_04879_));
 sky130_fd_sc_hd__nand2_2 _17641_ (.A(_04873_),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_2 _17642_ (.A(_04878_),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__or2_2 _17643_ (.A(_04878_),
    .B(_04880_),
    .X(_04882_));
 sky130_fd_sc_hd__a32o_2 _17644_ (.A1(_11712_),
    .A2(_04881_),
    .A3(_04882_),
    .B1(\systolic_inst.acc_wires[10][10] ),
    .B2(_11258_),
    .X(_01308_));
 sky130_fd_sc_hd__nor2_2 _17645_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[10][11] ),
    .Y(_04883_));
 sky130_fd_sc_hd__or2_2 _17646_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[10][11] ),
    .X(_04884_));
 sky130_fd_sc_hd__nand2_2 _17647_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[10][11] ),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_2 _17648_ (.A(_04884_),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__a21oi_2 _17649_ (.A1(_04876_),
    .A2(_04881_),
    .B1(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__a31o_2 _17650_ (.A1(_04876_),
    .A2(_04881_),
    .A3(_04886_),
    .B1(_11713_),
    .X(_04888_));
 sky130_fd_sc_hd__a2bb2o_2 _17651_ (.A1_N(_04888_),
    .A2_N(_04887_),
    .B1(\systolic_inst.acc_wires[10][11] ),
    .B2(_11258_),
    .X(_01309_));
 sky130_fd_sc_hd__nand3_2 _17652_ (.A(_04878_),
    .B(_04884_),
    .C(_04885_),
    .Y(_04889_));
 sky130_fd_sc_hd__inv_2 _17653_ (.A(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__and3b_2 _17654_ (.A_N(_04868_),
    .B(_04871_),
    .C(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__o2bb2a_2 _17655_ (.A1_N(_04867_),
    .A2_N(_04891_),
    .B1(_04879_),
    .B2(_04889_),
    .X(_04892_));
 sky130_fd_sc_hd__o21a_2 _17656_ (.A1(_04876_),
    .A2(_04883_),
    .B1(_04885_),
    .X(_04893_));
 sky130_fd_sc_hd__xnor2_2 _17657_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[10][12] ),
    .Y(_04894_));
 sky130_fd_sc_hd__and3_2 _17658_ (.A(_04892_),
    .B(_04893_),
    .C(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__a21oi_2 _17659_ (.A1(_04892_),
    .A2(_04893_),
    .B1(_04894_),
    .Y(_04896_));
 sky130_fd_sc_hd__nor2_2 _17660_ (.A(_04895_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__a22o_2 _17661_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][12] ),
    .B1(_11712_),
    .B2(_04897_),
    .X(_01310_));
 sky130_fd_sc_hd__xor2_2 _17662_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[10][13] ),
    .X(_04898_));
 sky130_fd_sc_hd__a211o_2 _17663_ (.A1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[10][12] ),
    .B1(_04896_),
    .C1(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__nand2b_2 _17664_ (.A_N(_04894_),
    .B(_04898_),
    .Y(_04900_));
 sky130_fd_sc_hd__a21o_2 _17665_ (.A1(_04892_),
    .A2(_04893_),
    .B1(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__and3_2 _17666_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[10][12] ),
    .C(_04898_),
    .X(_04902_));
 sky130_fd_sc_hd__nor2_2 _17667_ (.A(_11713_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__a32o_2 _17668_ (.A1(_04899_),
    .A2(_04901_),
    .A3(_04903_),
    .B1(\systolic_inst.acc_wires[10][13] ),
    .B2(_11258_),
    .X(_01311_));
 sky130_fd_sc_hd__or2_2 _17669_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[10][14] ),
    .X(_04904_));
 sky130_fd_sc_hd__nand2_2 _17670_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[10][14] ),
    .Y(_04905_));
 sky130_fd_sc_hd__and2_2 _17671_ (.A(_04904_),
    .B(_04905_),
    .X(_04906_));
 sky130_fd_sc_hd__nand2_2 _17672_ (.A(_04904_),
    .B(_04905_),
    .Y(_04907_));
 sky130_fd_sc_hd__a21oi_2 _17673_ (.A1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[10][13] ),
    .B1(_04902_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand2_2 _17674_ (.A(_04901_),
    .B(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__nand2_2 _17675_ (.A(_04906_),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__or2_2 _17676_ (.A(_04906_),
    .B(_04909_),
    .X(_04911_));
 sky130_fd_sc_hd__a32o_2 _17677_ (.A1(_11712_),
    .A2(_04910_),
    .A3(_04911_),
    .B1(\systolic_inst.acc_wires[10][14] ),
    .B2(_11258_),
    .X(_01312_));
 sky130_fd_sc_hd__nor2_2 _17678_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][15] ),
    .Y(_04912_));
 sky130_fd_sc_hd__and2_2 _17679_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][15] ),
    .X(_04913_));
 sky130_fd_sc_hd__or2_2 _17680_ (.A(_04912_),
    .B(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__a21oi_2 _17681_ (.A1(_04905_),
    .A2(_04910_),
    .B1(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__a31o_2 _17682_ (.A1(_04905_),
    .A2(_04910_),
    .A3(_04914_),
    .B1(_11713_),
    .X(_04916_));
 sky130_fd_sc_hd__a2bb2o_2 _17683_ (.A1_N(_04916_),
    .A2_N(_04915_),
    .B1(\systolic_inst.acc_wires[10][15] ),
    .B2(_11258_),
    .X(_01313_));
 sky130_fd_sc_hd__a211o_2 _17684_ (.A1(_04901_),
    .A2(_04908_),
    .B1(_04914_),
    .C1(_04907_),
    .X(_04917_));
 sky130_fd_sc_hd__o21ba_2 _17685_ (.A1(_04905_),
    .A2(_04912_),
    .B1_N(_04913_),
    .X(_04918_));
 sky130_fd_sc_hd__and2_2 _17686_ (.A(_04917_),
    .B(_04918_),
    .X(_04919_));
 sky130_fd_sc_hd__xnor2_2 _17687_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][16] ),
    .Y(_04920_));
 sky130_fd_sc_hd__nand2_2 _17688_ (.A(_04919_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__nor2_2 _17689_ (.A(_04919_),
    .B(_04920_),
    .Y(_04922_));
 sky130_fd_sc_hd__nor2_2 _17690_ (.A(_11713_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__a22o_2 _17691_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][16] ),
    .B1(_04921_),
    .B2(_04923_),
    .X(_01314_));
 sky130_fd_sc_hd__xor2_2 _17692_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][17] ),
    .X(_04924_));
 sky130_fd_sc_hd__inv_2 _17693_ (.A(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__a21oi_2 _17694_ (.A1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[10][16] ),
    .B1(_04922_),
    .Y(_04926_));
 sky130_fd_sc_hd__xnor2_2 _17695_ (.A(_04924_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__a22o_2 _17696_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][17] ),
    .B1(_11712_),
    .B2(_04927_),
    .X(_01315_));
 sky130_fd_sc_hd__or2_2 _17697_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][18] ),
    .X(_04928_));
 sky130_fd_sc_hd__nand2_2 _17698_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][18] ),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_2 _17699_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__o21a_2 _17700_ (.A1(\systolic_inst.acc_wires[10][16] ),
    .A2(\systolic_inst.acc_wires[10][17] ),
    .B1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .X(_04931_));
 sky130_fd_sc_hd__a21oi_2 _17701_ (.A1(_04922_),
    .A2(_04924_),
    .B1(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__xor2_2 _17702_ (.A(_04930_),
    .B(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__a22o_2 _17703_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][18] ),
    .B1(_11712_),
    .B2(_04933_),
    .X(_01316_));
 sky130_fd_sc_hd__xnor2_2 _17704_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][19] ),
    .Y(_04934_));
 sky130_fd_sc_hd__o21ai_2 _17705_ (.A1(_04930_),
    .A2(_04932_),
    .B1(_04929_),
    .Y(_04935_));
 sky130_fd_sc_hd__xnor2_2 _17706_ (.A(_04934_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__a22o_2 _17707_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][19] ),
    .B1(_11712_),
    .B2(_04936_),
    .X(_01317_));
 sky130_fd_sc_hd__or2_2 _17708_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][20] ),
    .X(_04937_));
 sky130_fd_sc_hd__nand2_2 _17709_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][20] ),
    .Y(_04938_));
 sky130_fd_sc_hd__and2_2 _17710_ (.A(_04937_),
    .B(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__or4_2 _17711_ (.A(_04920_),
    .B(_04925_),
    .C(_04930_),
    .D(_04934_),
    .X(_04940_));
 sky130_fd_sc_hd__nor2_2 _17712_ (.A(_04919_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__o41a_2 _17713_ (.A1(\systolic_inst.acc_wires[10][16] ),
    .A2(\systolic_inst.acc_wires[10][17] ),
    .A3(\systolic_inst.acc_wires[10][18] ),
    .A4(\systolic_inst.acc_wires[10][19] ),
    .B1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .X(_04942_));
 sky130_fd_sc_hd__or3_2 _17714_ (.A(_04939_),
    .B(_04941_),
    .C(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__o21ai_2 _17715_ (.A1(_04941_),
    .A2(_04942_),
    .B1(_04939_),
    .Y(_04944_));
 sky130_fd_sc_hd__a32o_2 _17716_ (.A1(_11712_),
    .A2(_04943_),
    .A3(_04944_),
    .B1(\systolic_inst.acc_wires[10][20] ),
    .B2(_11258_),
    .X(_01318_));
 sky130_fd_sc_hd__xnor2_2 _17717_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][21] ),
    .Y(_04945_));
 sky130_fd_sc_hd__inv_2 _17718_ (.A(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__a21oi_2 _17719_ (.A1(_04938_),
    .A2(_04944_),
    .B1(_04945_),
    .Y(_04947_));
 sky130_fd_sc_hd__a31o_2 _17720_ (.A1(_04938_),
    .A2(_04944_),
    .A3(_04945_),
    .B1(_11713_),
    .X(_04948_));
 sky130_fd_sc_hd__a2bb2o_2 _17721_ (.A1_N(_04948_),
    .A2_N(_04947_),
    .B1(\systolic_inst.acc_wires[10][21] ),
    .B2(_11258_),
    .X(_01319_));
 sky130_fd_sc_hd__or2_2 _17722_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][22] ),
    .X(_04949_));
 sky130_fd_sc_hd__nand2_2 _17723_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][22] ),
    .Y(_04950_));
 sky130_fd_sc_hd__and2_2 _17724_ (.A(_04949_),
    .B(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__o21a_2 _17725_ (.A1(\systolic_inst.acc_wires[10][20] ),
    .A2(\systolic_inst.acc_wires[10][21] ),
    .B1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .X(_04952_));
 sky130_fd_sc_hd__nor2_2 _17726_ (.A(_04944_),
    .B(_04945_),
    .Y(_04953_));
 sky130_fd_sc_hd__o21ai_2 _17727_ (.A1(_04952_),
    .A2(_04953_),
    .B1(_04951_),
    .Y(_04954_));
 sky130_fd_sc_hd__or3_2 _17728_ (.A(_04951_),
    .B(_04952_),
    .C(_04953_),
    .X(_04955_));
 sky130_fd_sc_hd__a32o_2 _17729_ (.A1(_11712_),
    .A2(_04954_),
    .A3(_04955_),
    .B1(\systolic_inst.acc_wires[10][22] ),
    .B2(_11258_),
    .X(_01320_));
 sky130_fd_sc_hd__xor2_2 _17730_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][23] ),
    .X(_04956_));
 sky130_fd_sc_hd__inv_2 _17731_ (.A(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__nand3_2 _17732_ (.A(_04950_),
    .B(_04954_),
    .C(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__a21o_2 _17733_ (.A1(_04950_),
    .A2(_04954_),
    .B1(_04957_),
    .X(_04959_));
 sky130_fd_sc_hd__a32o_2 _17734_ (.A1(_11712_),
    .A2(_04958_),
    .A3(_04959_),
    .B1(\systolic_inst.acc_wires[10][23] ),
    .B2(_11258_),
    .X(_01321_));
 sky130_fd_sc_hd__nand4_2 _17735_ (.A(_04939_),
    .B(_04946_),
    .C(_04951_),
    .D(_04956_),
    .Y(_04960_));
 sky130_fd_sc_hd__a211o_2 _17736_ (.A1(_04917_),
    .A2(_04918_),
    .B1(_04940_),
    .C1(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__o41a_2 _17737_ (.A1(\systolic_inst.acc_wires[10][20] ),
    .A2(\systolic_inst.acc_wires[10][21] ),
    .A3(\systolic_inst.acc_wires[10][22] ),
    .A4(\systolic_inst.acc_wires[10][23] ),
    .B1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .X(_04962_));
 sky130_fd_sc_hd__nor2_2 _17738_ (.A(_04942_),
    .B(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__nor2_2 _17739_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][24] ),
    .Y(_04964_));
 sky130_fd_sc_hd__and2_2 _17740_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][24] ),
    .X(_04965_));
 sky130_fd_sc_hd__or2_2 _17741_ (.A(_04964_),
    .B(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__a21oi_2 _17742_ (.A1(_04961_),
    .A2(_04963_),
    .B1(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__a31o_2 _17743_ (.A1(_04961_),
    .A2(_04963_),
    .A3(_04966_),
    .B1(_11713_),
    .X(_04968_));
 sky130_fd_sc_hd__a2bb2o_2 _17744_ (.A1_N(_04968_),
    .A2_N(_04967_),
    .B1(\systolic_inst.acc_wires[10][24] ),
    .B2(_11258_),
    .X(_01322_));
 sky130_fd_sc_hd__xor2_2 _17745_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][25] ),
    .X(_04969_));
 sky130_fd_sc_hd__or3_2 _17746_ (.A(_04965_),
    .B(_04967_),
    .C(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__o21ai_2 _17747_ (.A1(_04965_),
    .A2(_04967_),
    .B1(_04969_),
    .Y(_04971_));
 sky130_fd_sc_hd__a32o_2 _17748_ (.A1(_11712_),
    .A2(_04970_),
    .A3(_04971_),
    .B1(\systolic_inst.acc_wires[10][25] ),
    .B2(_11258_),
    .X(_01323_));
 sky130_fd_sc_hd__or2_2 _17749_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][26] ),
    .X(_04972_));
 sky130_fd_sc_hd__nand2_2 _17750_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][26] ),
    .Y(_04973_));
 sky130_fd_sc_hd__nand2_2 _17751_ (.A(_04972_),
    .B(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__o21a_2 _17752_ (.A1(\systolic_inst.acc_wires[10][24] ),
    .A2(\systolic_inst.acc_wires[10][25] ),
    .B1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .X(_04975_));
 sky130_fd_sc_hd__a21o_2 _17753_ (.A1(_04967_),
    .A2(_04969_),
    .B1(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__xnor2_2 _17754_ (.A(_04974_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__a22o_2 _17755_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][26] ),
    .B1(_11712_),
    .B2(_04977_),
    .X(_01324_));
 sky130_fd_sc_hd__xnor2_2 _17756_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][27] ),
    .Y(_04978_));
 sky130_fd_sc_hd__a21bo_2 _17757_ (.A1(_04972_),
    .A2(_04976_),
    .B1_N(_04973_),
    .X(_04979_));
 sky130_fd_sc_hd__xnor2_2 _17758_ (.A(_04978_),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__a22o_2 _17759_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][27] ),
    .B1(_11712_),
    .B2(_04980_),
    .X(_01325_));
 sky130_fd_sc_hd__nor2_2 _17760_ (.A(_04974_),
    .B(_04978_),
    .Y(_04981_));
 sky130_fd_sc_hd__o21a_2 _17761_ (.A1(\systolic_inst.acc_wires[10][26] ),
    .A2(\systolic_inst.acc_wires[10][27] ),
    .B1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .X(_04982_));
 sky130_fd_sc_hd__a311oi_2 _17762_ (.A1(_04967_),
    .A2(_04969_),
    .A3(_04981_),
    .B1(_04982_),
    .C1(_04975_),
    .Y(_04983_));
 sky130_fd_sc_hd__or2_2 _17763_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][28] ),
    .X(_04984_));
 sky130_fd_sc_hd__nand2_2 _17764_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][28] ),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_2 _17765_ (.A(_04984_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__xor2_2 _17766_ (.A(_04983_),
    .B(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__a22o_2 _17767_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][28] ),
    .B1(_11712_),
    .B2(_04987_),
    .X(_01326_));
 sky130_fd_sc_hd__xor2_2 _17768_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][29] ),
    .X(_04988_));
 sky130_fd_sc_hd__inv_2 _17769_ (.A(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__o21a_2 _17770_ (.A1(_04983_),
    .A2(_04986_),
    .B1(_04985_),
    .X(_04990_));
 sky130_fd_sc_hd__xnor2_2 _17771_ (.A(_04988_),
    .B(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__a22o_2 _17772_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[10][29] ),
    .B1(_11712_),
    .B2(_04991_),
    .X(_01327_));
 sky130_fd_sc_hd__o21ai_2 _17773_ (.A1(\systolic_inst.acc_wires[10][28] ),
    .A2(\systolic_inst.acc_wires[10][29] ),
    .B1(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .Y(_04992_));
 sky130_fd_sc_hd__o31a_2 _17774_ (.A1(_04983_),
    .A2(_04986_),
    .A3(_04989_),
    .B1(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__nand2_2 _17775_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][30] ),
    .Y(_04994_));
 sky130_fd_sc_hd__or2_2 _17776_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][30] ),
    .X(_04995_));
 sky130_fd_sc_hd__nand2_2 _17777_ (.A(_04994_),
    .B(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_2 _17778_ (.A(_04993_),
    .B(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__or2_2 _17779_ (.A(_04993_),
    .B(_04996_),
    .X(_04998_));
 sky130_fd_sc_hd__a32o_2 _17780_ (.A1(_11712_),
    .A2(_04997_),
    .A3(_04998_),
    .B1(\systolic_inst.acc_wires[10][30] ),
    .B2(_11258_),
    .X(_01328_));
 sky130_fd_sc_hd__xnor2_2 _17781_ (.A(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[10][31] ),
    .Y(_04999_));
 sky130_fd_sc_hd__a21oi_2 _17782_ (.A1(_04994_),
    .A2(_04998_),
    .B1(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__a31o_2 _17783_ (.A1(_04994_),
    .A2(_04998_),
    .A3(_04999_),
    .B1(_11713_),
    .X(_05001_));
 sky130_fd_sc_hd__a2bb2o_2 _17784_ (.A1_N(_05001_),
    .A2_N(_05000_),
    .B1(\systolic_inst.acc_wires[10][31] ),
    .B2(_11258_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _17785_ (.A0(\systolic_inst.A_outs[9][0] ),
    .A1(\systolic_inst.A_outs[8][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _17786_ (.A0(\systolic_inst.A_outs[9][1] ),
    .A1(\systolic_inst.A_outs[8][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _17787_ (.A0(\systolic_inst.A_outs[9][2] ),
    .A1(\systolic_inst.A_outs[8][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _17788_ (.A0(\systolic_inst.A_outs[9][3] ),
    .A1(\systolic_inst.A_outs[8][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _17789_ (.A0(\systolic_inst.A_outs[9][4] ),
    .A1(\systolic_inst.A_outs[8][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _17790_ (.A0(\systolic_inst.A_outs[9][5] ),
    .A1(\systolic_inst.A_outs[8][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _17791_ (.A0(\systolic_inst.A_outs[9][6] ),
    .A1(\systolic_inst.A_outs[8][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _17792_ (.A0(\systolic_inst.A_outs[9][7] ),
    .A1(\systolic_inst.A_outs[8][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _17793_ (.A0(\systolic_inst.B_outs[8][0] ),
    .A1(\systolic_inst.B_outs[4][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _17794_ (.A0(\systolic_inst.B_outs[8][1] ),
    .A1(\systolic_inst.B_outs[4][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _17795_ (.A0(\systolic_inst.B_outs[8][2] ),
    .A1(\systolic_inst.B_outs[4][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _17796_ (.A0(\systolic_inst.B_outs[8][3] ),
    .A1(\systolic_inst.B_outs[4][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _17797_ (.A0(\systolic_inst.B_outs[8][4] ),
    .A1(\systolic_inst.B_outs[4][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _17798_ (.A0(\systolic_inst.B_outs[8][5] ),
    .A1(\systolic_inst.B_outs[4][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _17799_ (.A0(\systolic_inst.B_outs[8][6] ),
    .A1(\systolic_inst.B_outs[4][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _17800_ (.A0(\systolic_inst.B_outs[8][7] ),
    .A1(\systolic_inst.B_outs[4][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01345_));
 sky130_fd_sc_hd__and3_2 _17801_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[9][0] ),
    .C(\systolic_inst.A_outs[9][0] ),
    .X(_05002_));
 sky130_fd_sc_hd__a21o_2 _17802_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[0] ),
    .B1(_05002_),
    .X(_01346_));
 sky130_fd_sc_hd__and4_2 _17803_ (.A(\systolic_inst.B_outs[9][0] ),
    .B(\systolic_inst.A_outs[9][0] ),
    .C(\systolic_inst.B_outs[9][1] ),
    .D(\systolic_inst.A_outs[9][1] ),
    .X(_05003_));
 sky130_fd_sc_hd__inv_2 _17804_ (.A(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__a22o_2 _17805_ (.A1(\systolic_inst.A_outs[9][0] ),
    .A2(\systolic_inst.B_outs[9][1] ),
    .B1(\systolic_inst.A_outs[9][1] ),
    .B2(\systolic_inst.B_outs[9][0] ),
    .X(_05005_));
 sky130_fd_sc_hd__and2_2 _17806_ (.A(\systolic_inst.ce_local ),
    .B(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__a22o_2 _17807_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[1] ),
    .B1(_05004_),
    .B2(_05006_),
    .X(_01347_));
 sky130_fd_sc_hd__nand2_2 _17808_ (.A(\systolic_inst.B_outs[9][1] ),
    .B(\systolic_inst.A_outs[9][1] ),
    .Y(_05007_));
 sky130_fd_sc_hd__nand2_2 _17809_ (.A(\systolic_inst.B_outs[9][0] ),
    .B(\systolic_inst.A_outs[9][2] ),
    .Y(_05008_));
 sky130_fd_sc_hd__and4_2 _17810_ (.A(\systolic_inst.B_outs[9][0] ),
    .B(\systolic_inst.B_outs[9][1] ),
    .C(\systolic_inst.A_outs[9][1] ),
    .D(\systolic_inst.A_outs[9][2] ),
    .X(_05009_));
 sky130_fd_sc_hd__a21o_2 _17811_ (.A1(_05007_),
    .A2(_05008_),
    .B1(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__xnor2_2 _17812_ (.A(_05003_),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__and2_2 _17813_ (.A(\systolic_inst.A_outs[9][0] ),
    .B(\systolic_inst.B_outs[9][2] ),
    .X(_05012_));
 sky130_fd_sc_hd__nand2_2 _17814_ (.A(_05011_),
    .B(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__o21a_2 _17815_ (.A1(_05011_),
    .A2(_05012_),
    .B1(\systolic_inst.ce_local ),
    .X(_05014_));
 sky130_fd_sc_hd__a22o_2 _17816_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[2] ),
    .B1(_05013_),
    .B2(_05014_),
    .X(_01348_));
 sky130_fd_sc_hd__a22oi_2 _17817_ (.A1(\systolic_inst.A_outs[9][1] ),
    .A2(\systolic_inst.B_outs[9][2] ),
    .B1(\systolic_inst.B_outs[9][3] ),
    .B2(\systolic_inst.A_outs[9][0] ),
    .Y(_05015_));
 sky130_fd_sc_hd__and4_2 _17818_ (.A(\systolic_inst.A_outs[9][0] ),
    .B(\systolic_inst.A_outs[9][1] ),
    .C(\systolic_inst.B_outs[9][2] ),
    .D(\systolic_inst.B_outs[9][3] ),
    .X(_05016_));
 sky130_fd_sc_hd__or2_2 _17819_ (.A(_05015_),
    .B(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__nand2_2 _17820_ (.A(\systolic_inst.B_outs[9][1] ),
    .B(\systolic_inst.A_outs[9][3] ),
    .Y(_05018_));
 sky130_fd_sc_hd__or2_2 _17821_ (.A(_05008_),
    .B(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__a22o_2 _17822_ (.A1(\systolic_inst.B_outs[9][1] ),
    .A2(\systolic_inst.A_outs[9][2] ),
    .B1(\systolic_inst.A_outs[9][3] ),
    .B2(\systolic_inst.B_outs[9][0] ),
    .X(_05020_));
 sky130_fd_sc_hd__nand3_2 _17823_ (.A(_05009_),
    .B(_05019_),
    .C(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__a21o_2 _17824_ (.A1(_05019_),
    .A2(_05020_),
    .B1(_05009_),
    .X(_05022_));
 sky130_fd_sc_hd__nand2_2 _17825_ (.A(_05021_),
    .B(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__or2_2 _17826_ (.A(_05017_),
    .B(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__xnor2_2 _17827_ (.A(_05017_),
    .B(_05023_),
    .Y(_05025_));
 sky130_fd_sc_hd__o21ai_2 _17828_ (.A1(_05004_),
    .A2(_05010_),
    .B1(_05013_),
    .Y(_05026_));
 sky130_fd_sc_hd__and2b_2 _17829_ (.A_N(_05025_),
    .B(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__xnor2_2 _17830_ (.A(_05025_),
    .B(_05026_),
    .Y(_05028_));
 sky130_fd_sc_hd__mux2_1 _17831_ (.A0(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[3] ),
    .A1(_05028_),
    .S(\systolic_inst.ce_local ),
    .X(_01349_));
 sky130_fd_sc_hd__and2_2 _17832_ (.A(\systolic_inst.B_outs[9][2] ),
    .B(\systolic_inst.A_outs[9][2] ),
    .X(_05029_));
 sky130_fd_sc_hd__nand4_2 _17833_ (.A(\systolic_inst.A_outs[9][0] ),
    .B(\systolic_inst.A_outs[9][1] ),
    .C(\systolic_inst.B_outs[9][3] ),
    .D(\systolic_inst.B_outs[9][4] ),
    .Y(_05030_));
 sky130_fd_sc_hd__a22o_2 _17834_ (.A1(\systolic_inst.A_outs[9][1] ),
    .A2(\systolic_inst.B_outs[9][3] ),
    .B1(\systolic_inst.B_outs[9][4] ),
    .B2(\systolic_inst.A_outs[9][0] ),
    .X(_05031_));
 sky130_fd_sc_hd__nand2_2 _17835_ (.A(_05030_),
    .B(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__xnor2_2 _17836_ (.A(_05029_),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__inv_2 _17837_ (.A(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand2_2 _17838_ (.A(\systolic_inst.B_outs[9][0] ),
    .B(\systolic_inst.A_outs[9][4] ),
    .Y(_05035_));
 sky130_fd_sc_hd__and4_2 _17839_ (.A(\systolic_inst.B_outs[9][0] ),
    .B(\systolic_inst.B_outs[9][1] ),
    .C(\systolic_inst.A_outs[9][3] ),
    .D(\systolic_inst.A_outs[9][4] ),
    .X(_05036_));
 sky130_fd_sc_hd__a21oi_2 _17840_ (.A1(_05018_),
    .A2(_05035_),
    .B1(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__xnor2_2 _17841_ (.A(_05016_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__nor2_2 _17842_ (.A(_05019_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__xnor2_2 _17843_ (.A(_05019_),
    .B(_05038_),
    .Y(_05040_));
 sky130_fd_sc_hd__nor2_2 _17844_ (.A(_05034_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__and2_2 _17845_ (.A(_05034_),
    .B(_05040_),
    .X(_05042_));
 sky130_fd_sc_hd__or2_2 _17846_ (.A(_05041_),
    .B(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__a21o_2 _17847_ (.A1(_05021_),
    .A2(_05024_),
    .B1(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__inv_2 _17848_ (.A(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand3_2 _17849_ (.A(_05021_),
    .B(_05024_),
    .C(_05043_),
    .Y(_05046_));
 sky130_fd_sc_hd__a21oi_2 _17850_ (.A1(_05044_),
    .A2(_05046_),
    .B1(_05027_),
    .Y(_05047_));
 sky130_fd_sc_hd__and3_2 _17851_ (.A(_05027_),
    .B(_05044_),
    .C(_05046_),
    .X(_05048_));
 sky130_fd_sc_hd__or3_2 _17852_ (.A(_11258_),
    .B(_05047_),
    .C(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__a21bo_2 _17853_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[4] ),
    .B1_N(_05049_),
    .X(_01350_));
 sky130_fd_sc_hd__a21oi_2 _17854_ (.A1(_05016_),
    .A2(_05037_),
    .B1(_05039_),
    .Y(_05050_));
 sky130_fd_sc_hd__a21bo_2 _17855_ (.A1(_05029_),
    .A2(_05031_),
    .B1_N(_05030_),
    .X(_05051_));
 sky130_fd_sc_hd__a22oi_2 _17856_ (.A1(\systolic_inst.B_outs[9][1] ),
    .A2(\systolic_inst.A_outs[9][4] ),
    .B1(\systolic_inst.A_outs[9][5] ),
    .B2(\systolic_inst.B_outs[9][0] ),
    .Y(_05052_));
 sky130_fd_sc_hd__and4_2 _17857_ (.A(\systolic_inst.B_outs[9][0] ),
    .B(\systolic_inst.B_outs[9][1] ),
    .C(\systolic_inst.A_outs[9][4] ),
    .D(\systolic_inst.A_outs[9][5] ),
    .X(_05053_));
 sky130_fd_sc_hd__or2_2 _17858_ (.A(_05052_),
    .B(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__nand2b_2 _17859_ (.A_N(_05054_),
    .B(_05051_),
    .Y(_05055_));
 sky130_fd_sc_hd__xnor2_2 _17860_ (.A(_05051_),
    .B(_05054_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_2 _17861_ (.A(_05036_),
    .B(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__xnor2_2 _17862_ (.A(_05036_),
    .B(_05056_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand2_2 _17863_ (.A(\systolic_inst.A_outs[9][0] ),
    .B(\systolic_inst.B_outs[9][5] ),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_2 _17864_ (.A(\systolic_inst.B_outs[9][2] ),
    .B(\systolic_inst.A_outs[9][3] ),
    .Y(_05060_));
 sky130_fd_sc_hd__and4_2 _17865_ (.A(\systolic_inst.A_outs[9][1] ),
    .B(\systolic_inst.A_outs[9][2] ),
    .C(\systolic_inst.B_outs[9][3] ),
    .D(\systolic_inst.B_outs[9][4] ),
    .X(_05061_));
 sky130_fd_sc_hd__a22o_2 _17866_ (.A1(\systolic_inst.A_outs[9][2] ),
    .A2(\systolic_inst.B_outs[9][3] ),
    .B1(\systolic_inst.B_outs[9][4] ),
    .B2(\systolic_inst.A_outs[9][1] ),
    .X(_05062_));
 sky130_fd_sc_hd__and2b_2 _17867_ (.A_N(_05061_),
    .B(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__xnor2_2 _17868_ (.A(_05060_),
    .B(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__nand2b_2 _17869_ (.A_N(_05059_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__xor2_2 _17870_ (.A(_05059_),
    .B(_05064_),
    .X(_05066_));
 sky130_fd_sc_hd__nor2_2 _17871_ (.A(_05058_),
    .B(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__inv_2 _17872_ (.A(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__and2_2 _17873_ (.A(_05058_),
    .B(_05066_),
    .X(_05069_));
 sky130_fd_sc_hd__nor2_2 _17874_ (.A(_05067_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__nand2_2 _17875_ (.A(_05041_),
    .B(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__or2_2 _17876_ (.A(_05041_),
    .B(_05070_),
    .X(_05072_));
 sky130_fd_sc_hd__and2_2 _17877_ (.A(_05071_),
    .B(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__nand2b_2 _17878_ (.A_N(_05050_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__xnor2_2 _17879_ (.A(_05050_),
    .B(_05073_),
    .Y(_05075_));
 sky130_fd_sc_hd__nor2_2 _17880_ (.A(_05045_),
    .B(_05048_),
    .Y(_05076_));
 sky130_fd_sc_hd__nand2b_2 _17881_ (.A_N(_05076_),
    .B(_05075_),
    .Y(_05077_));
 sky130_fd_sc_hd__o31a_2 _17882_ (.A1(_05045_),
    .A2(_05048_),
    .A3(_05075_),
    .B1(\systolic_inst.ce_local ),
    .X(_05078_));
 sky130_fd_sc_hd__a22o_2 _17883_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[5] ),
    .B1(_05077_),
    .B2(_05078_),
    .X(_01351_));
 sky130_fd_sc_hd__a31o_2 _17884_ (.A1(\systolic_inst.B_outs[9][2] ),
    .A2(\systolic_inst.A_outs[9][3] ),
    .A3(_05062_),
    .B1(_05061_),
    .X(_05079_));
 sky130_fd_sc_hd__a22oi_2 _17885_ (.A1(\systolic_inst.B_outs[9][1] ),
    .A2(\systolic_inst.A_outs[9][5] ),
    .B1(\systolic_inst.A_outs[9][6] ),
    .B2(\systolic_inst.B_outs[9][0] ),
    .Y(_05080_));
 sky130_fd_sc_hd__and4_2 _17886_ (.A(\systolic_inst.B_outs[9][0] ),
    .B(\systolic_inst.B_outs[9][1] ),
    .C(\systolic_inst.A_outs[9][5] ),
    .D(\systolic_inst.A_outs[9][6] ),
    .X(_05081_));
 sky130_fd_sc_hd__nor2_2 _17887_ (.A(_05080_),
    .B(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__xor2_2 _17888_ (.A(_05079_),
    .B(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__and2_2 _17889_ (.A(_05053_),
    .B(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__nor2_2 _17890_ (.A(_05053_),
    .B(_05083_),
    .Y(_05085_));
 sky130_fd_sc_hd__or2_2 _17891_ (.A(_05084_),
    .B(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__nand2_2 _17892_ (.A(\systolic_inst.B_outs[9][2] ),
    .B(\systolic_inst.A_outs[9][4] ),
    .Y(_05087_));
 sky130_fd_sc_hd__and4_2 _17893_ (.A(\systolic_inst.A_outs[9][2] ),
    .B(\systolic_inst.B_outs[9][3] ),
    .C(\systolic_inst.A_outs[9][3] ),
    .D(\systolic_inst.B_outs[9][4] ),
    .X(_05088_));
 sky130_fd_sc_hd__a22oi_2 _17894_ (.A1(\systolic_inst.B_outs[9][3] ),
    .A2(\systolic_inst.A_outs[9][3] ),
    .B1(\systolic_inst.B_outs[9][4] ),
    .B2(\systolic_inst.A_outs[9][2] ),
    .Y(_05089_));
 sky130_fd_sc_hd__or2_2 _17895_ (.A(_05088_),
    .B(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__xnor2_2 _17896_ (.A(_05087_),
    .B(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__a22oi_2 _17897_ (.A1(\systolic_inst.A_outs[9][1] ),
    .A2(\systolic_inst.B_outs[9][5] ),
    .B1(\systolic_inst.B_outs[9][6] ),
    .B2(\systolic_inst.A_outs[9][0] ),
    .Y(_05092_));
 sky130_fd_sc_hd__nand2_2 _17898_ (.A(\systolic_inst.A_outs[9][1] ),
    .B(\systolic_inst.B_outs[9][6] ),
    .Y(_05093_));
 sky130_fd_sc_hd__nor2_2 _17899_ (.A(_05059_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__nor2_2 _17900_ (.A(_05092_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__or3_2 _17901_ (.A(_05091_),
    .B(_05092_),
    .C(_05094_),
    .X(_05096_));
 sky130_fd_sc_hd__xor2_2 _17902_ (.A(_05091_),
    .B(_05095_),
    .X(_05097_));
 sky130_fd_sc_hd__xnor2_2 _17903_ (.A(_05065_),
    .B(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__xnor2_2 _17904_ (.A(_05086_),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__xnor2_2 _17905_ (.A(_05068_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__a21oi_2 _17906_ (.A1(_05055_),
    .A2(_05057_),
    .B1(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__and3_2 _17907_ (.A(_05055_),
    .B(_05057_),
    .C(_05100_),
    .X(_05102_));
 sky130_fd_sc_hd__a211oi_2 _17908_ (.A1(_05071_),
    .A2(_05074_),
    .B1(_05101_),
    .C1(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__o211a_2 _17909_ (.A1(_05101_),
    .A2(_05102_),
    .B1(_05071_),
    .C1(_05074_),
    .X(_05104_));
 sky130_fd_sc_hd__o21ai_2 _17910_ (.A1(_05103_),
    .A2(_05104_),
    .B1(_05077_),
    .Y(_05105_));
 sky130_fd_sc_hd__nor3_2 _17911_ (.A(_05077_),
    .B(_05103_),
    .C(_05104_),
    .Y(_05106_));
 sky130_fd_sc_hd__nor2_2 _17912_ (.A(_11258_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__a22o_2 _17913_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[6] ),
    .B1(_05105_),
    .B2(_05107_),
    .X(_01352_));
 sky130_fd_sc_hd__o21ba_2 _17914_ (.A1(_05068_),
    .A2(_05099_),
    .B1_N(_05101_),
    .X(_05108_));
 sky130_fd_sc_hd__a21oi_2 _17915_ (.A1(_05079_),
    .A2(_05082_),
    .B1(_05084_),
    .Y(_05109_));
 sky130_fd_sc_hd__o21ba_2 _17916_ (.A1(_05087_),
    .A2(_05089_),
    .B1_N(_05088_),
    .X(_05110_));
 sky130_fd_sc_hd__a22o_2 _17917_ (.A1(\systolic_inst.B_outs[9][1] ),
    .A2(\systolic_inst.A_outs[9][6] ),
    .B1(\systolic_inst.A_outs[9][7] ),
    .B2(\systolic_inst.B_outs[9][0] ),
    .X(_05111_));
 sky130_fd_sc_hd__nand4_2 _17918_ (.A(\systolic_inst.B_outs[9][0] ),
    .B(\systolic_inst.B_outs[9][1] ),
    .C(\systolic_inst.A_outs[9][6] ),
    .D(\systolic_inst.A_outs[9][7] ),
    .Y(_05112_));
 sky130_fd_sc_hd__nand2_2 _17919_ (.A(_05111_),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__xnor2_2 _17920_ (.A(_11263_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__nor2_2 _17921_ (.A(_05110_),
    .B(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__and2_2 _17922_ (.A(_05110_),
    .B(_05114_),
    .X(_05116_));
 sky130_fd_sc_hd__nor2_2 _17923_ (.A(_05115_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__xnor2_2 _17924_ (.A(_05081_),
    .B(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__nand2_2 _17925_ (.A(\systolic_inst.B_outs[9][2] ),
    .B(\systolic_inst.A_outs[9][5] ),
    .Y(_05119_));
 sky130_fd_sc_hd__and4_2 _17926_ (.A(\systolic_inst.B_outs[9][3] ),
    .B(\systolic_inst.A_outs[9][3] ),
    .C(\systolic_inst.B_outs[9][4] ),
    .D(\systolic_inst.A_outs[9][4] ),
    .X(_05120_));
 sky130_fd_sc_hd__a22oi_2 _17927_ (.A1(\systolic_inst.A_outs[9][3] ),
    .A2(\systolic_inst.B_outs[9][4] ),
    .B1(\systolic_inst.A_outs[9][4] ),
    .B2(\systolic_inst.B_outs[9][3] ),
    .Y(_05121_));
 sky130_fd_sc_hd__or2_2 _17928_ (.A(_05120_),
    .B(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__xnor2_2 _17929_ (.A(_05119_),
    .B(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__nand2_2 _17930_ (.A(\systolic_inst.A_outs[9][2] ),
    .B(\systolic_inst.B_outs[9][5] ),
    .Y(_05124_));
 sky130_fd_sc_hd__and2b_2 _17931_ (.A_N(\systolic_inst.A_outs[9][0] ),
    .B(\systolic_inst.B_outs[9][7] ),
    .X(_05125_));
 sky130_fd_sc_hd__and3_2 _17932_ (.A(\systolic_inst.A_outs[9][1] ),
    .B(\systolic_inst.B_outs[9][6] ),
    .C(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__xnor2_2 _17933_ (.A(_05093_),
    .B(_05125_),
    .Y(_05127_));
 sky130_fd_sc_hd__xnor2_2 _17934_ (.A(_05124_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__xnor2_2 _17935_ (.A(_05094_),
    .B(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__nor2_2 _17936_ (.A(_05123_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__xnor2_2 _17937_ (.A(_05123_),
    .B(_05129_),
    .Y(_05131_));
 sky130_fd_sc_hd__or2_2 _17938_ (.A(_05096_),
    .B(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__and2_2 _17939_ (.A(_05096_),
    .B(_05131_),
    .X(_05133_));
 sky130_fd_sc_hd__xor2_2 _17940_ (.A(_05096_),
    .B(_05131_),
    .X(_05134_));
 sky130_fd_sc_hd__xnor2_2 _17941_ (.A(_05118_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__o32a_2 _17942_ (.A1(_05084_),
    .A2(_05085_),
    .A3(_05098_),
    .B1(_05097_),
    .B2(_05065_),
    .X(_05136_));
 sky130_fd_sc_hd__nand2b_2 _17943_ (.A_N(_05136_),
    .B(_05135_),
    .Y(_05137_));
 sky130_fd_sc_hd__xnor2_2 _17944_ (.A(_05135_),
    .B(_05136_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2b_2 _17945_ (.A_N(_05109_),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__xnor2_2 _17946_ (.A(_05109_),
    .B(_05138_),
    .Y(_05140_));
 sky130_fd_sc_hd__and2b_2 _17947_ (.A_N(_05108_),
    .B(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__xnor2_2 _17948_ (.A(_05108_),
    .B(_05140_),
    .Y(_05142_));
 sky130_fd_sc_hd__nor3_2 _17949_ (.A(_05103_),
    .B(_05106_),
    .C(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__o21a_2 _17950_ (.A1(_05103_),
    .A2(_05106_),
    .B1(_05142_),
    .X(_05144_));
 sky130_fd_sc_hd__nand2_2 _17951_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[7] ),
    .Y(_05145_));
 sky130_fd_sc_hd__o31ai_2 _17952_ (.A1(_11258_),
    .A2(_05143_),
    .A3(_05144_),
    .B1(_05145_),
    .Y(_01353_));
 sky130_fd_sc_hd__a21o_2 _17953_ (.A1(_05081_),
    .A2(_05117_),
    .B1(_05115_),
    .X(_05146_));
 sky130_fd_sc_hd__a21bo_2 _17954_ (.A1(\systolic_inst.B_outs[9][7] ),
    .A2(_05111_),
    .B1_N(_05112_),
    .X(_05147_));
 sky130_fd_sc_hd__o21bai_2 _17955_ (.A1(_05119_),
    .A2(_05121_),
    .B1_N(_05120_),
    .Y(_05148_));
 sky130_fd_sc_hd__o21a_2 _17956_ (.A1(\systolic_inst.B_outs[9][0] ),
    .A2(\systolic_inst.B_outs[9][1] ),
    .B1(\systolic_inst.A_outs[9][7] ),
    .X(_05149_));
 sky130_fd_sc_hd__o21ai_2 _17957_ (.A1(\systolic_inst.B_outs[9][0] ),
    .A2(\systolic_inst.B_outs[9][1] ),
    .B1(\systolic_inst.A_outs[9][7] ),
    .Y(_05150_));
 sky130_fd_sc_hd__a21o_2 _17958_ (.A1(\systolic_inst.B_outs[9][0] ),
    .A2(\systolic_inst.B_outs[9][1] ),
    .B1(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__and2b_2 _17959_ (.A_N(_05151_),
    .B(_05148_),
    .X(_05152_));
 sky130_fd_sc_hd__xnor2_2 _17960_ (.A(_05148_),
    .B(_05151_),
    .Y(_05153_));
 sky130_fd_sc_hd__xnor2_2 _17961_ (.A(_05147_),
    .B(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__and4_2 _17962_ (.A(\systolic_inst.B_outs[9][3] ),
    .B(\systolic_inst.B_outs[9][4] ),
    .C(\systolic_inst.A_outs[9][4] ),
    .D(\systolic_inst.A_outs[9][5] ),
    .X(_05155_));
 sky130_fd_sc_hd__a22oi_2 _17963_ (.A1(\systolic_inst.B_outs[9][4] ),
    .A2(\systolic_inst.A_outs[9][4] ),
    .B1(\systolic_inst.A_outs[9][5] ),
    .B2(\systolic_inst.B_outs[9][3] ),
    .Y(_05156_));
 sky130_fd_sc_hd__nor2_2 _17964_ (.A(_05155_),
    .B(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2_2 _17965_ (.A(\systolic_inst.B_outs[9][2] ),
    .B(\systolic_inst.A_outs[9][6] ),
    .Y(_05158_));
 sky130_fd_sc_hd__xnor2_2 _17966_ (.A(_05157_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand2_2 _17967_ (.A(\systolic_inst.A_outs[9][3] ),
    .B(\systolic_inst.B_outs[9][5] ),
    .Y(_05160_));
 sky130_fd_sc_hd__and4b_2 _17968_ (.A_N(\systolic_inst.A_outs[9][1] ),
    .B(\systolic_inst.A_outs[9][2] ),
    .C(\systolic_inst.B_outs[9][6] ),
    .D(\systolic_inst.B_outs[9][7] ),
    .X(_05161_));
 sky130_fd_sc_hd__o2bb2a_2 _17969_ (.A1_N(\systolic_inst.A_outs[9][2] ),
    .A2_N(\systolic_inst.B_outs[9][6] ),
    .B1(_11263_),
    .B2(\systolic_inst.A_outs[9][1] ),
    .X(_05162_));
 sky130_fd_sc_hd__nor2_2 _17970_ (.A(_05161_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__xnor2_2 _17971_ (.A(_05160_),
    .B(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__a31oi_2 _17972_ (.A1(\systolic_inst.A_outs[9][2] ),
    .A2(\systolic_inst.B_outs[9][5] ),
    .A3(_05127_),
    .B1(_05126_),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2b_2 _17973_ (.A_N(_05165_),
    .B(_05164_),
    .Y(_05166_));
 sky130_fd_sc_hd__xnor2_2 _17974_ (.A(_05164_),
    .B(_05165_),
    .Y(_05167_));
 sky130_fd_sc_hd__nand2_2 _17975_ (.A(_05159_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__xnor2_2 _17976_ (.A(_05159_),
    .B(_05167_),
    .Y(_05169_));
 sky130_fd_sc_hd__a21oi_2 _17977_ (.A1(_05094_),
    .A2(_05128_),
    .B1(_05130_),
    .Y(_05170_));
 sky130_fd_sc_hd__xnor2_2 _17978_ (.A(_05169_),
    .B(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__or2_2 _17979_ (.A(_05154_),
    .B(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__xor2_2 _17980_ (.A(_05154_),
    .B(_05171_),
    .X(_05173_));
 sky130_fd_sc_hd__o21a_2 _17981_ (.A1(_05118_),
    .A2(_05133_),
    .B1(_05132_),
    .X(_05174_));
 sky130_fd_sc_hd__nand2b_2 _17982_ (.A_N(_05174_),
    .B(_05173_),
    .Y(_05175_));
 sky130_fd_sc_hd__xor2_2 _17983_ (.A(_05173_),
    .B(_05174_),
    .X(_05176_));
 sky130_fd_sc_hd__nand2b_2 _17984_ (.A_N(_05176_),
    .B(_05146_),
    .Y(_05177_));
 sky130_fd_sc_hd__xor2_2 _17985_ (.A(_05146_),
    .B(_05176_),
    .X(_05178_));
 sky130_fd_sc_hd__and2_2 _17986_ (.A(_05137_),
    .B(_05139_),
    .X(_05179_));
 sky130_fd_sc_hd__or2_2 _17987_ (.A(_05178_),
    .B(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__nand2_2 _17988_ (.A(_05178_),
    .B(_05179_),
    .Y(_05181_));
 sky130_fd_sc_hd__and2_2 _17989_ (.A(_05180_),
    .B(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__o21ai_2 _17990_ (.A1(_05141_),
    .A2(_05144_),
    .B1(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__or3_2 _17991_ (.A(_05141_),
    .B(_05144_),
    .C(_05182_),
    .X(_05184_));
 sky130_fd_sc_hd__and2_2 _17992_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[8] ),
    .X(_05185_));
 sky130_fd_sc_hd__a31o_2 _17993_ (.A1(\systolic_inst.ce_local ),
    .A2(_05183_),
    .A3(_05184_),
    .B1(_05185_),
    .X(_01354_));
 sky130_fd_sc_hd__a21o_2 _17994_ (.A1(_05147_),
    .A2(_05153_),
    .B1(_05152_),
    .X(_05186_));
 sky130_fd_sc_hd__o21ba_2 _17995_ (.A1(_05156_),
    .A2(_05158_),
    .B1_N(_05155_),
    .X(_05187_));
 sky130_fd_sc_hd__nor2_2 _17996_ (.A(_05150_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__and2_2 _17997_ (.A(_05150_),
    .B(_05187_),
    .X(_05189_));
 sky130_fd_sc_hd__or2_2 _17998_ (.A(_05188_),
    .B(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__nand2_2 _17999_ (.A(\systolic_inst.B_outs[9][2] ),
    .B(\systolic_inst.A_outs[9][7] ),
    .Y(_05191_));
 sky130_fd_sc_hd__a22oi_2 _18000_ (.A1(\systolic_inst.B_outs[9][4] ),
    .A2(\systolic_inst.A_outs[9][5] ),
    .B1(\systolic_inst.A_outs[9][6] ),
    .B2(\systolic_inst.B_outs[9][3] ),
    .Y(_05192_));
 sky130_fd_sc_hd__and4_2 _18001_ (.A(\systolic_inst.B_outs[9][3] ),
    .B(\systolic_inst.B_outs[9][4] ),
    .C(\systolic_inst.A_outs[9][5] ),
    .D(\systolic_inst.A_outs[9][6] ),
    .X(_05193_));
 sky130_fd_sc_hd__nor2_2 _18002_ (.A(_05192_),
    .B(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__xnor2_2 _18003_ (.A(_05191_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__nand2_2 _18004_ (.A(\systolic_inst.A_outs[9][4] ),
    .B(\systolic_inst.B_outs[9][5] ),
    .Y(_05196_));
 sky130_fd_sc_hd__and4b_2 _18005_ (.A_N(\systolic_inst.A_outs[9][2] ),
    .B(\systolic_inst.A_outs[9][3] ),
    .C(\systolic_inst.B_outs[9][6] ),
    .D(\systolic_inst.B_outs[9][7] ),
    .X(_05197_));
 sky130_fd_sc_hd__o2bb2a_2 _18006_ (.A1_N(\systolic_inst.A_outs[9][3] ),
    .A2_N(\systolic_inst.B_outs[9][6] ),
    .B1(_11263_),
    .B2(\systolic_inst.A_outs[9][2] ),
    .X(_05198_));
 sky130_fd_sc_hd__nor2_2 _18007_ (.A(_05197_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__xnor2_2 _18008_ (.A(_05196_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__o21ba_2 _18009_ (.A1(_05160_),
    .A2(_05162_),
    .B1_N(_05161_),
    .X(_05201_));
 sky130_fd_sc_hd__nand2b_2 _18010_ (.A_N(_05201_),
    .B(_05200_),
    .Y(_05202_));
 sky130_fd_sc_hd__xnor2_2 _18011_ (.A(_05200_),
    .B(_05201_),
    .Y(_05203_));
 sky130_fd_sc_hd__xnor2_2 _18012_ (.A(_05195_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__a21o_2 _18013_ (.A1(_05166_),
    .A2(_05168_),
    .B1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__nand3_2 _18014_ (.A(_05166_),
    .B(_05168_),
    .C(_05204_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_2 _18015_ (.A(_05205_),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__xor2_2 _18016_ (.A(_05190_),
    .B(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__o21a_2 _18017_ (.A1(_05169_),
    .A2(_05170_),
    .B1(_05172_),
    .X(_05209_));
 sky130_fd_sc_hd__nand2b_2 _18018_ (.A_N(_05209_),
    .B(_05208_),
    .Y(_05210_));
 sky130_fd_sc_hd__xnor2_2 _18019_ (.A(_05208_),
    .B(_05209_),
    .Y(_05211_));
 sky130_fd_sc_hd__xnor2_2 _18020_ (.A(_05186_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__a21o_2 _18021_ (.A1(_05175_),
    .A2(_05177_),
    .B1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__and3_2 _18022_ (.A(_05175_),
    .B(_05177_),
    .C(_05212_),
    .X(_05214_));
 sky130_fd_sc_hd__inv_2 _18023_ (.A(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__nand2_2 _18024_ (.A(_05213_),
    .B(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand2_2 _18025_ (.A(_05180_),
    .B(_05183_),
    .Y(_05217_));
 sky130_fd_sc_hd__xnor2_2 _18026_ (.A(_05216_),
    .B(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__mux2_1 _18027_ (.A0(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[9] ),
    .A1(_05218_),
    .S(\systolic_inst.ce_local ),
    .X(_01355_));
 sky130_fd_sc_hd__o21ba_2 _18028_ (.A1(_05191_),
    .A2(_05192_),
    .B1_N(_05193_),
    .X(_05219_));
 sky130_fd_sc_hd__nor2_2 _18029_ (.A(_05150_),
    .B(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__and2_2 _18030_ (.A(_05150_),
    .B(_05219_),
    .X(_05221_));
 sky130_fd_sc_hd__or2_2 _18031_ (.A(_05220_),
    .B(_05221_),
    .X(_05222_));
 sky130_fd_sc_hd__a22o_2 _18032_ (.A1(\systolic_inst.B_outs[9][4] ),
    .A2(\systolic_inst.A_outs[9][6] ),
    .B1(\systolic_inst.A_outs[9][7] ),
    .B2(\systolic_inst.B_outs[9][3] ),
    .X(_05223_));
 sky130_fd_sc_hd__and3_2 _18033_ (.A(\systolic_inst.B_outs[9][3] ),
    .B(\systolic_inst.B_outs[9][4] ),
    .C(\systolic_inst.A_outs[9][7] ),
    .X(_05224_));
 sky130_fd_sc_hd__a21bo_2 _18034_ (.A1(\systolic_inst.A_outs[9][6] ),
    .A2(_05224_),
    .B1_N(_05223_),
    .X(_05225_));
 sky130_fd_sc_hd__xor2_2 _18035_ (.A(_05191_),
    .B(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__nand2_2 _18036_ (.A(\systolic_inst.B_outs[9][5] ),
    .B(\systolic_inst.A_outs[9][5] ),
    .Y(_05227_));
 sky130_fd_sc_hd__and4b_2 _18037_ (.A_N(\systolic_inst.A_outs[9][3] ),
    .B(\systolic_inst.A_outs[9][4] ),
    .C(\systolic_inst.B_outs[9][6] ),
    .D(\systolic_inst.B_outs[9][7] ),
    .X(_05228_));
 sky130_fd_sc_hd__o2bb2a_2 _18038_ (.A1_N(\systolic_inst.A_outs[9][4] ),
    .A2_N(\systolic_inst.B_outs[9][6] ),
    .B1(_11263_),
    .B2(\systolic_inst.A_outs[9][3] ),
    .X(_05229_));
 sky130_fd_sc_hd__nor2_2 _18039_ (.A(_05228_),
    .B(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__xnor2_2 _18040_ (.A(_05227_),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__o21ba_2 _18041_ (.A1(_05196_),
    .A2(_05198_),
    .B1_N(_05197_),
    .X(_05232_));
 sky130_fd_sc_hd__nand2b_2 _18042_ (.A_N(_05232_),
    .B(_05231_),
    .Y(_05233_));
 sky130_fd_sc_hd__xnor2_2 _18043_ (.A(_05231_),
    .B(_05232_),
    .Y(_05234_));
 sky130_fd_sc_hd__nand2_2 _18044_ (.A(_05226_),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__or2_2 _18045_ (.A(_05226_),
    .B(_05234_),
    .X(_05236_));
 sky130_fd_sc_hd__nand2_2 _18046_ (.A(_05235_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__a21bo_2 _18047_ (.A1(_05195_),
    .A2(_05203_),
    .B1_N(_05202_),
    .X(_05238_));
 sky130_fd_sc_hd__nand2b_2 _18048_ (.A_N(_05237_),
    .B(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__xor2_2 _18049_ (.A(_05237_),
    .B(_05238_),
    .X(_05240_));
 sky130_fd_sc_hd__xor2_2 _18050_ (.A(_05222_),
    .B(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__o21a_2 _18051_ (.A1(_05190_),
    .A2(_05207_),
    .B1(_05205_),
    .X(_05242_));
 sky130_fd_sc_hd__nand2b_2 _18052_ (.A_N(_05242_),
    .B(_05241_),
    .Y(_05243_));
 sky130_fd_sc_hd__xnor2_2 _18053_ (.A(_05241_),
    .B(_05242_),
    .Y(_05244_));
 sky130_fd_sc_hd__nand2_2 _18054_ (.A(_05188_),
    .B(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__or2_2 _18055_ (.A(_05188_),
    .B(_05244_),
    .X(_05246_));
 sky130_fd_sc_hd__nand2_2 _18056_ (.A(_05245_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__a21boi_2 _18057_ (.A1(_05186_),
    .A2(_05211_),
    .B1_N(_05210_),
    .Y(_05248_));
 sky130_fd_sc_hd__nor2_2 _18058_ (.A(_05247_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__xnor2_2 _18059_ (.A(_05247_),
    .B(_05248_),
    .Y(_05250_));
 sky130_fd_sc_hd__a31o_2 _18060_ (.A1(_05180_),
    .A2(_05183_),
    .A3(_05213_),
    .B1(_05214_),
    .X(_05251_));
 sky130_fd_sc_hd__a311oi_2 _18061_ (.A1(_05180_),
    .A2(_05183_),
    .A3(_05213_),
    .B1(_05214_),
    .C1(_05250_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand2_2 _18062_ (.A(_05250_),
    .B(_05251_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2b_2 _18063_ (.A_N(_05252_),
    .B(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__nor2_2 _18064_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[10] ),
    .Y(_05255_));
 sky130_fd_sc_hd__a21oi_2 _18065_ (.A1(\systolic_inst.ce_local ),
    .A2(_05254_),
    .B1(_05255_),
    .Y(_01356_));
 sky130_fd_sc_hd__o2bb2a_2 _18066_ (.A1_N(\systolic_inst.A_outs[9][6] ),
    .A2_N(_05224_),
    .B1(_05225_),
    .B2(_05191_),
    .X(_05256_));
 sky130_fd_sc_hd__or2_2 _18067_ (.A(_05150_),
    .B(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__nand2_2 _18068_ (.A(_05150_),
    .B(_05256_),
    .Y(_05258_));
 sky130_fd_sc_hd__nand2_2 _18069_ (.A(_05257_),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__or2_2 _18070_ (.A(\systolic_inst.B_outs[9][3] ),
    .B(\systolic_inst.B_outs[9][4] ),
    .X(_05260_));
 sky130_fd_sc_hd__and3b_2 _18071_ (.A_N(_05224_),
    .B(_05260_),
    .C(\systolic_inst.A_outs[9][7] ),
    .X(_05261_));
 sky130_fd_sc_hd__xnor2_2 _18072_ (.A(_05191_),
    .B(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__nand2_2 _18073_ (.A(\systolic_inst.B_outs[9][5] ),
    .B(\systolic_inst.A_outs[9][6] ),
    .Y(_05263_));
 sky130_fd_sc_hd__and4b_2 _18074_ (.A_N(\systolic_inst.A_outs[9][4] ),
    .B(\systolic_inst.A_outs[9][5] ),
    .C(\systolic_inst.B_outs[9][6] ),
    .D(\systolic_inst.B_outs[9][7] ),
    .X(_05264_));
 sky130_fd_sc_hd__o2bb2a_2 _18075_ (.A1_N(\systolic_inst.A_outs[9][5] ),
    .A2_N(\systolic_inst.B_outs[9][6] ),
    .B1(_11263_),
    .B2(\systolic_inst.A_outs[9][4] ),
    .X(_05265_));
 sky130_fd_sc_hd__nor2_2 _18076_ (.A(_05264_),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__xnor2_2 _18077_ (.A(_05263_),
    .B(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__o21ba_2 _18078_ (.A1(_05227_),
    .A2(_05229_),
    .B1_N(_05228_),
    .X(_05268_));
 sky130_fd_sc_hd__nand2b_2 _18079_ (.A_N(_05268_),
    .B(_05267_),
    .Y(_05269_));
 sky130_fd_sc_hd__xnor2_2 _18080_ (.A(_05267_),
    .B(_05268_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2_2 _18081_ (.A(_05262_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__xnor2_2 _18082_ (.A(_05262_),
    .B(_05270_),
    .Y(_05272_));
 sky130_fd_sc_hd__a21o_2 _18083_ (.A1(_05233_),
    .A2(_05235_),
    .B1(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__nand3_2 _18084_ (.A(_05233_),
    .B(_05235_),
    .C(_05272_),
    .Y(_05274_));
 sky130_fd_sc_hd__nand2_2 _18085_ (.A(_05273_),
    .B(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__xor2_2 _18086_ (.A(_05259_),
    .B(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__o21a_2 _18087_ (.A1(_05222_),
    .A2(_05240_),
    .B1(_05239_),
    .X(_05277_));
 sky130_fd_sc_hd__and2b_2 _18088_ (.A_N(_05277_),
    .B(_05276_),
    .X(_05278_));
 sky130_fd_sc_hd__and2b_2 _18089_ (.A_N(_05276_),
    .B(_05277_),
    .X(_05279_));
 sky130_fd_sc_hd__nor2_2 _18090_ (.A(_05278_),
    .B(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__xnor2_2 _18091_ (.A(_05220_),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__nand3_2 _18092_ (.A(_05243_),
    .B(_05245_),
    .C(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__inv_2 _18093_ (.A(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__a21oi_2 _18094_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_05281_),
    .Y(_05284_));
 sky130_fd_sc_hd__nor2_2 _18095_ (.A(_05283_),
    .B(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__nor2_2 _18096_ (.A(_05249_),
    .B(_05252_),
    .Y(_05286_));
 sky130_fd_sc_hd__xnor2_2 _18097_ (.A(_05285_),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__mux2_1 _18098_ (.A0(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[11] ),
    .A1(_05287_),
    .S(\systolic_inst.ce_local ),
    .X(_01357_));
 sky130_fd_sc_hd__a31o_2 _18099_ (.A1(\systolic_inst.B_outs[9][2] ),
    .A2(\systolic_inst.A_outs[9][7] ),
    .A3(_05260_),
    .B1(_05224_),
    .X(_05288_));
 sky130_fd_sc_hd__or2_2 _18100_ (.A(_05149_),
    .B(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__nand2_2 _18101_ (.A(_05149_),
    .B(_05288_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand2_2 _18102_ (.A(_05289_),
    .B(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__inv_2 _18103_ (.A(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__o2bb2a_2 _18104_ (.A1_N(\systolic_inst.B_outs[9][6] ),
    .A2_N(\systolic_inst.A_outs[9][6] ),
    .B1(_11263_),
    .B2(\systolic_inst.A_outs[9][5] ),
    .X(_05293_));
 sky130_fd_sc_hd__and4b_2 _18105_ (.A_N(\systolic_inst.A_outs[9][5] ),
    .B(\systolic_inst.B_outs[9][6] ),
    .C(\systolic_inst.A_outs[9][6] ),
    .D(\systolic_inst.B_outs[9][7] ),
    .X(_05294_));
 sky130_fd_sc_hd__nor2_2 _18106_ (.A(_05293_),
    .B(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__nand2_2 _18107_ (.A(\systolic_inst.B_outs[9][5] ),
    .B(\systolic_inst.A_outs[9][7] ),
    .Y(_05296_));
 sky130_fd_sc_hd__xnor2_2 _18108_ (.A(_05295_),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__o21ba_2 _18109_ (.A1(_05263_),
    .A2(_05265_),
    .B1_N(_05264_),
    .X(_05298_));
 sky130_fd_sc_hd__nand2b_2 _18110_ (.A_N(_05298_),
    .B(_05297_),
    .Y(_05299_));
 sky130_fd_sc_hd__xnor2_2 _18111_ (.A(_05297_),
    .B(_05298_),
    .Y(_05300_));
 sky130_fd_sc_hd__xnor2_2 _18112_ (.A(_05262_),
    .B(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__a21o_2 _18113_ (.A1(_05269_),
    .A2(_05271_),
    .B1(_05301_),
    .X(_05302_));
 sky130_fd_sc_hd__nand3_2 _18114_ (.A(_05269_),
    .B(_05271_),
    .C(_05301_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand2_2 _18115_ (.A(_05302_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__xnor2_2 _18116_ (.A(_05292_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__o21a_2 _18117_ (.A1(_05259_),
    .A2(_05275_),
    .B1(_05273_),
    .X(_05306_));
 sky130_fd_sc_hd__and2b_2 _18118_ (.A_N(_05306_),
    .B(_05305_),
    .X(_05307_));
 sky130_fd_sc_hd__and2b_2 _18119_ (.A_N(_05305_),
    .B(_05306_),
    .X(_05308_));
 sky130_fd_sc_hd__nor2_2 _18120_ (.A(_05307_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__and2b_2 _18121_ (.A_N(_05257_),
    .B(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__xor2_2 _18122_ (.A(_05257_),
    .B(_05309_),
    .X(_05311_));
 sky130_fd_sc_hd__a21oi_2 _18123_ (.A1(_05220_),
    .A2(_05280_),
    .B1(_05278_),
    .Y(_05312_));
 sky130_fd_sc_hd__nor2_2 _18124_ (.A(_05311_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__and2_2 _18125_ (.A(_05311_),
    .B(_05312_),
    .X(_05314_));
 sky130_fd_sc_hd__nor2_2 _18126_ (.A(_05313_),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__o31a_2 _18127_ (.A1(_05249_),
    .A2(_05252_),
    .A3(_05284_),
    .B1(_05282_),
    .X(_05316_));
 sky130_fd_sc_hd__o311a_2 _18128_ (.A1(_05249_),
    .A2(_05252_),
    .A3(_05284_),
    .B1(_05315_),
    .C1(_05282_),
    .X(_05317_));
 sky130_fd_sc_hd__nor2_2 _18129_ (.A(_05315_),
    .B(_05316_),
    .Y(_05318_));
 sky130_fd_sc_hd__nor2_2 _18130_ (.A(_05317_),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__mux2_1 _18131_ (.A0(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[12] ),
    .A1(_05319_),
    .S(\systolic_inst.ce_local ),
    .X(_01358_));
 sky130_fd_sc_hd__nand2_2 _18132_ (.A(\systolic_inst.B_outs[9][6] ),
    .B(\systolic_inst.A_outs[9][7] ),
    .Y(_05320_));
 sky130_fd_sc_hd__or2_2 _18133_ (.A(\systolic_inst.A_outs[9][6] ),
    .B(_11263_),
    .X(_05321_));
 sky130_fd_sc_hd__and2_2 _18134_ (.A(_05320_),
    .B(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__nor2_2 _18135_ (.A(_05320_),
    .B(_05321_),
    .Y(_05323_));
 sky130_fd_sc_hd__nor2_2 _18136_ (.A(_05322_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__xnor2_2 _18137_ (.A(_05296_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__o21ba_2 _18138_ (.A1(_05293_),
    .A2(_05296_),
    .B1_N(_05294_),
    .X(_05326_));
 sky130_fd_sc_hd__nand2b_2 _18139_ (.A_N(_05326_),
    .B(_05325_),
    .Y(_05327_));
 sky130_fd_sc_hd__xnor2_2 _18140_ (.A(_05325_),
    .B(_05326_),
    .Y(_05328_));
 sky130_fd_sc_hd__nand2_2 _18141_ (.A(_05262_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__or2_2 _18142_ (.A(_05262_),
    .B(_05328_),
    .X(_05330_));
 sky130_fd_sc_hd__nand2_2 _18143_ (.A(_05329_),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__a21bo_2 _18144_ (.A1(_05262_),
    .A2(_05300_),
    .B1_N(_05299_),
    .X(_05332_));
 sky130_fd_sc_hd__nand2b_2 _18145_ (.A_N(_05331_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__xor2_2 _18146_ (.A(_05331_),
    .B(_05332_),
    .X(_05334_));
 sky130_fd_sc_hd__xnor2_2 _18147_ (.A(_05292_),
    .B(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__o21a_2 _18148_ (.A1(_05291_),
    .A2(_05304_),
    .B1(_05302_),
    .X(_05336_));
 sky130_fd_sc_hd__and2b_2 _18149_ (.A_N(_05336_),
    .B(_05335_),
    .X(_05337_));
 sky130_fd_sc_hd__and2b_2 _18150_ (.A_N(_05335_),
    .B(_05336_),
    .X(_05338_));
 sky130_fd_sc_hd__nor2_2 _18151_ (.A(_05337_),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__xnor2_2 _18152_ (.A(_05290_),
    .B(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__nor3_2 _18153_ (.A(_05307_),
    .B(_05310_),
    .C(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__o21a_2 _18154_ (.A1(_05307_),
    .A2(_05310_),
    .B1(_05340_),
    .X(_05342_));
 sky130_fd_sc_hd__nor2_2 _18155_ (.A(_05341_),
    .B(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__o21ai_2 _18156_ (.A1(_05313_),
    .A2(_05317_),
    .B1(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__o31a_2 _18157_ (.A1(_05313_),
    .A2(_05317_),
    .A3(_05343_),
    .B1(\systolic_inst.ce_local ),
    .X(_05345_));
 sky130_fd_sc_hd__a22o_2 _18158_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[13] ),
    .B1(_05344_),
    .B2(_05345_),
    .X(_01359_));
 sky130_fd_sc_hd__and2_2 _18159_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[14] ),
    .X(_05346_));
 sky130_fd_sc_hd__a31o_2 _18160_ (.A1(\systolic_inst.B_outs[9][5] ),
    .A2(\systolic_inst.A_outs[9][7] ),
    .A3(_05324_),
    .B1(_05323_),
    .X(_05347_));
 sky130_fd_sc_hd__nand3_2 _18161_ (.A(\systolic_inst.B_outs[9][5] ),
    .B(\systolic_inst.B_outs[9][6] ),
    .C(\systolic_inst.A_outs[9][7] ),
    .Y(_05348_));
 sky130_fd_sc_hd__o211a_2 _18162_ (.A1(_11263_),
    .A2(\systolic_inst.A_outs[9][7] ),
    .B1(_05296_),
    .C1(_05320_),
    .X(_05349_));
 sky130_fd_sc_hd__a21oi_2 _18163_ (.A1(_05347_),
    .A2(_05348_),
    .B1(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__or2_2 _18164_ (.A(_05262_),
    .B(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__nand2_2 _18165_ (.A(_05262_),
    .B(_05350_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_2 _18166_ (.A(_05351_),
    .B(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__a21oi_2 _18167_ (.A1(_05327_),
    .A2(_05329_),
    .B1(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__and3_2 _18168_ (.A(_05327_),
    .B(_05329_),
    .C(_05353_),
    .X(_05355_));
 sky130_fd_sc_hd__nor2_2 _18169_ (.A(_05354_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__xnor2_2 _18170_ (.A(_05291_),
    .B(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__o21a_2 _18171_ (.A1(_05291_),
    .A2(_05334_),
    .B1(_05333_),
    .X(_05358_));
 sky130_fd_sc_hd__and2b_2 _18172_ (.A_N(_05358_),
    .B(_05357_),
    .X(_05359_));
 sky130_fd_sc_hd__and2b_2 _18173_ (.A_N(_05357_),
    .B(_05358_),
    .X(_05360_));
 sky130_fd_sc_hd__nor2_2 _18174_ (.A(_05359_),
    .B(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__xnor2_2 _18175_ (.A(_05290_),
    .B(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__o21ba_2 _18176_ (.A1(_05290_),
    .A2(_05338_),
    .B1_N(_05337_),
    .X(_05363_));
 sky130_fd_sc_hd__nand2b_2 _18177_ (.A_N(_05363_),
    .B(_05362_),
    .Y(_05364_));
 sky130_fd_sc_hd__xnor2_2 _18178_ (.A(_05362_),
    .B(_05363_),
    .Y(_05365_));
 sky130_fd_sc_hd__and2_2 _18179_ (.A(_05317_),
    .B(_05343_),
    .X(_05366_));
 sky130_fd_sc_hd__and2b_2 _18180_ (.A_N(_05341_),
    .B(_05313_),
    .X(_05367_));
 sky130_fd_sc_hd__or4_2 _18181_ (.A(_05342_),
    .B(_05365_),
    .C(_05366_),
    .D(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__o31ai_2 _18182_ (.A1(_05342_),
    .A2(_05366_),
    .A3(_05367_),
    .B1(_05365_),
    .Y(_05369_));
 sky130_fd_sc_hd__a31o_2 _18183_ (.A1(\systolic_inst.ce_local ),
    .A2(_05368_),
    .A3(_05369_),
    .B1(_05346_),
    .X(_01360_));
 sky130_fd_sc_hd__a31o_2 _18184_ (.A1(_05149_),
    .A2(_05288_),
    .A3(_05361_),
    .B1(_05359_),
    .X(_05370_));
 sky130_fd_sc_hd__a21oi_2 _18185_ (.A1(_05292_),
    .A2(_05356_),
    .B1(_05354_),
    .Y(_05371_));
 sky130_fd_sc_hd__xnor2_2 _18186_ (.A(_05289_),
    .B(_05351_),
    .Y(_05372_));
 sky130_fd_sc_hd__xnor2_2 _18187_ (.A(_05371_),
    .B(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__xnor2_2 _18188_ (.A(_05370_),
    .B(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__and3_2 _18189_ (.A(\systolic_inst.ce_local ),
    .B(_05364_),
    .C(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__a22o_2 _18190_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B1(_05369_),
    .B2(_05375_),
    .X(_01361_));
 sky130_fd_sc_hd__a21o_2 _18191_ (.A1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[9][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_05376_));
 sky130_fd_sc_hd__a21oi_2 _18192_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[9][0] ),
    .Y(_05377_));
 sky130_fd_sc_hd__a21oi_2 _18193_ (.A1(\systolic_inst.ce_local ),
    .A2(_05376_),
    .B1(_05377_),
    .Y(_01362_));
 sky130_fd_sc_hd__and2_2 _18194_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[9][1] ),
    .X(_05378_));
 sky130_fd_sc_hd__nand2_2 _18195_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[9][1] ),
    .Y(_05379_));
 sky130_fd_sc_hd__or2_2 _18196_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[9][1] ),
    .X(_05380_));
 sky130_fd_sc_hd__and4_2 _18197_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[9][0] ),
    .C(_05379_),
    .D(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__inv_2 _18198_ (.A(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__a22o_2 _18199_ (.A1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[9][0] ),
    .B1(_05379_),
    .B2(_05380_),
    .X(_05383_));
 sky130_fd_sc_hd__a32o_2 _18200_ (.A1(_11712_),
    .A2(_05382_),
    .A3(_05383_),
    .B1(\systolic_inst.acc_wires[9][1] ),
    .B2(_11258_),
    .X(_01363_));
 sky130_fd_sc_hd__and2_2 _18201_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[9][2] ),
    .X(_05384_));
 sky130_fd_sc_hd__nand2_2 _18202_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[9][2] ),
    .Y(_05385_));
 sky130_fd_sc_hd__or2_2 _18203_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[9][2] ),
    .X(_05386_));
 sky130_fd_sc_hd__a211o_2 _18204_ (.A1(_05385_),
    .A2(_05386_),
    .B1(_05378_),
    .C1(_05381_),
    .X(_05387_));
 sky130_fd_sc_hd__o211a_2 _18205_ (.A1(_05378_),
    .A2(_05381_),
    .B1(_05385_),
    .C1(_05386_),
    .X(_05388_));
 sky130_fd_sc_hd__inv_2 _18206_ (.A(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__a32o_2 _18207_ (.A1(_11712_),
    .A2(_05387_),
    .A3(_05389_),
    .B1(\systolic_inst.acc_wires[9][2] ),
    .B2(_11258_),
    .X(_01364_));
 sky130_fd_sc_hd__and2_2 _18208_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[9][3] ),
    .X(_05390_));
 sky130_fd_sc_hd__nand2_2 _18209_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[9][3] ),
    .Y(_05391_));
 sky130_fd_sc_hd__or2_2 _18210_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[9][3] ),
    .X(_05392_));
 sky130_fd_sc_hd__a211o_2 _18211_ (.A1(_05391_),
    .A2(_05392_),
    .B1(_05384_),
    .C1(_05388_),
    .X(_05393_));
 sky130_fd_sc_hd__o211a_2 _18212_ (.A1(_05384_),
    .A2(_05388_),
    .B1(_05391_),
    .C1(_05392_),
    .X(_05394_));
 sky130_fd_sc_hd__inv_2 _18213_ (.A(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__a32o_2 _18214_ (.A1(_11712_),
    .A2(_05393_),
    .A3(_05395_),
    .B1(\systolic_inst.acc_wires[9][3] ),
    .B2(_11258_),
    .X(_01365_));
 sky130_fd_sc_hd__and2_2 _18215_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[9][4] ),
    .X(_05396_));
 sky130_fd_sc_hd__nand2_2 _18216_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[9][4] ),
    .Y(_05397_));
 sky130_fd_sc_hd__or2_2 _18217_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[9][4] ),
    .X(_05398_));
 sky130_fd_sc_hd__a211o_2 _18218_ (.A1(_05397_),
    .A2(_05398_),
    .B1(_05390_),
    .C1(_05394_),
    .X(_05399_));
 sky130_fd_sc_hd__o211a_2 _18219_ (.A1(_05390_),
    .A2(_05394_),
    .B1(_05397_),
    .C1(_05398_),
    .X(_05400_));
 sky130_fd_sc_hd__inv_2 _18220_ (.A(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__a32o_2 _18221_ (.A1(_11712_),
    .A2(_05399_),
    .A3(_05401_),
    .B1(\systolic_inst.acc_wires[9][4] ),
    .B2(_11258_),
    .X(_01366_));
 sky130_fd_sc_hd__and2_2 _18222_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[9][5] ),
    .X(_05402_));
 sky130_fd_sc_hd__nand2_2 _18223_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[9][5] ),
    .Y(_05403_));
 sky130_fd_sc_hd__or2_2 _18224_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[9][5] ),
    .X(_05404_));
 sky130_fd_sc_hd__a211o_2 _18225_ (.A1(_05403_),
    .A2(_05404_),
    .B1(_05396_),
    .C1(_05400_),
    .X(_05405_));
 sky130_fd_sc_hd__o211a_2 _18226_ (.A1(_05396_),
    .A2(_05400_),
    .B1(_05403_),
    .C1(_05404_),
    .X(_05406_));
 sky130_fd_sc_hd__inv_2 _18227_ (.A(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__a32o_2 _18228_ (.A1(_11712_),
    .A2(_05405_),
    .A3(_05407_),
    .B1(\systolic_inst.acc_wires[9][5] ),
    .B2(_11258_),
    .X(_01367_));
 sky130_fd_sc_hd__and2_2 _18229_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[9][6] ),
    .X(_05408_));
 sky130_fd_sc_hd__nand2_2 _18230_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[9][6] ),
    .Y(_05409_));
 sky130_fd_sc_hd__or2_2 _18231_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[9][6] ),
    .X(_05410_));
 sky130_fd_sc_hd__a211o_2 _18232_ (.A1(_05409_),
    .A2(_05410_),
    .B1(_05402_),
    .C1(_05406_),
    .X(_05411_));
 sky130_fd_sc_hd__o211a_2 _18233_ (.A1(_05402_),
    .A2(_05406_),
    .B1(_05409_),
    .C1(_05410_),
    .X(_05412_));
 sky130_fd_sc_hd__inv_2 _18234_ (.A(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__a32o_2 _18235_ (.A1(_11712_),
    .A2(_05411_),
    .A3(_05413_),
    .B1(\systolic_inst.acc_wires[9][6] ),
    .B2(_11258_),
    .X(_01368_));
 sky130_fd_sc_hd__nand2_2 _18236_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[9][7] ),
    .Y(_05414_));
 sky130_fd_sc_hd__or2_2 _18237_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[9][7] ),
    .X(_05415_));
 sky130_fd_sc_hd__a211o_2 _18238_ (.A1(_05414_),
    .A2(_05415_),
    .B1(_05408_),
    .C1(_05412_),
    .X(_05416_));
 sky130_fd_sc_hd__o211ai_2 _18239_ (.A1(_05408_),
    .A2(_05412_),
    .B1(_05414_),
    .C1(_05415_),
    .Y(_05417_));
 sky130_fd_sc_hd__a32o_2 _18240_ (.A1(_11712_),
    .A2(_05416_),
    .A3(_05417_),
    .B1(\systolic_inst.acc_wires[9][7] ),
    .B2(_11258_),
    .X(_01369_));
 sky130_fd_sc_hd__or2_2 _18241_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[9][8] ),
    .X(_05418_));
 sky130_fd_sc_hd__nand2_2 _18242_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[9][8] ),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2_2 _18243_ (.A(_05418_),
    .B(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__nand3_2 _18244_ (.A(_05414_),
    .B(_05417_),
    .C(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21o_2 _18245_ (.A1(_05414_),
    .A2(_05417_),
    .B1(_05420_),
    .X(_05422_));
 sky130_fd_sc_hd__a32o_2 _18246_ (.A1(_11712_),
    .A2(_05421_),
    .A3(_05422_),
    .B1(\systolic_inst.acc_wires[9][8] ),
    .B2(_11258_),
    .X(_01370_));
 sky130_fd_sc_hd__nor2_2 _18247_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[9][9] ),
    .Y(_05423_));
 sky130_fd_sc_hd__nand2_2 _18248_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[9][9] ),
    .Y(_05424_));
 sky130_fd_sc_hd__and2b_2 _18249_ (.A_N(_05423_),
    .B(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__nand2_2 _18250_ (.A(_05419_),
    .B(_05422_),
    .Y(_05426_));
 sky130_fd_sc_hd__or2_2 _18251_ (.A(_05425_),
    .B(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__a21bo_2 _18252_ (.A1(_05419_),
    .A2(_05422_),
    .B1_N(_05425_),
    .X(_05428_));
 sky130_fd_sc_hd__a32o_2 _18253_ (.A1(_11712_),
    .A2(_05427_),
    .A3(_05428_),
    .B1(\systolic_inst.acc_wires[9][9] ),
    .B2(_11258_),
    .X(_01371_));
 sky130_fd_sc_hd__or2_2 _18254_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[9][10] ),
    .X(_05429_));
 sky130_fd_sc_hd__nand2_2 _18255_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[9][10] ),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_2 _18256_ (.A(_05429_),
    .B(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__a21o_2 _18257_ (.A1(_05424_),
    .A2(_05428_),
    .B1(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__nand3_2 _18258_ (.A(_05424_),
    .B(_05428_),
    .C(_05431_),
    .Y(_05433_));
 sky130_fd_sc_hd__a32o_2 _18259_ (.A1(_11712_),
    .A2(_05432_),
    .A3(_05433_),
    .B1(\systolic_inst.acc_wires[9][10] ),
    .B2(_11258_),
    .X(_01372_));
 sky130_fd_sc_hd__or2_2 _18260_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[9][11] ),
    .X(_05434_));
 sky130_fd_sc_hd__nand2_2 _18261_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[9][11] ),
    .Y(_05435_));
 sky130_fd_sc_hd__nand2_2 _18262_ (.A(_05434_),
    .B(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__a21oi_2 _18263_ (.A1(_05430_),
    .A2(_05432_),
    .B1(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__a31o_2 _18264_ (.A1(_05430_),
    .A2(_05432_),
    .A3(_05436_),
    .B1(_11713_),
    .X(_05438_));
 sky130_fd_sc_hd__a2bb2o_2 _18265_ (.A1_N(_05438_),
    .A2_N(_05437_),
    .B1(\systolic_inst.acc_wires[9][11] ),
    .B2(_11258_),
    .X(_01373_));
 sky130_fd_sc_hd__nor2_2 _18266_ (.A(_05431_),
    .B(_05436_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand2_2 _18267_ (.A(_05425_),
    .B(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__a211o_2 _18268_ (.A1(_05414_),
    .A2(_05417_),
    .B1(_05420_),
    .C1(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__o21ai_2 _18269_ (.A1(_05419_),
    .A2(_05423_),
    .B1(_05424_),
    .Y(_05442_));
 sky130_fd_sc_hd__and3_2 _18270_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[9][10] ),
    .C(_05434_),
    .X(_05443_));
 sky130_fd_sc_hd__a221oi_2 _18271_ (.A1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[11] ),
    .A2(\systolic_inst.acc_wires[9][11] ),
    .B1(_05439_),
    .B2(_05442_),
    .C1(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__and2_2 _18272_ (.A(_05441_),
    .B(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__or2_2 _18273_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[9][12] ),
    .X(_05446_));
 sky130_fd_sc_hd__nand2_2 _18274_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[9][12] ),
    .Y(_05447_));
 sky130_fd_sc_hd__nand2_2 _18275_ (.A(_05446_),
    .B(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__xor2_2 _18276_ (.A(_05445_),
    .B(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__a22o_2 _18277_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[9][12] ),
    .B1(_11712_),
    .B2(_05449_),
    .X(_01374_));
 sky130_fd_sc_hd__or2_2 _18278_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[9][13] ),
    .X(_05450_));
 sky130_fd_sc_hd__nand2_2 _18279_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[9][13] ),
    .Y(_05451_));
 sky130_fd_sc_hd__nand2_2 _18280_ (.A(_05450_),
    .B(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__o211a_2 _18281_ (.A1(_05445_),
    .A2(_05448_),
    .B1(_05452_),
    .C1(_05447_),
    .X(_05453_));
 sky130_fd_sc_hd__a211o_2 _18282_ (.A1(_05441_),
    .A2(_05444_),
    .B1(_05448_),
    .C1(_05452_),
    .X(_05454_));
 sky130_fd_sc_hd__o211ai_2 _18283_ (.A1(_05447_),
    .A2(_05452_),
    .B1(_05454_),
    .C1(_11712_),
    .Y(_05455_));
 sky130_fd_sc_hd__a2bb2o_2 _18284_ (.A1_N(_05455_),
    .A2_N(_05453_),
    .B1(\systolic_inst.acc_wires[9][13] ),
    .B2(_11258_),
    .X(_01375_));
 sky130_fd_sc_hd__or2_2 _18285_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[9][14] ),
    .X(_05456_));
 sky130_fd_sc_hd__nand2_2 _18286_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[9][14] ),
    .Y(_05457_));
 sky130_fd_sc_hd__nand2_2 _18287_ (.A(_05456_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__o21a_2 _18288_ (.A1(_05447_),
    .A2(_05452_),
    .B1(_05451_),
    .X(_05459_));
 sky130_fd_sc_hd__a21o_2 _18289_ (.A1(_05454_),
    .A2(_05459_),
    .B1(_05458_),
    .X(_05460_));
 sky130_fd_sc_hd__nand3_2 _18290_ (.A(_05454_),
    .B(_05458_),
    .C(_05459_),
    .Y(_05461_));
 sky130_fd_sc_hd__a32o_2 _18291_ (.A1(_11712_),
    .A2(_05460_),
    .A3(_05461_),
    .B1(\systolic_inst.acc_wires[9][14] ),
    .B2(_11258_),
    .X(_01376_));
 sky130_fd_sc_hd__nor2_2 _18292_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][15] ),
    .Y(_05462_));
 sky130_fd_sc_hd__and2_2 _18293_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][15] ),
    .X(_05463_));
 sky130_fd_sc_hd__or2_2 _18294_ (.A(_05462_),
    .B(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__a21oi_2 _18295_ (.A1(_05457_),
    .A2(_05460_),
    .B1(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__a31o_2 _18296_ (.A1(_05457_),
    .A2(_05460_),
    .A3(_05464_),
    .B1(_11713_),
    .X(_05466_));
 sky130_fd_sc_hd__a2bb2o_2 _18297_ (.A1_N(_05466_),
    .A2_N(_05465_),
    .B1(\systolic_inst.acc_wires[9][15] ),
    .B2(_11258_),
    .X(_01377_));
 sky130_fd_sc_hd__a211o_2 _18298_ (.A1(_05454_),
    .A2(_05459_),
    .B1(_05464_),
    .C1(_05458_),
    .X(_05467_));
 sky130_fd_sc_hd__o21ba_2 _18299_ (.A1(_05457_),
    .A2(_05462_),
    .B1_N(_05463_),
    .X(_05468_));
 sky130_fd_sc_hd__and2_2 _18300_ (.A(_05467_),
    .B(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__or2_2 _18301_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][16] ),
    .X(_05470_));
 sky130_fd_sc_hd__nand2_2 _18302_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][16] ),
    .Y(_05471_));
 sky130_fd_sc_hd__nand2_2 _18303_ (.A(_05470_),
    .B(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2_2 _18304_ (.A(_05469_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__nor2_2 _18305_ (.A(_05469_),
    .B(_05472_),
    .Y(_05474_));
 sky130_fd_sc_hd__nor2_2 _18306_ (.A(_11713_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__a22o_2 _18307_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[9][16] ),
    .B1(_05473_),
    .B2(_05475_),
    .X(_01378_));
 sky130_fd_sc_hd__xor2_2 _18308_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][17] ),
    .X(_05476_));
 sky130_fd_sc_hd__o21a_2 _18309_ (.A1(_05469_),
    .A2(_05472_),
    .B1(_05471_),
    .X(_05477_));
 sky130_fd_sc_hd__xnor2_2 _18310_ (.A(_05476_),
    .B(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__a22o_2 _18311_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[9][17] ),
    .B1(_11712_),
    .B2(_05478_),
    .X(_01379_));
 sky130_fd_sc_hd__or2_2 _18312_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][18] ),
    .X(_05479_));
 sky130_fd_sc_hd__nand2_2 _18313_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][18] ),
    .Y(_05480_));
 sky130_fd_sc_hd__nand2_2 _18314_ (.A(_05479_),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__o21ai_2 _18315_ (.A1(\systolic_inst.acc_wires[9][16] ),
    .A2(\systolic_inst.acc_wires[9][17] ),
    .B1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .Y(_05482_));
 sky130_fd_sc_hd__nand2_2 _18316_ (.A(_05474_),
    .B(_05476_),
    .Y(_05483_));
 sky130_fd_sc_hd__a21o_2 _18317_ (.A1(_05482_),
    .A2(_05483_),
    .B1(_05481_),
    .X(_05484_));
 sky130_fd_sc_hd__nand3_2 _18318_ (.A(_05481_),
    .B(_05482_),
    .C(_05483_),
    .Y(_05485_));
 sky130_fd_sc_hd__a32o_2 _18319_ (.A1(_11712_),
    .A2(_05484_),
    .A3(_05485_),
    .B1(\systolic_inst.acc_wires[9][18] ),
    .B2(_11258_),
    .X(_01380_));
 sky130_fd_sc_hd__xnor2_2 _18320_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][19] ),
    .Y(_05486_));
 sky130_fd_sc_hd__a21oi_2 _18321_ (.A1(_05480_),
    .A2(_05484_),
    .B1(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__a31o_2 _18322_ (.A1(_05480_),
    .A2(_05484_),
    .A3(_05486_),
    .B1(_11713_),
    .X(_05488_));
 sky130_fd_sc_hd__a2bb2o_2 _18323_ (.A1_N(_05488_),
    .A2_N(_05487_),
    .B1(\systolic_inst.acc_wires[9][19] ),
    .B2(_11258_),
    .X(_01381_));
 sky130_fd_sc_hd__or2_2 _18324_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][20] ),
    .X(_05489_));
 sky130_fd_sc_hd__nand2_2 _18325_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][20] ),
    .Y(_05490_));
 sky130_fd_sc_hd__and2_2 _18326_ (.A(_05489_),
    .B(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__and3_2 _18327_ (.A(_05470_),
    .B(_05471_),
    .C(_05476_),
    .X(_05492_));
 sky130_fd_sc_hd__or3b_2 _18328_ (.A(_05481_),
    .B(_05486_),
    .C_N(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__nor2_2 _18329_ (.A(_05469_),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__o41a_2 _18330_ (.A1(\systolic_inst.acc_wires[9][16] ),
    .A2(\systolic_inst.acc_wires[9][17] ),
    .A3(\systolic_inst.acc_wires[9][18] ),
    .A4(\systolic_inst.acc_wires[9][19] ),
    .B1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .X(_05495_));
 sky130_fd_sc_hd__or3_2 _18331_ (.A(_05491_),
    .B(_05494_),
    .C(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__o21ai_2 _18332_ (.A1(_05494_),
    .A2(_05495_),
    .B1(_05491_),
    .Y(_05497_));
 sky130_fd_sc_hd__a32o_2 _18333_ (.A1(_11712_),
    .A2(_05496_),
    .A3(_05497_),
    .B1(\systolic_inst.acc_wires[9][20] ),
    .B2(_11258_),
    .X(_01382_));
 sky130_fd_sc_hd__xnor2_2 _18334_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][21] ),
    .Y(_05498_));
 sky130_fd_sc_hd__inv_2 _18335_ (.A(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__a21oi_2 _18336_ (.A1(_05490_),
    .A2(_05497_),
    .B1(_05498_),
    .Y(_05500_));
 sky130_fd_sc_hd__a31o_2 _18337_ (.A1(_05490_),
    .A2(_05497_),
    .A3(_05498_),
    .B1(_11713_),
    .X(_05501_));
 sky130_fd_sc_hd__a2bb2o_2 _18338_ (.A1_N(_05501_),
    .A2_N(_05500_),
    .B1(\systolic_inst.acc_wires[9][21] ),
    .B2(_11258_),
    .X(_01383_));
 sky130_fd_sc_hd__or2_2 _18339_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][22] ),
    .X(_05502_));
 sky130_fd_sc_hd__nand2_2 _18340_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][22] ),
    .Y(_05503_));
 sky130_fd_sc_hd__and2_2 _18341_ (.A(_05502_),
    .B(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__o21a_2 _18342_ (.A1(\systolic_inst.acc_wires[9][20] ),
    .A2(\systolic_inst.acc_wires[9][21] ),
    .B1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .X(_05505_));
 sky130_fd_sc_hd__nor2_2 _18343_ (.A(_05497_),
    .B(_05498_),
    .Y(_05506_));
 sky130_fd_sc_hd__o21ai_2 _18344_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_05504_),
    .Y(_05507_));
 sky130_fd_sc_hd__or3_2 _18345_ (.A(_05504_),
    .B(_05505_),
    .C(_05506_),
    .X(_05508_));
 sky130_fd_sc_hd__a32o_2 _18346_ (.A1(_11712_),
    .A2(_05507_),
    .A3(_05508_),
    .B1(\systolic_inst.acc_wires[9][22] ),
    .B2(_11258_),
    .X(_01384_));
 sky130_fd_sc_hd__xor2_2 _18347_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][23] ),
    .X(_05509_));
 sky130_fd_sc_hd__inv_2 _18348_ (.A(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__nand3_2 _18349_ (.A(_05503_),
    .B(_05507_),
    .C(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hd__a21o_2 _18350_ (.A1(_05503_),
    .A2(_05507_),
    .B1(_05510_),
    .X(_05512_));
 sky130_fd_sc_hd__a32o_2 _18351_ (.A1(_11712_),
    .A2(_05511_),
    .A3(_05512_),
    .B1(\systolic_inst.acc_wires[9][23] ),
    .B2(_11258_),
    .X(_01385_));
 sky130_fd_sc_hd__nand4_2 _18352_ (.A(_05491_),
    .B(_05499_),
    .C(_05504_),
    .D(_05509_),
    .Y(_05513_));
 sky130_fd_sc_hd__a211o_2 _18353_ (.A1(_05467_),
    .A2(_05468_),
    .B1(_05493_),
    .C1(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__o41a_2 _18354_ (.A1(\systolic_inst.acc_wires[9][20] ),
    .A2(\systolic_inst.acc_wires[9][21] ),
    .A3(\systolic_inst.acc_wires[9][22] ),
    .A4(\systolic_inst.acc_wires[9][23] ),
    .B1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .X(_05515_));
 sky130_fd_sc_hd__nor2_2 _18355_ (.A(_05495_),
    .B(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__nor2_2 _18356_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][24] ),
    .Y(_05517_));
 sky130_fd_sc_hd__and2_2 _18357_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][24] ),
    .X(_05518_));
 sky130_fd_sc_hd__or2_2 _18358_ (.A(_05517_),
    .B(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__a21oi_2 _18359_ (.A1(_05514_),
    .A2(_05516_),
    .B1(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__a31o_2 _18360_ (.A1(_05514_),
    .A2(_05516_),
    .A3(_05519_),
    .B1(_11713_),
    .X(_05521_));
 sky130_fd_sc_hd__a2bb2o_2 _18361_ (.A1_N(_05521_),
    .A2_N(_05520_),
    .B1(\systolic_inst.acc_wires[9][24] ),
    .B2(_11258_),
    .X(_01386_));
 sky130_fd_sc_hd__xor2_2 _18362_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][25] ),
    .X(_05522_));
 sky130_fd_sc_hd__or3_2 _18363_ (.A(_05518_),
    .B(_05520_),
    .C(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__o21ai_2 _18364_ (.A1(_05518_),
    .A2(_05520_),
    .B1(_05522_),
    .Y(_05524_));
 sky130_fd_sc_hd__a32o_2 _18365_ (.A1(_11712_),
    .A2(_05523_),
    .A3(_05524_),
    .B1(\systolic_inst.acc_wires[9][25] ),
    .B2(_11258_),
    .X(_01387_));
 sky130_fd_sc_hd__or2_2 _18366_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][26] ),
    .X(_05525_));
 sky130_fd_sc_hd__nand2_2 _18367_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][26] ),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_2 _18368_ (.A(_05525_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__o21a_2 _18369_ (.A1(\systolic_inst.acc_wires[9][24] ),
    .A2(\systolic_inst.acc_wires[9][25] ),
    .B1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .X(_05528_));
 sky130_fd_sc_hd__a21o_2 _18370_ (.A1(_05520_),
    .A2(_05522_),
    .B1(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__xnor2_2 _18371_ (.A(_05527_),
    .B(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__a22o_2 _18372_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[9][26] ),
    .B1(_11712_),
    .B2(_05530_),
    .X(_01388_));
 sky130_fd_sc_hd__xnor2_2 _18373_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][27] ),
    .Y(_05531_));
 sky130_fd_sc_hd__a21bo_2 _18374_ (.A1(_05525_),
    .A2(_05529_),
    .B1_N(_05526_),
    .X(_05532_));
 sky130_fd_sc_hd__xnor2_2 _18375_ (.A(_05531_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__a22o_2 _18376_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[9][27] ),
    .B1(_11712_),
    .B2(_05533_),
    .X(_01389_));
 sky130_fd_sc_hd__nor2_2 _18377_ (.A(_05527_),
    .B(_05531_),
    .Y(_05534_));
 sky130_fd_sc_hd__o21a_2 _18378_ (.A1(\systolic_inst.acc_wires[9][26] ),
    .A2(\systolic_inst.acc_wires[9][27] ),
    .B1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .X(_05535_));
 sky130_fd_sc_hd__a311oi_2 _18379_ (.A1(_05520_),
    .A2(_05522_),
    .A3(_05534_),
    .B1(_05535_),
    .C1(_05528_),
    .Y(_05536_));
 sky130_fd_sc_hd__or2_2 _18380_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][28] ),
    .X(_05537_));
 sky130_fd_sc_hd__nand2_2 _18381_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][28] ),
    .Y(_05538_));
 sky130_fd_sc_hd__nand2_2 _18382_ (.A(_05537_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__or2_2 _18383_ (.A(_05536_),
    .B(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__nand2_2 _18384_ (.A(_05536_),
    .B(_05539_),
    .Y(_05541_));
 sky130_fd_sc_hd__a32o_2 _18385_ (.A1(_11712_),
    .A2(_05540_),
    .A3(_05541_),
    .B1(\systolic_inst.acc_wires[9][28] ),
    .B2(_11258_),
    .X(_01390_));
 sky130_fd_sc_hd__xor2_2 _18386_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][29] ),
    .X(_05542_));
 sky130_fd_sc_hd__inv_2 _18387_ (.A(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__o21a_2 _18388_ (.A1(_05536_),
    .A2(_05539_),
    .B1(_05538_),
    .X(_05544_));
 sky130_fd_sc_hd__xnor2_2 _18389_ (.A(_05542_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__a22o_2 _18390_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[9][29] ),
    .B1(_11712_),
    .B2(_05545_),
    .X(_01391_));
 sky130_fd_sc_hd__o21ai_2 _18391_ (.A1(\systolic_inst.acc_wires[9][28] ),
    .A2(\systolic_inst.acc_wires[9][29] ),
    .B1(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .Y(_05546_));
 sky130_fd_sc_hd__o31a_2 _18392_ (.A1(_05536_),
    .A2(_05539_),
    .A3(_05543_),
    .B1(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__nand2_2 _18393_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][30] ),
    .Y(_05548_));
 sky130_fd_sc_hd__or2_2 _18394_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][30] ),
    .X(_05549_));
 sky130_fd_sc_hd__nand2_2 _18395_ (.A(_05548_),
    .B(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__nand2_2 _18396_ (.A(_05547_),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__or2_2 _18397_ (.A(_05547_),
    .B(_05550_),
    .X(_05552_));
 sky130_fd_sc_hd__a32o_2 _18398_ (.A1(_11712_),
    .A2(_05551_),
    .A3(_05552_),
    .B1(\systolic_inst.acc_wires[9][30] ),
    .B2(_11258_),
    .X(_01392_));
 sky130_fd_sc_hd__xnor2_2 _18399_ (.A(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[9][31] ),
    .Y(_05553_));
 sky130_fd_sc_hd__a21oi_2 _18400_ (.A1(_05548_),
    .A2(_05552_),
    .B1(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__a31o_2 _18401_ (.A1(_05548_),
    .A2(_05552_),
    .A3(_05553_),
    .B1(_11713_),
    .X(_05555_));
 sky130_fd_sc_hd__a2bb2o_2 _18402_ (.A1_N(_05555_),
    .A2_N(_05554_),
    .B1(\systolic_inst.acc_wires[9][31] ),
    .B2(_11258_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _18403_ (.A0(\systolic_inst.A_outs[8][0] ),
    .A1(\systolic_inst.A_shift[16][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _18404_ (.A0(\systolic_inst.A_outs[8][1] ),
    .A1(\systolic_inst.A_shift[16][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _18405_ (.A0(\systolic_inst.A_outs[8][2] ),
    .A1(\systolic_inst.A_shift[16][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _18406_ (.A0(\systolic_inst.A_outs[8][3] ),
    .A1(\systolic_inst.A_shift[16][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _18407_ (.A0(\systolic_inst.A_outs[8][4] ),
    .A1(\systolic_inst.A_shift[16][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _18408_ (.A0(\systolic_inst.A_outs[8][5] ),
    .A1(\systolic_inst.A_shift[16][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _18409_ (.A0(\systolic_inst.A_outs[8][6] ),
    .A1(\systolic_inst.A_shift[16][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _18410_ (.A0(\systolic_inst.A_outs[8][7] ),
    .A1(\systolic_inst.A_shift[16][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _18411_ (.A0(\systolic_inst.B_outs[7][0] ),
    .A1(\systolic_inst.B_outs[3][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _18412_ (.A0(\systolic_inst.B_outs[7][1] ),
    .A1(\systolic_inst.B_outs[3][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _18413_ (.A0(\systolic_inst.B_outs[7][2] ),
    .A1(\systolic_inst.B_outs[3][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _18414_ (.A0(\systolic_inst.B_outs[7][3] ),
    .A1(\systolic_inst.B_outs[3][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _18415_ (.A0(\systolic_inst.B_outs[7][4] ),
    .A1(\systolic_inst.B_outs[3][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _18416_ (.A0(\systolic_inst.B_outs[7][5] ),
    .A1(\systolic_inst.B_outs[3][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _18417_ (.A0(\systolic_inst.B_outs[7][6] ),
    .A1(\systolic_inst.B_outs[3][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _18418_ (.A0(\systolic_inst.B_outs[7][7] ),
    .A1(\systolic_inst.B_outs[3][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01409_));
 sky130_fd_sc_hd__and3_2 _18419_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[8][0] ),
    .C(\systolic_inst.A_outs[8][0] ),
    .X(_05556_));
 sky130_fd_sc_hd__a21o_2 _18420_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[0] ),
    .B1(_05556_),
    .X(_01410_));
 sky130_fd_sc_hd__and4_2 _18421_ (.A(\systolic_inst.B_outs[8][0] ),
    .B(\systolic_inst.A_outs[8][0] ),
    .C(\systolic_inst.B_outs[8][1] ),
    .D(\systolic_inst.A_outs[8][1] ),
    .X(_05557_));
 sky130_fd_sc_hd__a22o_2 _18422_ (.A1(\systolic_inst.A_outs[8][0] ),
    .A2(\systolic_inst.B_outs[8][1] ),
    .B1(\systolic_inst.A_outs[8][1] ),
    .B2(\systolic_inst.B_outs[8][0] ),
    .X(_05558_));
 sky130_fd_sc_hd__nand2_2 _18423_ (.A(\systolic_inst.ce_local ),
    .B(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__a2bb2o_2 _18424_ (.A1_N(_05559_),
    .A2_N(_05557_),
    .B1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01411_));
 sky130_fd_sc_hd__and2_2 _18425_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[2] ),
    .X(_05560_));
 sky130_fd_sc_hd__a22oi_2 _18426_ (.A1(\systolic_inst.B_outs[8][1] ),
    .A2(\systolic_inst.A_outs[8][1] ),
    .B1(\systolic_inst.A_outs[8][2] ),
    .B2(\systolic_inst.B_outs[8][0] ),
    .Y(_05561_));
 sky130_fd_sc_hd__and4_2 _18427_ (.A(\systolic_inst.B_outs[8][0] ),
    .B(\systolic_inst.B_outs[8][1] ),
    .C(\systolic_inst.A_outs[8][1] ),
    .D(\systolic_inst.A_outs[8][2] ),
    .X(_05562_));
 sky130_fd_sc_hd__or2_2 _18428_ (.A(_05561_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__or3b_2 _18429_ (.A(_05561_),
    .B(_05562_),
    .C_N(_05557_),
    .X(_05564_));
 sky130_fd_sc_hd__xnor2_2 _18430_ (.A(_05557_),
    .B(_05563_),
    .Y(_05565_));
 sky130_fd_sc_hd__nand3_2 _18431_ (.A(\systolic_inst.A_outs[8][0] ),
    .B(\systolic_inst.B_outs[8][2] ),
    .C(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__a21o_2 _18432_ (.A1(\systolic_inst.A_outs[8][0] ),
    .A2(\systolic_inst.B_outs[8][2] ),
    .B1(_05565_),
    .X(_05567_));
 sky130_fd_sc_hd__a31o_2 _18433_ (.A1(\systolic_inst.ce_local ),
    .A2(_05566_),
    .A3(_05567_),
    .B1(_05560_),
    .X(_01412_));
 sky130_fd_sc_hd__a22oi_2 _18434_ (.A1(\systolic_inst.A_outs[8][1] ),
    .A2(\systolic_inst.B_outs[8][2] ),
    .B1(\systolic_inst.B_outs[8][3] ),
    .B2(\systolic_inst.A_outs[8][0] ),
    .Y(_05568_));
 sky130_fd_sc_hd__and4_2 _18435_ (.A(\systolic_inst.A_outs[8][0] ),
    .B(\systolic_inst.A_outs[8][1] ),
    .C(\systolic_inst.B_outs[8][2] ),
    .D(\systolic_inst.B_outs[8][3] ),
    .X(_05569_));
 sky130_fd_sc_hd__nor2_2 _18436_ (.A(_05568_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__a22o_2 _18437_ (.A1(\systolic_inst.B_outs[8][1] ),
    .A2(\systolic_inst.A_outs[8][2] ),
    .B1(\systolic_inst.A_outs[8][3] ),
    .B2(\systolic_inst.B_outs[8][0] ),
    .X(_05571_));
 sky130_fd_sc_hd__nand4_2 _18438_ (.A(\systolic_inst.B_outs[8][0] ),
    .B(\systolic_inst.B_outs[8][1] ),
    .C(\systolic_inst.A_outs[8][2] ),
    .D(\systolic_inst.A_outs[8][3] ),
    .Y(_05572_));
 sky130_fd_sc_hd__nand3_2 _18439_ (.A(_05562_),
    .B(_05571_),
    .C(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__a21o_2 _18440_ (.A1(_05571_),
    .A2(_05572_),
    .B1(_05562_),
    .X(_05574_));
 sky130_fd_sc_hd__and2_2 _18441_ (.A(_05573_),
    .B(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__nand2_2 _18442_ (.A(_05570_),
    .B(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__xnor2_2 _18443_ (.A(_05570_),
    .B(_05575_),
    .Y(_05577_));
 sky130_fd_sc_hd__and3_2 _18444_ (.A(_05564_),
    .B(_05566_),
    .C(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__a21oi_2 _18445_ (.A1(_05564_),
    .A2(_05566_),
    .B1(_05577_),
    .Y(_05579_));
 sky130_fd_sc_hd__nand2_2 _18446_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[3] ),
    .Y(_05580_));
 sky130_fd_sc_hd__o31ai_2 _18447_ (.A1(_11258_),
    .A2(_05578_),
    .A3(_05579_),
    .B1(_05580_),
    .Y(_01413_));
 sky130_fd_sc_hd__and2_2 _18448_ (.A(\systolic_inst.B_outs[8][2] ),
    .B(\systolic_inst.A_outs[8][2] ),
    .X(_05581_));
 sky130_fd_sc_hd__nand4_2 _18449_ (.A(\systolic_inst.A_outs[8][0] ),
    .B(\systolic_inst.A_outs[8][1] ),
    .C(\systolic_inst.B_outs[8][3] ),
    .D(\systolic_inst.B_outs[8][4] ),
    .Y(_05582_));
 sky130_fd_sc_hd__a22o_2 _18450_ (.A1(\systolic_inst.A_outs[8][1] ),
    .A2(\systolic_inst.B_outs[8][3] ),
    .B1(\systolic_inst.B_outs[8][4] ),
    .B2(\systolic_inst.A_outs[8][0] ),
    .X(_05583_));
 sky130_fd_sc_hd__nand2_2 _18451_ (.A(_05582_),
    .B(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__xnor2_2 _18452_ (.A(_05581_),
    .B(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__a22o_2 _18453_ (.A1(\systolic_inst.B_outs[8][1] ),
    .A2(\systolic_inst.A_outs[8][3] ),
    .B1(\systolic_inst.A_outs[8][4] ),
    .B2(\systolic_inst.B_outs[8][0] ),
    .X(_05586_));
 sky130_fd_sc_hd__and3_2 _18454_ (.A(\systolic_inst.B_outs[8][0] ),
    .B(\systolic_inst.B_outs[8][1] ),
    .C(\systolic_inst.A_outs[8][3] ),
    .X(_05587_));
 sky130_fd_sc_hd__nand2_2 _18455_ (.A(\systolic_inst.A_outs[8][4] ),
    .B(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__and3_2 _18456_ (.A(_05569_),
    .B(_05586_),
    .C(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__a21oi_2 _18457_ (.A1(_05586_),
    .A2(_05588_),
    .B1(_05569_),
    .Y(_05590_));
 sky130_fd_sc_hd__nor3_2 _18458_ (.A(_05572_),
    .B(_05589_),
    .C(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__or3_2 _18459_ (.A(_05572_),
    .B(_05589_),
    .C(_05590_),
    .X(_05592_));
 sky130_fd_sc_hd__o21ai_2 _18460_ (.A1(_05589_),
    .A2(_05590_),
    .B1(_05572_),
    .Y(_05593_));
 sky130_fd_sc_hd__and3_2 _18461_ (.A(_05585_),
    .B(_05592_),
    .C(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__a21oi_2 _18462_ (.A1(_05592_),
    .A2(_05593_),
    .B1(_05585_),
    .Y(_05595_));
 sky130_fd_sc_hd__a211o_2 _18463_ (.A1(_05573_),
    .A2(_05576_),
    .B1(_05594_),
    .C1(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__o211ai_2 _18464_ (.A1(_05594_),
    .A2(_05595_),
    .B1(_05573_),
    .C1(_05576_),
    .Y(_05597_));
 sky130_fd_sc_hd__a21oi_2 _18465_ (.A1(_05596_),
    .A2(_05597_),
    .B1(_05579_),
    .Y(_05598_));
 sky130_fd_sc_hd__and3_2 _18466_ (.A(_05579_),
    .B(_05596_),
    .C(_05597_),
    .X(_05599_));
 sky130_fd_sc_hd__or3_2 _18467_ (.A(_11258_),
    .B(_05598_),
    .C(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__a21bo_2 _18468_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[4] ),
    .B1_N(_05600_),
    .X(_01414_));
 sky130_fd_sc_hd__a21bo_2 _18469_ (.A1(_05581_),
    .A2(_05583_),
    .B1_N(_05582_),
    .X(_05601_));
 sky130_fd_sc_hd__a22oi_2 _18470_ (.A1(\systolic_inst.B_outs[8][1] ),
    .A2(\systolic_inst.A_outs[8][4] ),
    .B1(\systolic_inst.A_outs[8][5] ),
    .B2(\systolic_inst.B_outs[8][0] ),
    .Y(_05602_));
 sky130_fd_sc_hd__and4_2 _18471_ (.A(\systolic_inst.B_outs[8][0] ),
    .B(\systolic_inst.B_outs[8][1] ),
    .C(\systolic_inst.A_outs[8][4] ),
    .D(\systolic_inst.A_outs[8][5] ),
    .X(_05603_));
 sky130_fd_sc_hd__nor2_2 _18472_ (.A(_05602_),
    .B(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__xor2_2 _18473_ (.A(_05601_),
    .B(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__xor2_2 _18474_ (.A(_05588_),
    .B(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__and4_2 _18475_ (.A(\systolic_inst.A_outs[8][1] ),
    .B(\systolic_inst.A_outs[8][2] ),
    .C(\systolic_inst.B_outs[8][3] ),
    .D(\systolic_inst.B_outs[8][4] ),
    .X(_05607_));
 sky130_fd_sc_hd__a22oi_2 _18476_ (.A1(\systolic_inst.A_outs[8][2] ),
    .A2(\systolic_inst.B_outs[8][3] ),
    .B1(\systolic_inst.B_outs[8][4] ),
    .B2(\systolic_inst.A_outs[8][1] ),
    .Y(_05608_));
 sky130_fd_sc_hd__a22o_2 _18477_ (.A1(\systolic_inst.A_outs[8][2] ),
    .A2(\systolic_inst.B_outs[8][3] ),
    .B1(\systolic_inst.B_outs[8][4] ),
    .B2(\systolic_inst.A_outs[8][1] ),
    .X(_05609_));
 sky130_fd_sc_hd__and4b_2 _18478_ (.A_N(_05607_),
    .B(_05609_),
    .C(\systolic_inst.B_outs[8][2] ),
    .D(\systolic_inst.A_outs[8][3] ),
    .X(_05610_));
 sky130_fd_sc_hd__o2bb2a_2 _18479_ (.A1_N(\systolic_inst.B_outs[8][2] ),
    .A2_N(\systolic_inst.A_outs[8][3] ),
    .B1(_05607_),
    .B2(_05608_),
    .X(_05611_));
 sky130_fd_sc_hd__and4bb_2 _18480_ (.A_N(_05610_),
    .B_N(_05611_),
    .C(\systolic_inst.A_outs[8][0] ),
    .D(\systolic_inst.B_outs[8][5] ),
    .X(_05612_));
 sky130_fd_sc_hd__o2bb2a_2 _18481_ (.A1_N(\systolic_inst.A_outs[8][0] ),
    .A2_N(\systolic_inst.B_outs[8][5] ),
    .B1(_05610_),
    .B2(_05611_),
    .X(_05613_));
 sky130_fd_sc_hd__or2_2 _18482_ (.A(_05612_),
    .B(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__nor2_2 _18483_ (.A(_05606_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__xor2_2 _18484_ (.A(_05606_),
    .B(_05614_),
    .X(_05616_));
 sky130_fd_sc_hd__nand2_2 _18485_ (.A(_05594_),
    .B(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hd__xor2_2 _18486_ (.A(_05594_),
    .B(_05616_),
    .X(_05618_));
 sky130_fd_sc_hd__o21ai_2 _18487_ (.A1(_05589_),
    .A2(_05591_),
    .B1(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__or3_2 _18488_ (.A(_05589_),
    .B(_05591_),
    .C(_05618_),
    .X(_05620_));
 sky130_fd_sc_hd__and2_2 _18489_ (.A(_05619_),
    .B(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__a21bo_2 _18490_ (.A1(_05579_),
    .A2(_05597_),
    .B1_N(_05596_),
    .X(_05622_));
 sky130_fd_sc_hd__nand2_2 _18491_ (.A(_05621_),
    .B(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__o21a_2 _18492_ (.A1(_05621_),
    .A2(_05622_),
    .B1(\systolic_inst.ce_local ),
    .X(_05624_));
 sky130_fd_sc_hd__a22o_2 _18493_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[5] ),
    .B1(_05623_),
    .B2(_05624_),
    .X(_01415_));
 sky130_fd_sc_hd__a32o_2 _18494_ (.A1(\systolic_inst.A_outs[8][4] ),
    .A2(_05587_),
    .A3(_05605_),
    .B1(_05604_),
    .B2(_05601_),
    .X(_05625_));
 sky130_fd_sc_hd__a31o_2 _18495_ (.A1(\systolic_inst.B_outs[8][2] ),
    .A2(\systolic_inst.A_outs[8][3] ),
    .A3(_05609_),
    .B1(_05607_),
    .X(_05626_));
 sky130_fd_sc_hd__a22oi_2 _18496_ (.A1(\systolic_inst.B_outs[8][1] ),
    .A2(\systolic_inst.A_outs[8][5] ),
    .B1(\systolic_inst.A_outs[8][6] ),
    .B2(\systolic_inst.B_outs[8][0] ),
    .Y(_05627_));
 sky130_fd_sc_hd__and4_2 _18497_ (.A(\systolic_inst.B_outs[8][0] ),
    .B(\systolic_inst.B_outs[8][1] ),
    .C(\systolic_inst.A_outs[8][5] ),
    .D(\systolic_inst.A_outs[8][6] ),
    .X(_05628_));
 sky130_fd_sc_hd__or2_2 _18498_ (.A(_05627_),
    .B(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__and2b_2 _18499_ (.A_N(_05629_),
    .B(_05626_),
    .X(_05630_));
 sky130_fd_sc_hd__xnor2_2 _18500_ (.A(_05626_),
    .B(_05629_),
    .Y(_05631_));
 sky130_fd_sc_hd__xor2_2 _18501_ (.A(_05603_),
    .B(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__nand4_2 _18502_ (.A(\systolic_inst.A_outs[8][2] ),
    .B(\systolic_inst.B_outs[8][3] ),
    .C(\systolic_inst.A_outs[8][3] ),
    .D(\systolic_inst.B_outs[8][4] ),
    .Y(_05633_));
 sky130_fd_sc_hd__a22o_2 _18503_ (.A1(\systolic_inst.B_outs[8][3] ),
    .A2(\systolic_inst.A_outs[8][3] ),
    .B1(\systolic_inst.B_outs[8][4] ),
    .B2(\systolic_inst.A_outs[8][2] ),
    .X(_05634_));
 sky130_fd_sc_hd__nand4_2 _18504_ (.A(\systolic_inst.B_outs[8][2] ),
    .B(\systolic_inst.A_outs[8][4] ),
    .C(_05633_),
    .D(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__a22o_2 _18505_ (.A1(\systolic_inst.B_outs[8][2] ),
    .A2(\systolic_inst.A_outs[8][4] ),
    .B1(_05633_),
    .B2(_05634_),
    .X(_05636_));
 sky130_fd_sc_hd__a22oi_2 _18506_ (.A1(\systolic_inst.A_outs[8][1] ),
    .A2(\systolic_inst.B_outs[8][5] ),
    .B1(\systolic_inst.B_outs[8][6] ),
    .B2(\systolic_inst.A_outs[8][0] ),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_2 _18507_ (.A(\systolic_inst.A_outs[8][1] ),
    .B(\systolic_inst.B_outs[8][6] ),
    .Y(_05638_));
 sky130_fd_sc_hd__and4_2 _18508_ (.A(\systolic_inst.A_outs[8][0] ),
    .B(\systolic_inst.A_outs[8][1] ),
    .C(\systolic_inst.B_outs[8][5] ),
    .D(\systolic_inst.B_outs[8][6] ),
    .X(_05639_));
 sky130_fd_sc_hd__nor2_2 _18509_ (.A(_05637_),
    .B(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__nand3_2 _18510_ (.A(_05635_),
    .B(_05636_),
    .C(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__a21o_2 _18511_ (.A1(_05635_),
    .A2(_05636_),
    .B1(_05640_),
    .X(_05642_));
 sky130_fd_sc_hd__and3_2 _18512_ (.A(_05612_),
    .B(_05641_),
    .C(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__a21oi_2 _18513_ (.A1(_05641_),
    .A2(_05642_),
    .B1(_05612_),
    .Y(_05644_));
 sky130_fd_sc_hd__or3b_2 _18514_ (.A(_05643_),
    .B(_05644_),
    .C_N(_05632_),
    .X(_05645_));
 sky130_fd_sc_hd__o21bai_2 _18515_ (.A1(_05643_),
    .A2(_05644_),
    .B1_N(_05632_),
    .Y(_05646_));
 sky130_fd_sc_hd__nand3_2 _18516_ (.A(_05615_),
    .B(_05645_),
    .C(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__a21o_2 _18517_ (.A1(_05645_),
    .A2(_05646_),
    .B1(_05615_),
    .X(_05648_));
 sky130_fd_sc_hd__and3_2 _18518_ (.A(_05625_),
    .B(_05647_),
    .C(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__a21oi_2 _18519_ (.A1(_05647_),
    .A2(_05648_),
    .B1(_05625_),
    .Y(_05650_));
 sky130_fd_sc_hd__a211oi_2 _18520_ (.A1(_05617_),
    .A2(_05619_),
    .B1(_05649_),
    .C1(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__o211a_2 _18521_ (.A1(_05649_),
    .A2(_05650_),
    .B1(_05617_),
    .C1(_05619_),
    .X(_05652_));
 sky130_fd_sc_hd__nor2_2 _18522_ (.A(_05651_),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__xnor2_2 _18523_ (.A(_05623_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__mux2_1 _18524_ (.A0(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[6] ),
    .A1(_05654_),
    .S(\systolic_inst.ce_local ),
    .X(_01416_));
 sky130_fd_sc_hd__a21boi_2 _18525_ (.A1(_05625_),
    .A2(_05648_),
    .B1_N(_05647_),
    .Y(_05655_));
 sky130_fd_sc_hd__a21oi_2 _18526_ (.A1(_05603_),
    .A2(_05631_),
    .B1(_05630_),
    .Y(_05656_));
 sky130_fd_sc_hd__nand2_2 _18527_ (.A(_05633_),
    .B(_05635_),
    .Y(_05657_));
 sky130_fd_sc_hd__a22o_2 _18528_ (.A1(\systolic_inst.B_outs[8][1] ),
    .A2(\systolic_inst.A_outs[8][6] ),
    .B1(\systolic_inst.A_outs[8][7] ),
    .B2(\systolic_inst.B_outs[8][0] ),
    .X(_05658_));
 sky130_fd_sc_hd__nand4_2 _18529_ (.A(\systolic_inst.B_outs[8][0] ),
    .B(\systolic_inst.B_outs[8][1] ),
    .C(\systolic_inst.A_outs[8][6] ),
    .D(\systolic_inst.A_outs[8][7] ),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2_2 _18530_ (.A(_05658_),
    .B(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__xnor2_2 _18531_ (.A(_11259_),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__nand2b_2 _18532_ (.A_N(_05661_),
    .B(_05657_),
    .Y(_05662_));
 sky130_fd_sc_hd__xnor2_2 _18533_ (.A(_05657_),
    .B(_05661_),
    .Y(_05663_));
 sky130_fd_sc_hd__xnor2_2 _18534_ (.A(_05628_),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__nand2_2 _18535_ (.A(\systolic_inst.B_outs[8][2] ),
    .B(\systolic_inst.A_outs[8][5] ),
    .Y(_05665_));
 sky130_fd_sc_hd__and4_2 _18536_ (.A(\systolic_inst.B_outs[8][3] ),
    .B(\systolic_inst.A_outs[8][3] ),
    .C(\systolic_inst.B_outs[8][4] ),
    .D(\systolic_inst.A_outs[8][4] ),
    .X(_05666_));
 sky130_fd_sc_hd__a22oi_2 _18537_ (.A1(\systolic_inst.A_outs[8][3] ),
    .A2(\systolic_inst.B_outs[8][4] ),
    .B1(\systolic_inst.A_outs[8][4] ),
    .B2(\systolic_inst.B_outs[8][3] ),
    .Y(_05667_));
 sky130_fd_sc_hd__or2_2 _18538_ (.A(_05666_),
    .B(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__xnor2_2 _18539_ (.A(_05665_),
    .B(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__nand2_2 _18540_ (.A(\systolic_inst.A_outs[8][2] ),
    .B(\systolic_inst.B_outs[8][5] ),
    .Y(_05670_));
 sky130_fd_sc_hd__and2b_2 _18541_ (.A_N(\systolic_inst.A_outs[8][0] ),
    .B(\systolic_inst.B_outs[8][7] ),
    .X(_05671_));
 sky130_fd_sc_hd__and3_2 _18542_ (.A(\systolic_inst.A_outs[8][1] ),
    .B(\systolic_inst.B_outs[8][6] ),
    .C(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__xnor2_2 _18543_ (.A(_05638_),
    .B(_05671_),
    .Y(_05673_));
 sky130_fd_sc_hd__xnor2_2 _18544_ (.A(_05670_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__xnor2_2 _18545_ (.A(_05639_),
    .B(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__nor2_2 _18546_ (.A(_05669_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__xnor2_2 _18547_ (.A(_05669_),
    .B(_05675_),
    .Y(_05677_));
 sky130_fd_sc_hd__or2_2 _18548_ (.A(_05641_),
    .B(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__and2_2 _18549_ (.A(_05641_),
    .B(_05677_),
    .X(_05679_));
 sky130_fd_sc_hd__xor2_2 _18550_ (.A(_05641_),
    .B(_05677_),
    .X(_05680_));
 sky130_fd_sc_hd__xnor2_2 _18551_ (.A(_05664_),
    .B(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__and2b_2 _18552_ (.A_N(_05643_),
    .B(_05645_),
    .X(_05682_));
 sky130_fd_sc_hd__nand2b_2 _18553_ (.A_N(_05682_),
    .B(_05681_),
    .Y(_05683_));
 sky130_fd_sc_hd__xnor2_2 _18554_ (.A(_05681_),
    .B(_05682_),
    .Y(_05684_));
 sky130_fd_sc_hd__nand2b_2 _18555_ (.A_N(_05656_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__xnor2_2 _18556_ (.A(_05656_),
    .B(_05684_),
    .Y(_05686_));
 sky130_fd_sc_hd__and2b_2 _18557_ (.A_N(_05655_),
    .B(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__xnor2_2 _18558_ (.A(_05655_),
    .B(_05686_),
    .Y(_05688_));
 sky130_fd_sc_hd__a31o_2 _18559_ (.A1(_05621_),
    .A2(_05622_),
    .A3(_05653_),
    .B1(_05651_),
    .X(_05689_));
 sky130_fd_sc_hd__xor2_2 _18560_ (.A(_05688_),
    .B(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__mux2_1 _18561_ (.A0(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[7] ),
    .A1(_05690_),
    .S(\systolic_inst.ce_local ),
    .X(_01417_));
 sky130_fd_sc_hd__a21bo_2 _18562_ (.A1(_05628_),
    .A2(_05663_),
    .B1_N(_05662_),
    .X(_05691_));
 sky130_fd_sc_hd__a21bo_2 _18563_ (.A1(\systolic_inst.B_outs[8][7] ),
    .A2(_05658_),
    .B1_N(_05659_),
    .X(_05692_));
 sky130_fd_sc_hd__o21bai_2 _18564_ (.A1(_05665_),
    .A2(_05667_),
    .B1_N(_05666_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21a_2 _18565_ (.A1(\systolic_inst.B_outs[8][0] ),
    .A2(\systolic_inst.B_outs[8][1] ),
    .B1(\systolic_inst.A_outs[8][7] ),
    .X(_05694_));
 sky130_fd_sc_hd__o21ai_2 _18566_ (.A1(\systolic_inst.B_outs[8][0] ),
    .A2(\systolic_inst.B_outs[8][1] ),
    .B1(\systolic_inst.A_outs[8][7] ),
    .Y(_05695_));
 sky130_fd_sc_hd__a21o_2 _18567_ (.A1(\systolic_inst.B_outs[8][0] ),
    .A2(\systolic_inst.B_outs[8][1] ),
    .B1(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__and2b_2 _18568_ (.A_N(_05696_),
    .B(_05693_),
    .X(_05697_));
 sky130_fd_sc_hd__xnor2_2 _18569_ (.A(_05693_),
    .B(_05696_),
    .Y(_05698_));
 sky130_fd_sc_hd__xnor2_2 _18570_ (.A(_05692_),
    .B(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__and4_2 _18571_ (.A(\systolic_inst.B_outs[8][3] ),
    .B(\systolic_inst.B_outs[8][4] ),
    .C(\systolic_inst.A_outs[8][4] ),
    .D(\systolic_inst.A_outs[8][5] ),
    .X(_05700_));
 sky130_fd_sc_hd__a22oi_2 _18572_ (.A1(\systolic_inst.B_outs[8][4] ),
    .A2(\systolic_inst.A_outs[8][4] ),
    .B1(\systolic_inst.A_outs[8][5] ),
    .B2(\systolic_inst.B_outs[8][3] ),
    .Y(_05701_));
 sky130_fd_sc_hd__nor2_2 _18573_ (.A(_05700_),
    .B(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__nand2_2 _18574_ (.A(\systolic_inst.B_outs[8][2] ),
    .B(\systolic_inst.A_outs[8][6] ),
    .Y(_05703_));
 sky130_fd_sc_hd__xnor2_2 _18575_ (.A(_05702_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__nand2_2 _18576_ (.A(\systolic_inst.A_outs[8][3] ),
    .B(\systolic_inst.B_outs[8][5] ),
    .Y(_05705_));
 sky130_fd_sc_hd__and4b_2 _18577_ (.A_N(\systolic_inst.A_outs[8][1] ),
    .B(\systolic_inst.A_outs[8][2] ),
    .C(\systolic_inst.B_outs[8][6] ),
    .D(\systolic_inst.B_outs[8][7] ),
    .X(_05706_));
 sky130_fd_sc_hd__a2bb2o_2 _18578_ (.A1_N(\systolic_inst.A_outs[8][1] ),
    .A2_N(_11259_),
    .B1(\systolic_inst.B_outs[8][6] ),
    .B2(\systolic_inst.A_outs[8][2] ),
    .X(_05707_));
 sky130_fd_sc_hd__and2b_2 _18579_ (.A_N(_05706_),
    .B(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__xnor2_2 _18580_ (.A(_05705_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__a31o_2 _18581_ (.A1(\systolic_inst.A_outs[8][2] ),
    .A2(\systolic_inst.B_outs[8][5] ),
    .A3(_05673_),
    .B1(_05672_),
    .X(_05710_));
 sky130_fd_sc_hd__and2_2 _18582_ (.A(_05709_),
    .B(_05710_),
    .X(_05711_));
 sky130_fd_sc_hd__xor2_2 _18583_ (.A(_05709_),
    .B(_05710_),
    .X(_05712_));
 sky130_fd_sc_hd__xor2_2 _18584_ (.A(_05704_),
    .B(_05712_),
    .X(_05713_));
 sky130_fd_sc_hd__a21oi_2 _18585_ (.A1(_05639_),
    .A2(_05674_),
    .B1(_05676_),
    .Y(_05714_));
 sky130_fd_sc_hd__and2b_2 _18586_ (.A_N(_05714_),
    .B(_05713_),
    .X(_05715_));
 sky130_fd_sc_hd__xor2_2 _18587_ (.A(_05713_),
    .B(_05714_),
    .X(_05716_));
 sky130_fd_sc_hd__xor2_2 _18588_ (.A(_05699_),
    .B(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__o21a_2 _18589_ (.A1(_05664_),
    .A2(_05679_),
    .B1(_05678_),
    .X(_05718_));
 sky130_fd_sc_hd__nand2b_2 _18590_ (.A_N(_05718_),
    .B(_05717_),
    .Y(_05719_));
 sky130_fd_sc_hd__xor2_2 _18591_ (.A(_05717_),
    .B(_05718_),
    .X(_05720_));
 sky130_fd_sc_hd__nand2b_2 _18592_ (.A_N(_05720_),
    .B(_05691_),
    .Y(_05721_));
 sky130_fd_sc_hd__xor2_2 _18593_ (.A(_05691_),
    .B(_05720_),
    .X(_05722_));
 sky130_fd_sc_hd__and2_2 _18594_ (.A(_05683_),
    .B(_05685_),
    .X(_05723_));
 sky130_fd_sc_hd__or2_2 _18595_ (.A(_05722_),
    .B(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__xor2_2 _18596_ (.A(_05722_),
    .B(_05723_),
    .X(_05725_));
 sky130_fd_sc_hd__a21o_2 _18597_ (.A1(_05688_),
    .A2(_05689_),
    .B1(_05687_),
    .X(_05726_));
 sky130_fd_sc_hd__nand2_2 _18598_ (.A(_05725_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__or2_2 _18599_ (.A(_05725_),
    .B(_05726_),
    .X(_05728_));
 sky130_fd_sc_hd__and2_2 _18600_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[8] ),
    .X(_05729_));
 sky130_fd_sc_hd__a31o_2 _18601_ (.A1(\systolic_inst.ce_local ),
    .A2(_05727_),
    .A3(_05728_),
    .B1(_05729_),
    .X(_01418_));
 sky130_fd_sc_hd__a21o_2 _18602_ (.A1(_05692_),
    .A2(_05698_),
    .B1(_05697_),
    .X(_05730_));
 sky130_fd_sc_hd__o21ba_2 _18603_ (.A1(_05701_),
    .A2(_05703_),
    .B1_N(_05700_),
    .X(_05731_));
 sky130_fd_sc_hd__nor2_2 _18604_ (.A(_05695_),
    .B(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__and2_2 _18605_ (.A(_05695_),
    .B(_05731_),
    .X(_05733_));
 sky130_fd_sc_hd__or2_2 _18606_ (.A(_05732_),
    .B(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__nand2_2 _18607_ (.A(\systolic_inst.B_outs[8][2] ),
    .B(\systolic_inst.A_outs[8][7] ),
    .Y(_05735_));
 sky130_fd_sc_hd__a22oi_2 _18608_ (.A1(\systolic_inst.B_outs[8][4] ),
    .A2(\systolic_inst.A_outs[8][5] ),
    .B1(\systolic_inst.A_outs[8][6] ),
    .B2(\systolic_inst.B_outs[8][3] ),
    .Y(_05736_));
 sky130_fd_sc_hd__and4_2 _18609_ (.A(\systolic_inst.B_outs[8][3] ),
    .B(\systolic_inst.B_outs[8][4] ),
    .C(\systolic_inst.A_outs[8][5] ),
    .D(\systolic_inst.A_outs[8][6] ),
    .X(_05737_));
 sky130_fd_sc_hd__nor2_2 _18610_ (.A(_05736_),
    .B(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__xnor2_2 _18611_ (.A(_05735_),
    .B(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__nand2_2 _18612_ (.A(\systolic_inst.B_outs[8][5] ),
    .B(\systolic_inst.A_outs[8][4] ),
    .Y(_05740_));
 sky130_fd_sc_hd__and4b_2 _18613_ (.A_N(\systolic_inst.A_outs[8][2] ),
    .B(\systolic_inst.A_outs[8][3] ),
    .C(\systolic_inst.B_outs[8][6] ),
    .D(\systolic_inst.B_outs[8][7] ),
    .X(_05741_));
 sky130_fd_sc_hd__o2bb2a_2 _18614_ (.A1_N(\systolic_inst.A_outs[8][3] ),
    .A2_N(\systolic_inst.B_outs[8][6] ),
    .B1(_11259_),
    .B2(\systolic_inst.A_outs[8][2] ),
    .X(_05742_));
 sky130_fd_sc_hd__nor2_2 _18615_ (.A(_05741_),
    .B(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__xnor2_2 _18616_ (.A(_05740_),
    .B(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__a31oi_2 _18617_ (.A1(\systolic_inst.A_outs[8][3] ),
    .A2(\systolic_inst.B_outs[8][5] ),
    .A3(_05707_),
    .B1(_05706_),
    .Y(_05745_));
 sky130_fd_sc_hd__nand2b_2 _18618_ (.A_N(_05745_),
    .B(_05744_),
    .Y(_05746_));
 sky130_fd_sc_hd__xnor2_2 _18619_ (.A(_05744_),
    .B(_05745_),
    .Y(_05747_));
 sky130_fd_sc_hd__xnor2_2 _18620_ (.A(_05739_),
    .B(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__a21o_2 _18621_ (.A1(_05704_),
    .A2(_05712_),
    .B1(_05711_),
    .X(_05749_));
 sky130_fd_sc_hd__and2b_2 _18622_ (.A_N(_05748_),
    .B(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__xor2_2 _18623_ (.A(_05748_),
    .B(_05749_),
    .X(_05751_));
 sky130_fd_sc_hd__xor2_2 _18624_ (.A(_05734_),
    .B(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__o21ba_2 _18625_ (.A1(_05699_),
    .A2(_05716_),
    .B1_N(_05715_),
    .X(_05753_));
 sky130_fd_sc_hd__nand2b_2 _18626_ (.A_N(_05753_),
    .B(_05752_),
    .Y(_05754_));
 sky130_fd_sc_hd__xnor2_2 _18627_ (.A(_05752_),
    .B(_05753_),
    .Y(_05755_));
 sky130_fd_sc_hd__xnor2_2 _18628_ (.A(_05730_),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__a21o_2 _18629_ (.A1(_05719_),
    .A2(_05721_),
    .B1(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__and3_2 _18630_ (.A(_05719_),
    .B(_05721_),
    .C(_05756_),
    .X(_05758_));
 sky130_fd_sc_hd__inv_2 _18631_ (.A(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__nand2_2 _18632_ (.A(_05757_),
    .B(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__a21o_2 _18633_ (.A1(_05724_),
    .A2(_05727_),
    .B1(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__a31oi_2 _18634_ (.A1(_05724_),
    .A2(_05727_),
    .A3(_05760_),
    .B1(_11258_),
    .Y(_05762_));
 sky130_fd_sc_hd__a22o_2 _18635_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[9] ),
    .B1(_05761_),
    .B2(_05762_),
    .X(_01419_));
 sky130_fd_sc_hd__o21ba_2 _18636_ (.A1(_05735_),
    .A2(_05736_),
    .B1_N(_05737_),
    .X(_05763_));
 sky130_fd_sc_hd__nor2_2 _18637_ (.A(_05695_),
    .B(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__and2_2 _18638_ (.A(_05695_),
    .B(_05763_),
    .X(_05765_));
 sky130_fd_sc_hd__or2_2 _18639_ (.A(_05764_),
    .B(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__a22o_2 _18640_ (.A1(\systolic_inst.B_outs[8][4] ),
    .A2(\systolic_inst.A_outs[8][6] ),
    .B1(\systolic_inst.A_outs[8][7] ),
    .B2(\systolic_inst.B_outs[8][3] ),
    .X(_05767_));
 sky130_fd_sc_hd__and3_2 _18641_ (.A(\systolic_inst.B_outs[8][3] ),
    .B(\systolic_inst.B_outs[8][4] ),
    .C(\systolic_inst.A_outs[8][7] ),
    .X(_05768_));
 sky130_fd_sc_hd__a21bo_2 _18642_ (.A1(\systolic_inst.A_outs[8][6] ),
    .A2(_05768_),
    .B1_N(_05767_),
    .X(_05769_));
 sky130_fd_sc_hd__xor2_2 _18643_ (.A(_05735_),
    .B(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__nand2_2 _18644_ (.A(\systolic_inst.B_outs[8][5] ),
    .B(\systolic_inst.A_outs[8][5] ),
    .Y(_05771_));
 sky130_fd_sc_hd__and4b_2 _18645_ (.A_N(\systolic_inst.A_outs[8][3] ),
    .B(\systolic_inst.A_outs[8][4] ),
    .C(\systolic_inst.B_outs[8][6] ),
    .D(\systolic_inst.B_outs[8][7] ),
    .X(_05772_));
 sky130_fd_sc_hd__o2bb2a_2 _18646_ (.A1_N(\systolic_inst.A_outs[8][4] ),
    .A2_N(\systolic_inst.B_outs[8][6] ),
    .B1(_11259_),
    .B2(\systolic_inst.A_outs[8][3] ),
    .X(_05773_));
 sky130_fd_sc_hd__nor2_2 _18647_ (.A(_05772_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__xnor2_2 _18648_ (.A(_05771_),
    .B(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__o21ba_2 _18649_ (.A1(_05740_),
    .A2(_05742_),
    .B1_N(_05741_),
    .X(_05776_));
 sky130_fd_sc_hd__nand2b_2 _18650_ (.A_N(_05776_),
    .B(_05775_),
    .Y(_05777_));
 sky130_fd_sc_hd__xnor2_2 _18651_ (.A(_05775_),
    .B(_05776_),
    .Y(_05778_));
 sky130_fd_sc_hd__nand2_2 _18652_ (.A(_05770_),
    .B(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__or2_2 _18653_ (.A(_05770_),
    .B(_05778_),
    .X(_05780_));
 sky130_fd_sc_hd__nand2_2 _18654_ (.A(_05779_),
    .B(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__a21bo_2 _18655_ (.A1(_05739_),
    .A2(_05747_),
    .B1_N(_05746_),
    .X(_05782_));
 sky130_fd_sc_hd__nand2b_2 _18656_ (.A_N(_05781_),
    .B(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__xor2_2 _18657_ (.A(_05781_),
    .B(_05782_),
    .X(_05784_));
 sky130_fd_sc_hd__xor2_2 _18658_ (.A(_05766_),
    .B(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__o21ba_2 _18659_ (.A1(_05734_),
    .A2(_05751_),
    .B1_N(_05750_),
    .X(_05786_));
 sky130_fd_sc_hd__nand2b_2 _18660_ (.A_N(_05786_),
    .B(_05785_),
    .Y(_05787_));
 sky130_fd_sc_hd__xnor2_2 _18661_ (.A(_05785_),
    .B(_05786_),
    .Y(_05788_));
 sky130_fd_sc_hd__nand2_2 _18662_ (.A(_05732_),
    .B(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__xnor2_2 _18663_ (.A(_05732_),
    .B(_05788_),
    .Y(_05790_));
 sky130_fd_sc_hd__a21boi_2 _18664_ (.A1(_05730_),
    .A2(_05755_),
    .B1_N(_05754_),
    .Y(_05791_));
 sky130_fd_sc_hd__nor2_2 _18665_ (.A(_05790_),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__and2_2 _18666_ (.A(_05790_),
    .B(_05791_),
    .X(_05793_));
 sky130_fd_sc_hd__or2_2 _18667_ (.A(_05792_),
    .B(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__or3b_2 _18668_ (.A(_05758_),
    .B(_05727_),
    .C_N(_05757_),
    .X(_05795_));
 sky130_fd_sc_hd__a21o_2 _18669_ (.A1(_05724_),
    .A2(_05757_),
    .B1(_05758_),
    .X(_05796_));
 sky130_fd_sc_hd__a21oi_2 _18670_ (.A1(_05795_),
    .A2(_05796_),
    .B1(_05794_),
    .Y(_05797_));
 sky130_fd_sc_hd__and3_2 _18671_ (.A(_05794_),
    .B(_05795_),
    .C(_05796_),
    .X(_05798_));
 sky130_fd_sc_hd__nand2_2 _18672_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[10] ),
    .Y(_05799_));
 sky130_fd_sc_hd__o31ai_2 _18673_ (.A1(_11258_),
    .A2(_05797_),
    .A3(_05798_),
    .B1(_05799_),
    .Y(_01420_));
 sky130_fd_sc_hd__o2bb2a_2 _18674_ (.A1_N(\systolic_inst.A_outs[8][6] ),
    .A2_N(_05768_),
    .B1(_05769_),
    .B2(_05735_),
    .X(_05800_));
 sky130_fd_sc_hd__or2_2 _18675_ (.A(_05695_),
    .B(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__nand2_2 _18676_ (.A(_05695_),
    .B(_05800_),
    .Y(_05802_));
 sky130_fd_sc_hd__nand2_2 _18677_ (.A(_05801_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__or2_2 _18678_ (.A(\systolic_inst.B_outs[8][3] ),
    .B(\systolic_inst.B_outs[8][4] ),
    .X(_05804_));
 sky130_fd_sc_hd__and3b_2 _18679_ (.A_N(_05768_),
    .B(_05804_),
    .C(\systolic_inst.A_outs[8][7] ),
    .X(_05805_));
 sky130_fd_sc_hd__xnor2_2 _18680_ (.A(_05735_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__nand2_2 _18681_ (.A(\systolic_inst.B_outs[8][5] ),
    .B(\systolic_inst.A_outs[8][6] ),
    .Y(_05807_));
 sky130_fd_sc_hd__and4b_2 _18682_ (.A_N(\systolic_inst.A_outs[8][4] ),
    .B(\systolic_inst.A_outs[8][5] ),
    .C(\systolic_inst.B_outs[8][6] ),
    .D(\systolic_inst.B_outs[8][7] ),
    .X(_05808_));
 sky130_fd_sc_hd__o2bb2a_2 _18683_ (.A1_N(\systolic_inst.A_outs[8][5] ),
    .A2_N(\systolic_inst.B_outs[8][6] ),
    .B1(_11259_),
    .B2(\systolic_inst.A_outs[8][4] ),
    .X(_05809_));
 sky130_fd_sc_hd__or2_2 _18684_ (.A(_05808_),
    .B(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__xor2_2 _18685_ (.A(_05807_),
    .B(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__o21ba_2 _18686_ (.A1(_05771_),
    .A2(_05773_),
    .B1_N(_05772_),
    .X(_05812_));
 sky130_fd_sc_hd__nand2b_2 _18687_ (.A_N(_05812_),
    .B(_05811_),
    .Y(_05813_));
 sky130_fd_sc_hd__xnor2_2 _18688_ (.A(_05811_),
    .B(_05812_),
    .Y(_05814_));
 sky130_fd_sc_hd__nand2_2 _18689_ (.A(_05806_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__xnor2_2 _18690_ (.A(_05806_),
    .B(_05814_),
    .Y(_05816_));
 sky130_fd_sc_hd__a21o_2 _18691_ (.A1(_05777_),
    .A2(_05779_),
    .B1(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__nand3_2 _18692_ (.A(_05777_),
    .B(_05779_),
    .C(_05816_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_2 _18693_ (.A(_05817_),
    .B(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__xor2_2 _18694_ (.A(_05803_),
    .B(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__o21a_2 _18695_ (.A1(_05766_),
    .A2(_05784_),
    .B1(_05783_),
    .X(_05821_));
 sky130_fd_sc_hd__and2b_2 _18696_ (.A_N(_05821_),
    .B(_05820_),
    .X(_05822_));
 sky130_fd_sc_hd__xnor2_2 _18697_ (.A(_05820_),
    .B(_05821_),
    .Y(_05823_));
 sky130_fd_sc_hd__xnor2_2 _18698_ (.A(_05764_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__nand3_2 _18699_ (.A(_05787_),
    .B(_05789_),
    .C(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__inv_2 _18700_ (.A(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__a21oi_2 _18701_ (.A1(_05787_),
    .A2(_05789_),
    .B1(_05824_),
    .Y(_05827_));
 sky130_fd_sc_hd__nor2_2 _18702_ (.A(_05826_),
    .B(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__or3_2 _18703_ (.A(_05792_),
    .B(_05797_),
    .C(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__o21ai_2 _18704_ (.A1(_05792_),
    .A2(_05797_),
    .B1(_05828_),
    .Y(_05830_));
 sky130_fd_sc_hd__and2_2 _18705_ (.A(_11258_),
    .B(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[11] ),
    .X(_05831_));
 sky130_fd_sc_hd__a31o_2 _18706_ (.A1(\systolic_inst.ce_local ),
    .A2(_05829_),
    .A3(_05830_),
    .B1(_05831_),
    .X(_01421_));
 sky130_fd_sc_hd__a31o_2 _18707_ (.A1(\systolic_inst.B_outs[8][2] ),
    .A2(\systolic_inst.A_outs[8][7] ),
    .A3(_05804_),
    .B1(_05768_),
    .X(_05832_));
 sky130_fd_sc_hd__or2_2 _18708_ (.A(_05694_),
    .B(_05832_),
    .X(_05833_));
 sky130_fd_sc_hd__nand2_2 _18709_ (.A(_05694_),
    .B(_05832_),
    .Y(_05834_));
 sky130_fd_sc_hd__nand2_2 _18710_ (.A(_05833_),
    .B(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__o2bb2a_2 _18711_ (.A1_N(\systolic_inst.B_outs[8][6] ),
    .A2_N(\systolic_inst.A_outs[8][6] ),
    .B1(_11259_),
    .B2(\systolic_inst.A_outs[8][5] ),
    .X(_05836_));
 sky130_fd_sc_hd__and4b_2 _18712_ (.A_N(\systolic_inst.A_outs[8][5] ),
    .B(\systolic_inst.B_outs[8][6] ),
    .C(\systolic_inst.A_outs[8][6] ),
    .D(\systolic_inst.B_outs[8][7] ),
    .X(_05837_));
 sky130_fd_sc_hd__nor2_2 _18713_ (.A(_05836_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2_2 _18714_ (.A(\systolic_inst.B_outs[8][5] ),
    .B(\systolic_inst.A_outs[8][7] ),
    .Y(_05839_));
 sky130_fd_sc_hd__xnor2_2 _18715_ (.A(_05838_),
    .B(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__o21ba_2 _18716_ (.A1(_05807_),
    .A2(_05809_),
    .B1_N(_05808_),
    .X(_05841_));
 sky130_fd_sc_hd__nand2b_2 _18717_ (.A_N(_05841_),
    .B(_05840_),
    .Y(_05842_));
 sky130_fd_sc_hd__xnor2_2 _18718_ (.A(_05840_),
    .B(_05841_),
    .Y(_05843_));
 sky130_fd_sc_hd__xnor2_2 _18719_ (.A(_05806_),
    .B(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__a21o_2 _18720_ (.A1(_05813_),
    .A2(_05815_),
    .B1(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__nand3_2 _18721_ (.A(_05813_),
    .B(_05815_),
    .C(_05844_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_2 _18722_ (.A(_05845_),
    .B(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__xor2_2 _18723_ (.A(_05835_),
    .B(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__o21a_2 _18724_ (.A1(_05803_),
    .A2(_05819_),
    .B1(_05817_),
    .X(_05849_));
 sky130_fd_sc_hd__and2b_2 _18725_ (.A_N(_05849_),
    .B(_05848_),
    .X(_05850_));
 sky130_fd_sc_hd__xnor2_2 _18726_ (.A(_05848_),
    .B(_05849_),
    .Y(_05851_));
 sky130_fd_sc_hd__and2b_2 _18727_ (.A_N(_05801_),
    .B(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__xor2_2 _18728_ (.A(_05801_),
    .B(_05851_),
    .X(_05853_));
 sky130_fd_sc_hd__a21oi_2 _18729_ (.A1(_05764_),
    .A2(_05823_),
    .B1(_05822_),
    .Y(_05854_));
 sky130_fd_sc_hd__or2_2 _18730_ (.A(_05853_),
    .B(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__inv_2 _18731_ (.A(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_2 _18732_ (.A(_05853_),
    .B(_05854_),
    .Y(_05857_));
 sky130_fd_sc_hd__nand2_2 _18733_ (.A(_05855_),
    .B(_05857_),
    .Y(_05858_));
 sky130_fd_sc_hd__inv_2 _18734_ (.A(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__o31a_2 _18735_ (.A1(_05792_),
    .A2(_05797_),
    .A3(_05827_),
    .B1(_05825_),
    .X(_05860_));
 sky130_fd_sc_hd__o311a_2 _18736_ (.A1(_05792_),
    .A2(_05797_),
    .A3(_05827_),
    .B1(_05859_),
    .C1(_05825_),
    .X(_05861_));
 sky130_fd_sc_hd__nor2_2 _18737_ (.A(_05859_),
    .B(_05860_),
    .Y(_05862_));
 sky130_fd_sc_hd__nor2_2 _18738_ (.A(_05861_),
    .B(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__mux2_1 _18739_ (.A0(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[12] ),
    .A1(_05863_),
    .S(\systolic_inst.ce_local ),
    .X(_01422_));
 sky130_fd_sc_hd__nand2_2 _18740_ (.A(\systolic_inst.B_outs[8][6] ),
    .B(\systolic_inst.A_outs[8][7] ),
    .Y(_05864_));
 sky130_fd_sc_hd__or2_2 _18741_ (.A(\systolic_inst.A_outs[8][6] ),
    .B(_11259_),
    .X(_05865_));
 sky130_fd_sc_hd__and2_2 _18742_ (.A(_05864_),
    .B(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__nor2_2 _18743_ (.A(_05864_),
    .B(_05865_),
    .Y(_05867_));
 sky130_fd_sc_hd__nor2_2 _18744_ (.A(_05866_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__xnor2_2 _18745_ (.A(_05839_),
    .B(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__o21ba_2 _18746_ (.A1(_05836_),
    .A2(_05839_),
    .B1_N(_05837_),
    .X(_05870_));
 sky130_fd_sc_hd__nand2b_2 _18747_ (.A_N(_05870_),
    .B(_05869_),
    .Y(_05871_));
 sky130_fd_sc_hd__xnor2_2 _18748_ (.A(_05869_),
    .B(_05870_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand2_2 _18749_ (.A(_05806_),
    .B(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__or2_2 _18750_ (.A(_05806_),
    .B(_05872_),
    .X(_05874_));
 sky130_fd_sc_hd__nand2_2 _18751_ (.A(_05873_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__a21bo_2 _18752_ (.A1(_05806_),
    .A2(_05843_),
    .B1_N(_05842_),
    .X(_05876_));
 sky130_fd_sc_hd__nand2b_2 _18753_ (.A_N(_05875_),
    .B(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__xor2_2 _18754_ (.A(_05875_),
    .B(_05876_),
    .X(_05878_));
 sky130_fd_sc_hd__xor2_2 _18755_ (.A(_05835_),
    .B(_05878_),
    .X(_05879_));
 sky130_fd_sc_hd__o21a_2 _18756_ (.A1(_05835_),
    .A2(_05847_),
    .B1(_05845_),
    .X(_05880_));
 sky130_fd_sc_hd__and2b_2 _18757_ (.A_N(_05880_),
    .B(_05879_),
    .X(_05881_));
 sky130_fd_sc_hd__and2b_2 _18758_ (.A_N(_05879_),
    .B(_05880_),
    .X(_05882_));
 sky130_fd_sc_hd__nor2_2 _18759_ (.A(_05881_),
    .B(_05882_),
    .Y(_05883_));
 sky130_fd_sc_hd__xnor2_2 _18760_ (.A(_05834_),
    .B(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__o21a_2 _18761_ (.A1(_05850_),
    .A2(_05852_),
    .B1(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__nor3_2 _18762_ (.A(_05850_),
    .B(_05852_),
    .C(_05884_),
    .Y(_05886_));
 sky130_fd_sc_hd__inv_2 _18763_ (.A(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__nor2_2 _18764_ (.A(_05885_),
    .B(_05886_),
    .Y(_05888_));
 sky130_fd_sc_hd__or3_2 _18765_ (.A(_05856_),
    .B(_05861_),
    .C(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__o21ai_2 _18766_ (.A1(_05856_),
    .A2(_05861_),
    .B1(_05888_),
    .Y(_05890_));
 sky130_fd_sc_hd__and3_2 _18767_ (.A(\systolic_inst.ce_local ),
    .B(_05889_),
    .C(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__a21o_2 _18768_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[13] ),
    .B1(_05891_),
    .X(_01423_));
 sky130_fd_sc_hd__a31o_2 _18769_ (.A1(\systolic_inst.B_outs[8][5] ),
    .A2(\systolic_inst.A_outs[8][7] ),
    .A3(_05868_),
    .B1(_05867_),
    .X(_05892_));
 sky130_fd_sc_hd__nand3_2 _18770_ (.A(\systolic_inst.B_outs[8][5] ),
    .B(\systolic_inst.B_outs[8][6] ),
    .C(\systolic_inst.A_outs[8][7] ),
    .Y(_05893_));
 sky130_fd_sc_hd__o211a_2 _18771_ (.A1(_11259_),
    .A2(\systolic_inst.A_outs[8][7] ),
    .B1(_05839_),
    .C1(_05864_),
    .X(_05894_));
 sky130_fd_sc_hd__a21oi_2 _18772_ (.A1(_05892_),
    .A2(_05893_),
    .B1(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__or2_2 _18773_ (.A(_05806_),
    .B(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__nand2_2 _18774_ (.A(_05806_),
    .B(_05895_),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_2 _18775_ (.A(_05896_),
    .B(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__a21oi_2 _18776_ (.A1(_05871_),
    .A2(_05873_),
    .B1(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__and3_2 _18777_ (.A(_05871_),
    .B(_05873_),
    .C(_05898_),
    .X(_05900_));
 sky130_fd_sc_hd__nor2_2 _18778_ (.A(_05899_),
    .B(_05900_),
    .Y(_05901_));
 sky130_fd_sc_hd__xnor2_2 _18779_ (.A(_05835_),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__o21a_2 _18780_ (.A1(_05835_),
    .A2(_05878_),
    .B1(_05877_),
    .X(_05903_));
 sky130_fd_sc_hd__and2b_2 _18781_ (.A_N(_05903_),
    .B(_05902_),
    .X(_05904_));
 sky130_fd_sc_hd__and2b_2 _18782_ (.A_N(_05902_),
    .B(_05903_),
    .X(_05905_));
 sky130_fd_sc_hd__nor2_2 _18783_ (.A(_05904_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__xnor2_2 _18784_ (.A(_05834_),
    .B(_05906_),
    .Y(_05907_));
 sky130_fd_sc_hd__o21ba_2 _18785_ (.A1(_05834_),
    .A2(_05882_),
    .B1_N(_05881_),
    .X(_05908_));
 sky130_fd_sc_hd__nand2b_2 _18786_ (.A_N(_05908_),
    .B(_05907_),
    .Y(_05909_));
 sky130_fd_sc_hd__xnor2_2 _18787_ (.A(_05907_),
    .B(_05908_),
    .Y(_05910_));
 sky130_fd_sc_hd__o31a_2 _18788_ (.A1(_05856_),
    .A2(_05861_),
    .A3(_05885_),
    .B1(_05887_),
    .X(_05911_));
 sky130_fd_sc_hd__xor2_2 _18789_ (.A(_05910_),
    .B(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__mux2_1 _18790_ (.A0(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[14] ),
    .A1(_05912_),
    .S(\systolic_inst.ce_local ),
    .X(_01424_));
 sky130_fd_sc_hd__a31oi_2 _18791_ (.A1(_05694_),
    .A2(_05832_),
    .A3(_05906_),
    .B1(_05904_),
    .Y(_05913_));
 sky130_fd_sc_hd__a31o_2 _18792_ (.A1(_05833_),
    .A2(_05834_),
    .A3(_05901_),
    .B1(_05899_),
    .X(_05914_));
 sky130_fd_sc_hd__xnor2_2 _18793_ (.A(_05833_),
    .B(_05896_),
    .Y(_05915_));
 sky130_fd_sc_hd__xnor2_2 _18794_ (.A(_05914_),
    .B(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__xnor2_2 _18795_ (.A(_05913_),
    .B(_05916_),
    .Y(_05917_));
 sky130_fd_sc_hd__nand2_2 _18796_ (.A(_05909_),
    .B(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__a21oi_2 _18797_ (.A1(_05910_),
    .A2(_05911_),
    .B1(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__mux2_1 _18798_ (.A0(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .A1(_05919_),
    .S(\systolic_inst.ce_local ),
    .X(_01425_));
 sky130_fd_sc_hd__a21o_2 _18799_ (.A1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[8][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_05920_));
 sky130_fd_sc_hd__a21oi_2 _18800_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[8][0] ),
    .Y(_05921_));
 sky130_fd_sc_hd__a21oi_2 _18801_ (.A1(\systolic_inst.ce_local ),
    .A2(_05920_),
    .B1(_05921_),
    .Y(_01426_));
 sky130_fd_sc_hd__and2_2 _18802_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[8][1] ),
    .X(_05922_));
 sky130_fd_sc_hd__nand2_2 _18803_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[8][1] ),
    .Y(_05923_));
 sky130_fd_sc_hd__or2_2 _18804_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[8][1] ),
    .X(_05924_));
 sky130_fd_sc_hd__and4_2 _18805_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[8][0] ),
    .C(_05923_),
    .D(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__inv_2 _18806_ (.A(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__a22o_2 _18807_ (.A1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[8][0] ),
    .B1(_05923_),
    .B2(_05924_),
    .X(_05927_));
 sky130_fd_sc_hd__a32o_2 _18808_ (.A1(_11712_),
    .A2(_05926_),
    .A3(_05927_),
    .B1(\systolic_inst.acc_wires[8][1] ),
    .B2(_11258_),
    .X(_01427_));
 sky130_fd_sc_hd__and2_2 _18809_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[8][2] ),
    .X(_05928_));
 sky130_fd_sc_hd__nand2_2 _18810_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[8][2] ),
    .Y(_05929_));
 sky130_fd_sc_hd__or2_2 _18811_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[8][2] ),
    .X(_05930_));
 sky130_fd_sc_hd__a211o_2 _18812_ (.A1(_05929_),
    .A2(_05930_),
    .B1(_05922_),
    .C1(_05925_),
    .X(_05931_));
 sky130_fd_sc_hd__o211a_2 _18813_ (.A1(_05922_),
    .A2(_05925_),
    .B1(_05929_),
    .C1(_05930_),
    .X(_05932_));
 sky130_fd_sc_hd__inv_2 _18814_ (.A(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__a32o_2 _18815_ (.A1(_11712_),
    .A2(_05931_),
    .A3(_05933_),
    .B1(\systolic_inst.acc_wires[8][2] ),
    .B2(_11258_),
    .X(_01428_));
 sky130_fd_sc_hd__and2_2 _18816_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[8][3] ),
    .X(_05934_));
 sky130_fd_sc_hd__nand2_2 _18817_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[8][3] ),
    .Y(_05935_));
 sky130_fd_sc_hd__or2_2 _18818_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[8][3] ),
    .X(_05936_));
 sky130_fd_sc_hd__a211o_2 _18819_ (.A1(_05935_),
    .A2(_05936_),
    .B1(_05928_),
    .C1(_05932_),
    .X(_05937_));
 sky130_fd_sc_hd__o211a_2 _18820_ (.A1(_05928_),
    .A2(_05932_),
    .B1(_05935_),
    .C1(_05936_),
    .X(_05938_));
 sky130_fd_sc_hd__inv_2 _18821_ (.A(_05938_),
    .Y(_05939_));
 sky130_fd_sc_hd__a32o_2 _18822_ (.A1(_11712_),
    .A2(_05937_),
    .A3(_05939_),
    .B1(\systolic_inst.acc_wires[8][3] ),
    .B2(_11258_),
    .X(_01429_));
 sky130_fd_sc_hd__and2_2 _18823_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[8][4] ),
    .X(_05940_));
 sky130_fd_sc_hd__nand2_2 _18824_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[8][4] ),
    .Y(_05941_));
 sky130_fd_sc_hd__or2_2 _18825_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[8][4] ),
    .X(_05942_));
 sky130_fd_sc_hd__a211o_2 _18826_ (.A1(_05941_),
    .A2(_05942_),
    .B1(_05934_),
    .C1(_05938_),
    .X(_05943_));
 sky130_fd_sc_hd__o211a_2 _18827_ (.A1(_05934_),
    .A2(_05938_),
    .B1(_05941_),
    .C1(_05942_),
    .X(_05944_));
 sky130_fd_sc_hd__inv_2 _18828_ (.A(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__a32o_2 _18829_ (.A1(_11712_),
    .A2(_05943_),
    .A3(_05945_),
    .B1(\systolic_inst.acc_wires[8][4] ),
    .B2(_11258_),
    .X(_01430_));
 sky130_fd_sc_hd__and2_2 _18830_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[8][5] ),
    .X(_05946_));
 sky130_fd_sc_hd__nand2_2 _18831_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[8][5] ),
    .Y(_05947_));
 sky130_fd_sc_hd__or2_2 _18832_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[8][5] ),
    .X(_05948_));
 sky130_fd_sc_hd__a211o_2 _18833_ (.A1(_05947_),
    .A2(_05948_),
    .B1(_05940_),
    .C1(_05944_),
    .X(_05949_));
 sky130_fd_sc_hd__o211a_2 _18834_ (.A1(_05940_),
    .A2(_05944_),
    .B1(_05947_),
    .C1(_05948_),
    .X(_05950_));
 sky130_fd_sc_hd__inv_2 _18835_ (.A(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__a32o_2 _18836_ (.A1(_11712_),
    .A2(_05949_),
    .A3(_05951_),
    .B1(\systolic_inst.acc_wires[8][5] ),
    .B2(_11258_),
    .X(_01431_));
 sky130_fd_sc_hd__nand2_2 _18837_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[8][6] ),
    .Y(_05952_));
 sky130_fd_sc_hd__or2_2 _18838_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[8][6] ),
    .X(_05953_));
 sky130_fd_sc_hd__o211ai_2 _18839_ (.A1(_05946_),
    .A2(_05950_),
    .B1(_05952_),
    .C1(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__a211o_2 _18840_ (.A1(_05952_),
    .A2(_05953_),
    .B1(_05946_),
    .C1(_05950_),
    .X(_05955_));
 sky130_fd_sc_hd__a32o_2 _18841_ (.A1(_11712_),
    .A2(_05954_),
    .A3(_05955_),
    .B1(\systolic_inst.acc_wires[8][6] ),
    .B2(_11258_),
    .X(_01432_));
 sky130_fd_sc_hd__nand2_2 _18842_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[8][7] ),
    .Y(_05956_));
 sky130_fd_sc_hd__or2_2 _18843_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[8][7] ),
    .X(_05957_));
 sky130_fd_sc_hd__nand2_2 _18844_ (.A(_05956_),
    .B(_05957_),
    .Y(_05958_));
 sky130_fd_sc_hd__nand3_2 _18845_ (.A(_05952_),
    .B(_05954_),
    .C(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__a21o_2 _18846_ (.A1(_05952_),
    .A2(_05954_),
    .B1(_05958_),
    .X(_05960_));
 sky130_fd_sc_hd__a32o_2 _18847_ (.A1(_11712_),
    .A2(_05959_),
    .A3(_05960_),
    .B1(\systolic_inst.acc_wires[8][7] ),
    .B2(_11258_),
    .X(_01433_));
 sky130_fd_sc_hd__or2_2 _18848_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[8][8] ),
    .X(_05961_));
 sky130_fd_sc_hd__nand2_2 _18849_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[8][8] ),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2_2 _18850_ (.A(_05961_),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__a21o_2 _18851_ (.A1(_05956_),
    .A2(_05960_),
    .B1(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__nand3_2 _18852_ (.A(_05956_),
    .B(_05960_),
    .C(_05963_),
    .Y(_05965_));
 sky130_fd_sc_hd__a32o_2 _18853_ (.A1(_11712_),
    .A2(_05964_),
    .A3(_05965_),
    .B1(\systolic_inst.acc_wires[8][8] ),
    .B2(_11258_),
    .X(_01434_));
 sky130_fd_sc_hd__nor2_2 _18854_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[8][9] ),
    .Y(_05966_));
 sky130_fd_sc_hd__nand2_2 _18855_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[8][9] ),
    .Y(_05967_));
 sky130_fd_sc_hd__and2b_2 _18856_ (.A_N(_05966_),
    .B(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__nand2_2 _18857_ (.A(_05962_),
    .B(_05964_),
    .Y(_05969_));
 sky130_fd_sc_hd__or2_2 _18858_ (.A(_05968_),
    .B(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__a21bo_2 _18859_ (.A1(_05962_),
    .A2(_05964_),
    .B1_N(_05968_),
    .X(_05971_));
 sky130_fd_sc_hd__a32o_2 _18860_ (.A1(_11712_),
    .A2(_05970_),
    .A3(_05971_),
    .B1(\systolic_inst.acc_wires[8][9] ),
    .B2(_11258_),
    .X(_01435_));
 sky130_fd_sc_hd__or2_2 _18861_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[8][10] ),
    .X(_05972_));
 sky130_fd_sc_hd__nand2_2 _18862_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[8][10] ),
    .Y(_05973_));
 sky130_fd_sc_hd__nand2_2 _18863_ (.A(_05972_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__nand3_2 _18864_ (.A(_05967_),
    .B(_05971_),
    .C(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__a21o_2 _18865_ (.A1(_05967_),
    .A2(_05971_),
    .B1(_05974_),
    .X(_05976_));
 sky130_fd_sc_hd__a32o_2 _18866_ (.A1(_11712_),
    .A2(_05975_),
    .A3(_05976_),
    .B1(\systolic_inst.acc_wires[8][10] ),
    .B2(_11258_),
    .X(_01436_));
 sky130_fd_sc_hd__or2_2 _18867_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[8][11] ),
    .X(_05977_));
 sky130_fd_sc_hd__nand2_2 _18868_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[8][11] ),
    .Y(_05978_));
 sky130_fd_sc_hd__nand2_2 _18869_ (.A(_05977_),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__a21oi_2 _18870_ (.A1(_05973_),
    .A2(_05976_),
    .B1(_05979_),
    .Y(_05980_));
 sky130_fd_sc_hd__a31o_2 _18871_ (.A1(_05973_),
    .A2(_05976_),
    .A3(_05979_),
    .B1(_11713_),
    .X(_05981_));
 sky130_fd_sc_hd__a2bb2o_2 _18872_ (.A1_N(_05981_),
    .A2_N(_05980_),
    .B1(\systolic_inst.acc_wires[8][11] ),
    .B2(_11258_),
    .X(_01437_));
 sky130_fd_sc_hd__nor2_2 _18873_ (.A(_05974_),
    .B(_05979_),
    .Y(_05982_));
 sky130_fd_sc_hd__nand2_2 _18874_ (.A(_05968_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__a211o_2 _18875_ (.A1(_05956_),
    .A2(_05960_),
    .B1(_05963_),
    .C1(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__o21ai_2 _18876_ (.A1(_05962_),
    .A2(_05966_),
    .B1(_05967_),
    .Y(_05985_));
 sky130_fd_sc_hd__and3_2 _18877_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[8][10] ),
    .C(_05977_),
    .X(_05986_));
 sky130_fd_sc_hd__a221oi_2 _18878_ (.A1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[11] ),
    .A2(\systolic_inst.acc_wires[8][11] ),
    .B1(_05982_),
    .B2(_05985_),
    .C1(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__or2_2 _18879_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[8][12] ),
    .X(_05988_));
 sky130_fd_sc_hd__nand2_2 _18880_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[8][12] ),
    .Y(_05989_));
 sky130_fd_sc_hd__nand2_2 _18881_ (.A(_05988_),
    .B(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__a21oi_2 _18882_ (.A1(_05984_),
    .A2(_05987_),
    .B1(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__a31o_2 _18883_ (.A1(_05984_),
    .A2(_05987_),
    .A3(_05990_),
    .B1(_11713_),
    .X(_05992_));
 sky130_fd_sc_hd__a2bb2o_2 _18884_ (.A1_N(_05992_),
    .A2_N(_05991_),
    .B1(\systolic_inst.acc_wires[8][12] ),
    .B2(_11258_),
    .X(_01438_));
 sky130_fd_sc_hd__or2_2 _18885_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[8][13] ),
    .X(_05993_));
 sky130_fd_sc_hd__nand2_2 _18886_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[8][13] ),
    .Y(_05994_));
 sky130_fd_sc_hd__nand2_2 _18887_ (.A(_05993_),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand2_2 _18888_ (.A(_05989_),
    .B(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__a211o_2 _18889_ (.A1(_05984_),
    .A2(_05987_),
    .B1(_05990_),
    .C1(_05995_),
    .X(_05997_));
 sky130_fd_sc_hd__or2_2 _18890_ (.A(_05989_),
    .B(_05995_),
    .X(_05998_));
 sky130_fd_sc_hd__o211a_2 _18891_ (.A1(_05991_),
    .A2(_05996_),
    .B1(_05997_),
    .C1(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__a22o_2 _18892_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[8][13] ),
    .B1(_11712_),
    .B2(_05999_),
    .X(_01439_));
 sky130_fd_sc_hd__or2_2 _18893_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[8][14] ),
    .X(_06000_));
 sky130_fd_sc_hd__nand2_2 _18894_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[8][14] ),
    .Y(_06001_));
 sky130_fd_sc_hd__and2_2 _18895_ (.A(_06000_),
    .B(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__and2_2 _18896_ (.A(_05994_),
    .B(_05998_),
    .X(_06003_));
 sky130_fd_sc_hd__nand2_2 _18897_ (.A(_05997_),
    .B(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__nand2_2 _18898_ (.A(_06002_),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__or2_2 _18899_ (.A(_06002_),
    .B(_06004_),
    .X(_06006_));
 sky130_fd_sc_hd__a32o_2 _18900_ (.A1(_11712_),
    .A2(_06005_),
    .A3(_06006_),
    .B1(\systolic_inst.acc_wires[8][14] ),
    .B2(_11258_),
    .X(_01440_));
 sky130_fd_sc_hd__nor2_2 _18901_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][15] ),
    .Y(_06007_));
 sky130_fd_sc_hd__and2_2 _18902_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][15] ),
    .X(_06008_));
 sky130_fd_sc_hd__a211o_2 _18903_ (.A1(_06001_),
    .A2(_06005_),
    .B1(_06007_),
    .C1(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__o211ai_2 _18904_ (.A1(_06007_),
    .A2(_06008_),
    .B1(_06001_),
    .C1(_06005_),
    .Y(_06010_));
 sky130_fd_sc_hd__a32o_2 _18905_ (.A1(_11712_),
    .A2(_06009_),
    .A3(_06010_),
    .B1(\systolic_inst.acc_wires[8][15] ),
    .B2(_11258_),
    .X(_01441_));
 sky130_fd_sc_hd__or3b_2 _18906_ (.A(_06007_),
    .B(_06008_),
    .C_N(_06002_),
    .X(_06011_));
 sky130_fd_sc_hd__a21o_2 _18907_ (.A1(_05997_),
    .A2(_06003_),
    .B1(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__o21ba_2 _18908_ (.A1(_06001_),
    .A2(_06007_),
    .B1_N(_06008_),
    .X(_06013_));
 sky130_fd_sc_hd__and2_2 _18909_ (.A(_06012_),
    .B(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__or2_2 _18910_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][16] ),
    .X(_06015_));
 sky130_fd_sc_hd__nand2_2 _18911_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][16] ),
    .Y(_06016_));
 sky130_fd_sc_hd__nand2_2 _18912_ (.A(_06015_),
    .B(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand2_2 _18913_ (.A(_06014_),
    .B(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__nor2_2 _18914_ (.A(_06014_),
    .B(_06017_),
    .Y(_06019_));
 sky130_fd_sc_hd__or2_2 _18915_ (.A(_06014_),
    .B(_06017_),
    .X(_06020_));
 sky130_fd_sc_hd__a32o_2 _18916_ (.A1(_11712_),
    .A2(_06018_),
    .A3(_06020_),
    .B1(\systolic_inst.acc_wires[8][16] ),
    .B2(_11258_),
    .X(_01442_));
 sky130_fd_sc_hd__xor2_2 _18917_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][17] ),
    .X(_06021_));
 sky130_fd_sc_hd__inv_2 _18918_ (.A(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__o21a_2 _18919_ (.A1(_06014_),
    .A2(_06017_),
    .B1(_06016_),
    .X(_06023_));
 sky130_fd_sc_hd__xnor2_2 _18920_ (.A(_06021_),
    .B(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__a22o_2 _18921_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[8][17] ),
    .B1(_11712_),
    .B2(_06024_),
    .X(_01443_));
 sky130_fd_sc_hd__or2_2 _18922_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][18] ),
    .X(_06025_));
 sky130_fd_sc_hd__nand2_2 _18923_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][18] ),
    .Y(_06026_));
 sky130_fd_sc_hd__nand2_2 _18924_ (.A(_06025_),
    .B(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__o21ai_2 _18925_ (.A1(\systolic_inst.acc_wires[8][16] ),
    .A2(\systolic_inst.acc_wires[8][17] ),
    .B1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .Y(_06028_));
 sky130_fd_sc_hd__nand2_2 _18926_ (.A(_06019_),
    .B(_06021_),
    .Y(_06029_));
 sky130_fd_sc_hd__a21o_2 _18927_ (.A1(_06028_),
    .A2(_06029_),
    .B1(_06027_),
    .X(_06030_));
 sky130_fd_sc_hd__nand3_2 _18928_ (.A(_06027_),
    .B(_06028_),
    .C(_06029_),
    .Y(_06031_));
 sky130_fd_sc_hd__a32o_2 _18929_ (.A1(_11712_),
    .A2(_06030_),
    .A3(_06031_),
    .B1(\systolic_inst.acc_wires[8][18] ),
    .B2(_11258_),
    .X(_01444_));
 sky130_fd_sc_hd__xnor2_2 _18930_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][19] ),
    .Y(_06032_));
 sky130_fd_sc_hd__a21oi_2 _18931_ (.A1(_06026_),
    .A2(_06030_),
    .B1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__a31o_2 _18932_ (.A1(_06026_),
    .A2(_06030_),
    .A3(_06032_),
    .B1(_11713_),
    .X(_06034_));
 sky130_fd_sc_hd__a2bb2o_2 _18933_ (.A1_N(_06034_),
    .A2_N(_06033_),
    .B1(\systolic_inst.acc_wires[8][19] ),
    .B2(_11258_),
    .X(_01445_));
 sky130_fd_sc_hd__or2_2 _18934_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][20] ),
    .X(_06035_));
 sky130_fd_sc_hd__nand2_2 _18935_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][20] ),
    .Y(_06036_));
 sky130_fd_sc_hd__and2_2 _18936_ (.A(_06035_),
    .B(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__or4_2 _18937_ (.A(_06017_),
    .B(_06022_),
    .C(_06027_),
    .D(_06032_),
    .X(_06038_));
 sky130_fd_sc_hd__nor2_2 _18938_ (.A(_06014_),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__o41a_2 _18939_ (.A1(\systolic_inst.acc_wires[8][16] ),
    .A2(\systolic_inst.acc_wires[8][17] ),
    .A3(\systolic_inst.acc_wires[8][18] ),
    .A4(\systolic_inst.acc_wires[8][19] ),
    .B1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .X(_06040_));
 sky130_fd_sc_hd__or3_2 _18940_ (.A(_06037_),
    .B(_06039_),
    .C(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__o21ai_2 _18941_ (.A1(_06039_),
    .A2(_06040_),
    .B1(_06037_),
    .Y(_06042_));
 sky130_fd_sc_hd__a32o_2 _18942_ (.A1(_11712_),
    .A2(_06041_),
    .A3(_06042_),
    .B1(\systolic_inst.acc_wires[8][20] ),
    .B2(_11258_),
    .X(_01446_));
 sky130_fd_sc_hd__xnor2_2 _18943_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][21] ),
    .Y(_06043_));
 sky130_fd_sc_hd__inv_2 _18944_ (.A(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__a21oi_2 _18945_ (.A1(_06036_),
    .A2(_06042_),
    .B1(_06043_),
    .Y(_06045_));
 sky130_fd_sc_hd__a31o_2 _18946_ (.A1(_06036_),
    .A2(_06042_),
    .A3(_06043_),
    .B1(_11713_),
    .X(_06046_));
 sky130_fd_sc_hd__a2bb2o_2 _18947_ (.A1_N(_06046_),
    .A2_N(_06045_),
    .B1(\systolic_inst.acc_wires[8][21] ),
    .B2(_11258_),
    .X(_01447_));
 sky130_fd_sc_hd__or2_2 _18948_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][22] ),
    .X(_06047_));
 sky130_fd_sc_hd__nand2_2 _18949_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][22] ),
    .Y(_06048_));
 sky130_fd_sc_hd__and2_2 _18950_ (.A(_06047_),
    .B(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__o21a_2 _18951_ (.A1(\systolic_inst.acc_wires[8][20] ),
    .A2(\systolic_inst.acc_wires[8][21] ),
    .B1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .X(_06050_));
 sky130_fd_sc_hd__nor2_2 _18952_ (.A(_06042_),
    .B(_06043_),
    .Y(_06051_));
 sky130_fd_sc_hd__o21ai_2 _18953_ (.A1(_06050_),
    .A2(_06051_),
    .B1(_06049_),
    .Y(_06052_));
 sky130_fd_sc_hd__or3_2 _18954_ (.A(_06049_),
    .B(_06050_),
    .C(_06051_),
    .X(_06053_));
 sky130_fd_sc_hd__a32o_2 _18955_ (.A1(_11712_),
    .A2(_06052_),
    .A3(_06053_),
    .B1(\systolic_inst.acc_wires[8][22] ),
    .B2(_11258_),
    .X(_01448_));
 sky130_fd_sc_hd__xor2_2 _18956_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][23] ),
    .X(_06054_));
 sky130_fd_sc_hd__inv_2 _18957_ (.A(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__nand3_2 _18958_ (.A(_06048_),
    .B(_06052_),
    .C(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__a21o_2 _18959_ (.A1(_06048_),
    .A2(_06052_),
    .B1(_06055_),
    .X(_06057_));
 sky130_fd_sc_hd__a32o_2 _18960_ (.A1(_11712_),
    .A2(_06056_),
    .A3(_06057_),
    .B1(\systolic_inst.acc_wires[8][23] ),
    .B2(_11258_),
    .X(_01449_));
 sky130_fd_sc_hd__nand4_2 _18961_ (.A(_06037_),
    .B(_06044_),
    .C(_06049_),
    .D(_06054_),
    .Y(_06058_));
 sky130_fd_sc_hd__a211o_2 _18962_ (.A1(_06012_),
    .A2(_06013_),
    .B1(_06038_),
    .C1(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__o41a_2 _18963_ (.A1(\systolic_inst.acc_wires[8][20] ),
    .A2(\systolic_inst.acc_wires[8][21] ),
    .A3(\systolic_inst.acc_wires[8][22] ),
    .A4(\systolic_inst.acc_wires[8][23] ),
    .B1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .X(_06060_));
 sky130_fd_sc_hd__nor2_2 _18964_ (.A(_06040_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__nor2_2 _18965_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][24] ),
    .Y(_06062_));
 sky130_fd_sc_hd__and2_2 _18966_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][24] ),
    .X(_06063_));
 sky130_fd_sc_hd__or2_2 _18967_ (.A(_06062_),
    .B(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__a21oi_2 _18968_ (.A1(_06059_),
    .A2(_06061_),
    .B1(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__a31o_2 _18969_ (.A1(_06059_),
    .A2(_06061_),
    .A3(_06064_),
    .B1(_11713_),
    .X(_06066_));
 sky130_fd_sc_hd__a2bb2o_2 _18970_ (.A1_N(_06066_),
    .A2_N(_06065_),
    .B1(\systolic_inst.acc_wires[8][24] ),
    .B2(_11258_),
    .X(_01450_));
 sky130_fd_sc_hd__xor2_2 _18971_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][25] ),
    .X(_06067_));
 sky130_fd_sc_hd__or3_2 _18972_ (.A(_06063_),
    .B(_06065_),
    .C(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__o21ai_2 _18973_ (.A1(_06063_),
    .A2(_06065_),
    .B1(_06067_),
    .Y(_06069_));
 sky130_fd_sc_hd__a32o_2 _18974_ (.A1(_11712_),
    .A2(_06068_),
    .A3(_06069_),
    .B1(\systolic_inst.acc_wires[8][25] ),
    .B2(_11258_),
    .X(_01451_));
 sky130_fd_sc_hd__or2_2 _18975_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][26] ),
    .X(_06070_));
 sky130_fd_sc_hd__nand2_2 _18976_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][26] ),
    .Y(_06071_));
 sky130_fd_sc_hd__nand2_2 _18977_ (.A(_06070_),
    .B(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__o21a_2 _18978_ (.A1(\systolic_inst.acc_wires[8][24] ),
    .A2(\systolic_inst.acc_wires[8][25] ),
    .B1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .X(_06073_));
 sky130_fd_sc_hd__a21o_2 _18979_ (.A1(_06065_),
    .A2(_06067_),
    .B1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__xnor2_2 _18980_ (.A(_06072_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__a22o_2 _18981_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[8][26] ),
    .B1(_11712_),
    .B2(_06075_),
    .X(_01452_));
 sky130_fd_sc_hd__xnor2_2 _18982_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][27] ),
    .Y(_06076_));
 sky130_fd_sc_hd__a21bo_2 _18983_ (.A1(_06070_),
    .A2(_06074_),
    .B1_N(_06071_),
    .X(_06077_));
 sky130_fd_sc_hd__xnor2_2 _18984_ (.A(_06076_),
    .B(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__a22o_2 _18985_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[8][27] ),
    .B1(_11712_),
    .B2(_06078_),
    .X(_01453_));
 sky130_fd_sc_hd__nor2_2 _18986_ (.A(_06072_),
    .B(_06076_),
    .Y(_06079_));
 sky130_fd_sc_hd__o21a_2 _18987_ (.A1(\systolic_inst.acc_wires[8][26] ),
    .A2(\systolic_inst.acc_wires[8][27] ),
    .B1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .X(_06080_));
 sky130_fd_sc_hd__a311oi_2 _18988_ (.A1(_06065_),
    .A2(_06067_),
    .A3(_06079_),
    .B1(_06080_),
    .C1(_06073_),
    .Y(_06081_));
 sky130_fd_sc_hd__or2_2 _18989_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][28] ),
    .X(_06082_));
 sky130_fd_sc_hd__nand2_2 _18990_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][28] ),
    .Y(_06083_));
 sky130_fd_sc_hd__nand2_2 _18991_ (.A(_06082_),
    .B(_06083_),
    .Y(_06084_));
 sky130_fd_sc_hd__xor2_2 _18992_ (.A(_06081_),
    .B(_06084_),
    .X(_06085_));
 sky130_fd_sc_hd__a22o_2 _18993_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[8][28] ),
    .B1(_11712_),
    .B2(_06085_),
    .X(_01454_));
 sky130_fd_sc_hd__xor2_2 _18994_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][29] ),
    .X(_06086_));
 sky130_fd_sc_hd__inv_2 _18995_ (.A(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__o21a_2 _18996_ (.A1(_06081_),
    .A2(_06084_),
    .B1(_06083_),
    .X(_06088_));
 sky130_fd_sc_hd__xnor2_2 _18997_ (.A(_06086_),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__a22o_2 _18998_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[8][29] ),
    .B1(_11712_),
    .B2(_06089_),
    .X(_01455_));
 sky130_fd_sc_hd__o21ai_2 _18999_ (.A1(\systolic_inst.acc_wires[8][28] ),
    .A2(\systolic_inst.acc_wires[8][29] ),
    .B1(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .Y(_06090_));
 sky130_fd_sc_hd__o31a_2 _19000_ (.A1(_06081_),
    .A2(_06084_),
    .A3(_06087_),
    .B1(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__nand2_2 _19001_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][30] ),
    .Y(_06092_));
 sky130_fd_sc_hd__or2_2 _19002_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][30] ),
    .X(_06093_));
 sky130_fd_sc_hd__nand2_2 _19003_ (.A(_06092_),
    .B(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__nand2_2 _19004_ (.A(_06091_),
    .B(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__or2_2 _19005_ (.A(_06091_),
    .B(_06094_),
    .X(_06096_));
 sky130_fd_sc_hd__a32o_2 _19006_ (.A1(_11712_),
    .A2(_06095_),
    .A3(_06096_),
    .B1(\systolic_inst.acc_wires[8][30] ),
    .B2(_11258_),
    .X(_01456_));
 sky130_fd_sc_hd__xnor2_2 _19007_ (.A(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[8][31] ),
    .Y(_06097_));
 sky130_fd_sc_hd__a21oi_2 _19008_ (.A1(_06092_),
    .A2(_06096_),
    .B1(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__a31o_2 _19009_ (.A1(_06092_),
    .A2(_06096_),
    .A3(_06097_),
    .B1(_11713_),
    .X(_06099_));
 sky130_fd_sc_hd__a2bb2o_2 _19010_ (.A1_N(_06099_),
    .A2_N(_06098_),
    .B1(\systolic_inst.acc_wires[8][31] ),
    .B2(_11258_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _19011_ (.A0(\systolic_inst.A_outs[7][0] ),
    .A1(\systolic_inst.A_outs[6][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _19012_ (.A0(\systolic_inst.A_outs[7][1] ),
    .A1(\systolic_inst.A_outs[6][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _19013_ (.A0(\systolic_inst.A_outs[7][2] ),
    .A1(\systolic_inst.A_outs[6][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _19014_ (.A0(\systolic_inst.A_outs[7][3] ),
    .A1(\systolic_inst.A_outs[6][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _19015_ (.A0(\systolic_inst.A_outs[7][4] ),
    .A1(\systolic_inst.A_outs[6][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _19016_ (.A0(\systolic_inst.A_outs[7][5] ),
    .A1(\systolic_inst.A_outs[6][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _19017_ (.A0(\systolic_inst.A_outs[7][6] ),
    .A1(\systolic_inst.A_outs[6][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _19018_ (.A0(\systolic_inst.A_outs[7][7] ),
    .A1(\systolic_inst.A_outs[6][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _19019_ (.A0(\systolic_inst.B_outs[6][0] ),
    .A1(\systolic_inst.B_outs[2][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _19020_ (.A0(\systolic_inst.B_outs[6][1] ),
    .A1(\systolic_inst.B_outs[2][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _19021_ (.A0(\systolic_inst.B_outs[6][2] ),
    .A1(\systolic_inst.B_outs[2][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _19022_ (.A0(\systolic_inst.B_outs[6][3] ),
    .A1(\systolic_inst.B_outs[2][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _19023_ (.A0(\systolic_inst.B_outs[6][4] ),
    .A1(\systolic_inst.B_outs[2][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _19024_ (.A0(\systolic_inst.B_outs[6][5] ),
    .A1(\systolic_inst.B_outs[2][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _19025_ (.A0(\systolic_inst.B_outs[6][6] ),
    .A1(\systolic_inst.B_outs[2][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _19026_ (.A0(\systolic_inst.B_outs[6][7] ),
    .A1(\systolic_inst.B_outs[2][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01473_));
 sky130_fd_sc_hd__and3_2 _19027_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[7][0] ),
    .C(\systolic_inst.A_outs[7][0] ),
    .X(_06100_));
 sky130_fd_sc_hd__a21o_2 _19028_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[0] ),
    .B1(_06100_),
    .X(_01474_));
 sky130_fd_sc_hd__and4_2 _19029_ (.A(\systolic_inst.B_outs[7][0] ),
    .B(\systolic_inst.A_outs[7][0] ),
    .C(\systolic_inst.B_outs[7][1] ),
    .D(\systolic_inst.A_outs[7][1] ),
    .X(_06101_));
 sky130_fd_sc_hd__a22o_2 _19030_ (.A1(\systolic_inst.A_outs[7][0] ),
    .A2(\systolic_inst.B_outs[7][1] ),
    .B1(\systolic_inst.A_outs[7][1] ),
    .B2(\systolic_inst.B_outs[7][0] ),
    .X(_06102_));
 sky130_fd_sc_hd__nand2_2 _19031_ (.A(\systolic_inst.ce_local ),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__a2bb2o_2 _19032_ (.A1_N(_06103_),
    .A2_N(_06101_),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01475_));
 sky130_fd_sc_hd__and2_2 _19033_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[2] ),
    .X(_06104_));
 sky130_fd_sc_hd__a22oi_2 _19034_ (.A1(\systolic_inst.B_outs[7][1] ),
    .A2(\systolic_inst.A_outs[7][1] ),
    .B1(\systolic_inst.A_outs[7][2] ),
    .B2(\systolic_inst.B_outs[7][0] ),
    .Y(_06105_));
 sky130_fd_sc_hd__and4_2 _19035_ (.A(\systolic_inst.B_outs[7][0] ),
    .B(\systolic_inst.B_outs[7][1] ),
    .C(\systolic_inst.A_outs[7][1] ),
    .D(\systolic_inst.A_outs[7][2] ),
    .X(_06106_));
 sky130_fd_sc_hd__or2_2 _19036_ (.A(_06105_),
    .B(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__or3b_2 _19037_ (.A(_06105_),
    .B(_06106_),
    .C_N(_06101_),
    .X(_06108_));
 sky130_fd_sc_hd__xnor2_2 _19038_ (.A(_06101_),
    .B(_06107_),
    .Y(_06109_));
 sky130_fd_sc_hd__nand3_2 _19039_ (.A(\systolic_inst.A_outs[7][0] ),
    .B(\systolic_inst.B_outs[7][2] ),
    .C(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__a21o_2 _19040_ (.A1(\systolic_inst.A_outs[7][0] ),
    .A2(\systolic_inst.B_outs[7][2] ),
    .B1(_06109_),
    .X(_06111_));
 sky130_fd_sc_hd__a31o_2 _19041_ (.A1(\systolic_inst.ce_local ),
    .A2(_06110_),
    .A3(_06111_),
    .B1(_06104_),
    .X(_01476_));
 sky130_fd_sc_hd__a22oi_2 _19042_ (.A1(\systolic_inst.A_outs[7][1] ),
    .A2(\systolic_inst.B_outs[7][2] ),
    .B1(\systolic_inst.B_outs[7][3] ),
    .B2(\systolic_inst.A_outs[7][0] ),
    .Y(_06112_));
 sky130_fd_sc_hd__and4_2 _19043_ (.A(\systolic_inst.A_outs[7][0] ),
    .B(\systolic_inst.A_outs[7][1] ),
    .C(\systolic_inst.B_outs[7][2] ),
    .D(\systolic_inst.B_outs[7][3] ),
    .X(_06113_));
 sky130_fd_sc_hd__nor2_2 _19044_ (.A(_06112_),
    .B(_06113_),
    .Y(_06114_));
 sky130_fd_sc_hd__nand4_2 _19045_ (.A(\systolic_inst.B_outs[7][0] ),
    .B(\systolic_inst.B_outs[7][1] ),
    .C(\systolic_inst.A_outs[7][2] ),
    .D(\systolic_inst.A_outs[7][3] ),
    .Y(_06115_));
 sky130_fd_sc_hd__a22o_2 _19046_ (.A1(\systolic_inst.B_outs[7][1] ),
    .A2(\systolic_inst.A_outs[7][2] ),
    .B1(\systolic_inst.A_outs[7][3] ),
    .B2(\systolic_inst.B_outs[7][0] ),
    .X(_06116_));
 sky130_fd_sc_hd__nand3_2 _19047_ (.A(_06106_),
    .B(_06115_),
    .C(_06116_),
    .Y(_06117_));
 sky130_fd_sc_hd__a21o_2 _19048_ (.A1(_06115_),
    .A2(_06116_),
    .B1(_06106_),
    .X(_06118_));
 sky130_fd_sc_hd__and2_2 _19049_ (.A(_06117_),
    .B(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__nand2_2 _19050_ (.A(_06114_),
    .B(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__xnor2_2 _19051_ (.A(_06114_),
    .B(_06119_),
    .Y(_06121_));
 sky130_fd_sc_hd__and3_2 _19052_ (.A(_06108_),
    .B(_06110_),
    .C(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__a21oi_2 _19053_ (.A1(_06108_),
    .A2(_06110_),
    .B1(_06121_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_2 _19054_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[3] ),
    .Y(_06124_));
 sky130_fd_sc_hd__o31ai_2 _19055_ (.A1(_11258_),
    .A2(_06122_),
    .A3(_06123_),
    .B1(_06124_),
    .Y(_01477_));
 sky130_fd_sc_hd__and2_2 _19056_ (.A(\systolic_inst.B_outs[7][2] ),
    .B(\systolic_inst.A_outs[7][2] ),
    .X(_06125_));
 sky130_fd_sc_hd__nand4_2 _19057_ (.A(\systolic_inst.A_outs[7][0] ),
    .B(\systolic_inst.A_outs[7][1] ),
    .C(\systolic_inst.B_outs[7][3] ),
    .D(\systolic_inst.B_outs[7][4] ),
    .Y(_06126_));
 sky130_fd_sc_hd__a22o_2 _19058_ (.A1(\systolic_inst.A_outs[7][1] ),
    .A2(\systolic_inst.B_outs[7][3] ),
    .B1(\systolic_inst.B_outs[7][4] ),
    .B2(\systolic_inst.A_outs[7][0] ),
    .X(_06127_));
 sky130_fd_sc_hd__nand2_2 _19059_ (.A(_06126_),
    .B(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__xnor2_2 _19060_ (.A(_06125_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__a22o_2 _19061_ (.A1(\systolic_inst.B_outs[7][1] ),
    .A2(\systolic_inst.A_outs[7][3] ),
    .B1(\systolic_inst.A_outs[7][4] ),
    .B2(\systolic_inst.B_outs[7][0] ),
    .X(_06130_));
 sky130_fd_sc_hd__and3_2 _19062_ (.A(\systolic_inst.B_outs[7][0] ),
    .B(\systolic_inst.B_outs[7][1] ),
    .C(\systolic_inst.A_outs[7][3] ),
    .X(_06131_));
 sky130_fd_sc_hd__nand2_2 _19063_ (.A(\systolic_inst.A_outs[7][4] ),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__and3_2 _19064_ (.A(_06113_),
    .B(_06130_),
    .C(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__a21oi_2 _19065_ (.A1(_06130_),
    .A2(_06132_),
    .B1(_06113_),
    .Y(_06134_));
 sky130_fd_sc_hd__o21ai_2 _19066_ (.A1(_06133_),
    .A2(_06134_),
    .B1(_06115_),
    .Y(_06135_));
 sky130_fd_sc_hd__or3_2 _19067_ (.A(_06115_),
    .B(_06133_),
    .C(_06134_),
    .X(_06136_));
 sky130_fd_sc_hd__and3_2 _19068_ (.A(_06129_),
    .B(_06135_),
    .C(_06136_),
    .X(_06137_));
 sky130_fd_sc_hd__a21oi_2 _19069_ (.A1(_06135_),
    .A2(_06136_),
    .B1(_06129_),
    .Y(_06138_));
 sky130_fd_sc_hd__a211o_2 _19070_ (.A1(_06117_),
    .A2(_06120_),
    .B1(_06137_),
    .C1(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__o211ai_2 _19071_ (.A1(_06137_),
    .A2(_06138_),
    .B1(_06117_),
    .C1(_06120_),
    .Y(_06140_));
 sky130_fd_sc_hd__a21oi_2 _19072_ (.A1(_06139_),
    .A2(_06140_),
    .B1(_06123_),
    .Y(_06141_));
 sky130_fd_sc_hd__and3_2 _19073_ (.A(_06123_),
    .B(_06139_),
    .C(_06140_),
    .X(_06142_));
 sky130_fd_sc_hd__or3_2 _19074_ (.A(_11258_),
    .B(_06141_),
    .C(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__a21bo_2 _19075_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[4] ),
    .B1_N(_06143_),
    .X(_01478_));
 sky130_fd_sc_hd__and2b_2 _19076_ (.A_N(_06133_),
    .B(_06136_),
    .X(_06144_));
 sky130_fd_sc_hd__a21bo_2 _19077_ (.A1(_06125_),
    .A2(_06127_),
    .B1_N(_06126_),
    .X(_06145_));
 sky130_fd_sc_hd__a22oi_2 _19078_ (.A1(\systolic_inst.B_outs[7][1] ),
    .A2(\systolic_inst.A_outs[7][4] ),
    .B1(\systolic_inst.A_outs[7][5] ),
    .B2(\systolic_inst.B_outs[7][0] ),
    .Y(_06146_));
 sky130_fd_sc_hd__and4_2 _19079_ (.A(\systolic_inst.B_outs[7][0] ),
    .B(\systolic_inst.B_outs[7][1] ),
    .C(\systolic_inst.A_outs[7][4] ),
    .D(\systolic_inst.A_outs[7][5] ),
    .X(_06147_));
 sky130_fd_sc_hd__nor2_2 _19080_ (.A(_06146_),
    .B(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__xor2_2 _19081_ (.A(_06145_),
    .B(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__xor2_2 _19082_ (.A(_06132_),
    .B(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__and4_2 _19083_ (.A(\systolic_inst.A_outs[7][1] ),
    .B(\systolic_inst.A_outs[7][2] ),
    .C(\systolic_inst.B_outs[7][3] ),
    .D(\systolic_inst.B_outs[7][4] ),
    .X(_06151_));
 sky130_fd_sc_hd__a22oi_2 _19084_ (.A1(\systolic_inst.A_outs[7][2] ),
    .A2(\systolic_inst.B_outs[7][3] ),
    .B1(\systolic_inst.B_outs[7][4] ),
    .B2(\systolic_inst.A_outs[7][1] ),
    .Y(_06152_));
 sky130_fd_sc_hd__a22o_2 _19085_ (.A1(\systolic_inst.A_outs[7][2] ),
    .A2(\systolic_inst.B_outs[7][3] ),
    .B1(\systolic_inst.B_outs[7][4] ),
    .B2(\systolic_inst.A_outs[7][1] ),
    .X(_06153_));
 sky130_fd_sc_hd__and4b_2 _19086_ (.A_N(_06151_),
    .B(_06153_),
    .C(\systolic_inst.B_outs[7][2] ),
    .D(\systolic_inst.A_outs[7][3] ),
    .X(_06154_));
 sky130_fd_sc_hd__o2bb2a_2 _19087_ (.A1_N(\systolic_inst.B_outs[7][2] ),
    .A2_N(\systolic_inst.A_outs[7][3] ),
    .B1(_06151_),
    .B2(_06152_),
    .X(_06155_));
 sky130_fd_sc_hd__and4bb_2 _19088_ (.A_N(_06154_),
    .B_N(_06155_),
    .C(\systolic_inst.A_outs[7][0] ),
    .D(\systolic_inst.B_outs[7][5] ),
    .X(_06156_));
 sky130_fd_sc_hd__o2bb2a_2 _19089_ (.A1_N(\systolic_inst.A_outs[7][0] ),
    .A2_N(\systolic_inst.B_outs[7][5] ),
    .B1(_06154_),
    .B2(_06155_),
    .X(_06157_));
 sky130_fd_sc_hd__or2_2 _19090_ (.A(_06156_),
    .B(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__nor2_2 _19091_ (.A(_06150_),
    .B(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__xor2_2 _19092_ (.A(_06150_),
    .B(_06158_),
    .X(_06160_));
 sky130_fd_sc_hd__nand2_2 _19093_ (.A(_06137_),
    .B(_06160_),
    .Y(_06161_));
 sky130_fd_sc_hd__xor2_2 _19094_ (.A(_06137_),
    .B(_06160_),
    .X(_06162_));
 sky130_fd_sc_hd__nand2b_2 _19095_ (.A_N(_06144_),
    .B(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__xnor2_2 _19096_ (.A(_06144_),
    .B(_06162_),
    .Y(_06164_));
 sky130_fd_sc_hd__a21bo_2 _19097_ (.A1(_06123_),
    .A2(_06140_),
    .B1_N(_06139_),
    .X(_06165_));
 sky130_fd_sc_hd__nand2_2 _19098_ (.A(_06164_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__o21a_2 _19099_ (.A1(_06164_),
    .A2(_06165_),
    .B1(\systolic_inst.ce_local ),
    .X(_06167_));
 sky130_fd_sc_hd__a22o_2 _19100_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[5] ),
    .B1(_06166_),
    .B2(_06167_),
    .X(_01479_));
 sky130_fd_sc_hd__a32o_2 _19101_ (.A1(\systolic_inst.A_outs[7][4] ),
    .A2(_06131_),
    .A3(_06149_),
    .B1(_06148_),
    .B2(_06145_),
    .X(_06168_));
 sky130_fd_sc_hd__a31o_2 _19102_ (.A1(\systolic_inst.B_outs[7][2] ),
    .A2(\systolic_inst.A_outs[7][3] ),
    .A3(_06153_),
    .B1(_06151_),
    .X(_06169_));
 sky130_fd_sc_hd__a22oi_2 _19103_ (.A1(\systolic_inst.B_outs[7][1] ),
    .A2(\systolic_inst.A_outs[7][5] ),
    .B1(\systolic_inst.A_outs[7][6] ),
    .B2(\systolic_inst.B_outs[7][0] ),
    .Y(_06170_));
 sky130_fd_sc_hd__and4_2 _19104_ (.A(\systolic_inst.B_outs[7][0] ),
    .B(\systolic_inst.B_outs[7][1] ),
    .C(\systolic_inst.A_outs[7][5] ),
    .D(\systolic_inst.A_outs[7][6] ),
    .X(_06171_));
 sky130_fd_sc_hd__or2_2 _19105_ (.A(_06170_),
    .B(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__and2b_2 _19106_ (.A_N(_06172_),
    .B(_06169_),
    .X(_06173_));
 sky130_fd_sc_hd__xnor2_2 _19107_ (.A(_06169_),
    .B(_06172_),
    .Y(_06174_));
 sky130_fd_sc_hd__xor2_2 _19108_ (.A(_06147_),
    .B(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__nand4_2 _19109_ (.A(\systolic_inst.A_outs[7][2] ),
    .B(\systolic_inst.B_outs[7][3] ),
    .C(\systolic_inst.A_outs[7][3] ),
    .D(\systolic_inst.B_outs[7][4] ),
    .Y(_06176_));
 sky130_fd_sc_hd__a22o_2 _19110_ (.A1(\systolic_inst.B_outs[7][3] ),
    .A2(\systolic_inst.A_outs[7][3] ),
    .B1(\systolic_inst.B_outs[7][4] ),
    .B2(\systolic_inst.A_outs[7][2] ),
    .X(_06177_));
 sky130_fd_sc_hd__nand4_2 _19111_ (.A(\systolic_inst.B_outs[7][2] ),
    .B(\systolic_inst.A_outs[7][4] ),
    .C(_06176_),
    .D(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__a22o_2 _19112_ (.A1(\systolic_inst.B_outs[7][2] ),
    .A2(\systolic_inst.A_outs[7][4] ),
    .B1(_06176_),
    .B2(_06177_),
    .X(_06179_));
 sky130_fd_sc_hd__a22oi_2 _19113_ (.A1(\systolic_inst.A_outs[7][1] ),
    .A2(\systolic_inst.B_outs[7][5] ),
    .B1(\systolic_inst.B_outs[7][6] ),
    .B2(\systolic_inst.A_outs[7][0] ),
    .Y(_06180_));
 sky130_fd_sc_hd__nand2_2 _19114_ (.A(\systolic_inst.A_outs[7][1] ),
    .B(\systolic_inst.B_outs[7][6] ),
    .Y(_06181_));
 sky130_fd_sc_hd__and4_2 _19115_ (.A(\systolic_inst.A_outs[7][0] ),
    .B(\systolic_inst.A_outs[7][1] ),
    .C(\systolic_inst.B_outs[7][5] ),
    .D(\systolic_inst.B_outs[7][6] ),
    .X(_06182_));
 sky130_fd_sc_hd__nor2_2 _19116_ (.A(_06180_),
    .B(_06182_),
    .Y(_06183_));
 sky130_fd_sc_hd__nand3_2 _19117_ (.A(_06178_),
    .B(_06179_),
    .C(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__a21o_2 _19118_ (.A1(_06178_),
    .A2(_06179_),
    .B1(_06183_),
    .X(_06185_));
 sky130_fd_sc_hd__and3_2 _19119_ (.A(_06156_),
    .B(_06184_),
    .C(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__a21oi_2 _19120_ (.A1(_06184_),
    .A2(_06185_),
    .B1(_06156_),
    .Y(_06187_));
 sky130_fd_sc_hd__or3b_2 _19121_ (.A(_06186_),
    .B(_06187_),
    .C_N(_06175_),
    .X(_06188_));
 sky130_fd_sc_hd__o21bai_2 _19122_ (.A1(_06186_),
    .A2(_06187_),
    .B1_N(_06175_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand3_2 _19123_ (.A(_06159_),
    .B(_06188_),
    .C(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__a21o_2 _19124_ (.A1(_06188_),
    .A2(_06189_),
    .B1(_06159_),
    .X(_06191_));
 sky130_fd_sc_hd__and3_2 _19125_ (.A(_06168_),
    .B(_06190_),
    .C(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__a21oi_2 _19126_ (.A1(_06190_),
    .A2(_06191_),
    .B1(_06168_),
    .Y(_06193_));
 sky130_fd_sc_hd__a211oi_2 _19127_ (.A1(_06161_),
    .A2(_06163_),
    .B1(_06192_),
    .C1(_06193_),
    .Y(_06194_));
 sky130_fd_sc_hd__o211a_2 _19128_ (.A1(_06192_),
    .A2(_06193_),
    .B1(_06161_),
    .C1(_06163_),
    .X(_06195_));
 sky130_fd_sc_hd__nor2_2 _19129_ (.A(_06194_),
    .B(_06195_),
    .Y(_06196_));
 sky130_fd_sc_hd__xnor2_2 _19130_ (.A(_06166_),
    .B(_06196_),
    .Y(_06197_));
 sky130_fd_sc_hd__mux2_1 _19131_ (.A0(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[6] ),
    .A1(_06197_),
    .S(\systolic_inst.ce_local ),
    .X(_01480_));
 sky130_fd_sc_hd__a21boi_2 _19132_ (.A1(_06168_),
    .A2(_06191_),
    .B1_N(_06190_),
    .Y(_06198_));
 sky130_fd_sc_hd__a21oi_2 _19133_ (.A1(_06147_),
    .A2(_06174_),
    .B1(_06173_),
    .Y(_06199_));
 sky130_fd_sc_hd__nand2_2 _19134_ (.A(_06176_),
    .B(_06178_),
    .Y(_06200_));
 sky130_fd_sc_hd__a22o_2 _19135_ (.A1(\systolic_inst.B_outs[7][1] ),
    .A2(\systolic_inst.A_outs[7][6] ),
    .B1(\systolic_inst.A_outs[7][7] ),
    .B2(\systolic_inst.B_outs[7][0] ),
    .X(_06201_));
 sky130_fd_sc_hd__nand4_2 _19136_ (.A(\systolic_inst.B_outs[7][0] ),
    .B(\systolic_inst.B_outs[7][1] ),
    .C(\systolic_inst.A_outs[7][6] ),
    .D(\systolic_inst.A_outs[7][7] ),
    .Y(_06202_));
 sky130_fd_sc_hd__nand2_2 _19137_ (.A(_06201_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__xnor2_2 _19138_ (.A(_11261_),
    .B(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__nand2b_2 _19139_ (.A_N(_06204_),
    .B(_06200_),
    .Y(_06205_));
 sky130_fd_sc_hd__xnor2_2 _19140_ (.A(_06200_),
    .B(_06204_),
    .Y(_06206_));
 sky130_fd_sc_hd__xnor2_2 _19141_ (.A(_06171_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__nand2_2 _19142_ (.A(\systolic_inst.B_outs[7][2] ),
    .B(\systolic_inst.A_outs[7][5] ),
    .Y(_06208_));
 sky130_fd_sc_hd__and4_2 _19143_ (.A(\systolic_inst.B_outs[7][3] ),
    .B(\systolic_inst.A_outs[7][3] ),
    .C(\systolic_inst.B_outs[7][4] ),
    .D(\systolic_inst.A_outs[7][4] ),
    .X(_06209_));
 sky130_fd_sc_hd__a22oi_2 _19144_ (.A1(\systolic_inst.A_outs[7][3] ),
    .A2(\systolic_inst.B_outs[7][4] ),
    .B1(\systolic_inst.A_outs[7][4] ),
    .B2(\systolic_inst.B_outs[7][3] ),
    .Y(_06210_));
 sky130_fd_sc_hd__or2_2 _19145_ (.A(_06209_),
    .B(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__xnor2_2 _19146_ (.A(_06208_),
    .B(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2_2 _19147_ (.A(\systolic_inst.A_outs[7][2] ),
    .B(\systolic_inst.B_outs[7][5] ),
    .Y(_06213_));
 sky130_fd_sc_hd__and2b_2 _19148_ (.A_N(\systolic_inst.A_outs[7][0] ),
    .B(\systolic_inst.B_outs[7][7] ),
    .X(_06214_));
 sky130_fd_sc_hd__and3_2 _19149_ (.A(\systolic_inst.A_outs[7][1] ),
    .B(\systolic_inst.B_outs[7][6] ),
    .C(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__xnor2_2 _19150_ (.A(_06181_),
    .B(_06214_),
    .Y(_06216_));
 sky130_fd_sc_hd__xnor2_2 _19151_ (.A(_06213_),
    .B(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__xnor2_2 _19152_ (.A(_06182_),
    .B(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__nor2_2 _19153_ (.A(_06212_),
    .B(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__xnor2_2 _19154_ (.A(_06212_),
    .B(_06218_),
    .Y(_06220_));
 sky130_fd_sc_hd__or2_2 _19155_ (.A(_06184_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__and2_2 _19156_ (.A(_06184_),
    .B(_06220_),
    .X(_06222_));
 sky130_fd_sc_hd__xor2_2 _19157_ (.A(_06184_),
    .B(_06220_),
    .X(_06223_));
 sky130_fd_sc_hd__xnor2_2 _19158_ (.A(_06207_),
    .B(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__and2b_2 _19159_ (.A_N(_06186_),
    .B(_06188_),
    .X(_06225_));
 sky130_fd_sc_hd__and2b_2 _19160_ (.A_N(_06225_),
    .B(_06224_),
    .X(_06226_));
 sky130_fd_sc_hd__xnor2_2 _19161_ (.A(_06224_),
    .B(_06225_),
    .Y(_06227_));
 sky130_fd_sc_hd__and2b_2 _19162_ (.A_N(_06199_),
    .B(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__xnor2_2 _19163_ (.A(_06199_),
    .B(_06227_),
    .Y(_06229_));
 sky130_fd_sc_hd__and2b_2 _19164_ (.A_N(_06198_),
    .B(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__xnor2_2 _19165_ (.A(_06198_),
    .B(_06229_),
    .Y(_06231_));
 sky130_fd_sc_hd__a31o_2 _19166_ (.A1(_06164_),
    .A2(_06165_),
    .A3(_06196_),
    .B1(_06194_),
    .X(_06232_));
 sky130_fd_sc_hd__xor2_2 _19167_ (.A(_06231_),
    .B(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__mux2_1 _19168_ (.A0(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[7] ),
    .A1(_06233_),
    .S(\systolic_inst.ce_local ),
    .X(_01481_));
 sky130_fd_sc_hd__a21bo_2 _19169_ (.A1(_06171_),
    .A2(_06206_),
    .B1_N(_06205_),
    .X(_06234_));
 sky130_fd_sc_hd__a21bo_2 _19170_ (.A1(\systolic_inst.B_outs[7][7] ),
    .A2(_06201_),
    .B1_N(_06202_),
    .X(_06235_));
 sky130_fd_sc_hd__o21bai_2 _19171_ (.A1(_06208_),
    .A2(_06210_),
    .B1_N(_06209_),
    .Y(_06236_));
 sky130_fd_sc_hd__o21a_2 _19172_ (.A1(\systolic_inst.B_outs[7][0] ),
    .A2(\systolic_inst.B_outs[7][1] ),
    .B1(\systolic_inst.A_outs[7][7] ),
    .X(_06237_));
 sky130_fd_sc_hd__o21ai_2 _19173_ (.A1(\systolic_inst.B_outs[7][0] ),
    .A2(\systolic_inst.B_outs[7][1] ),
    .B1(\systolic_inst.A_outs[7][7] ),
    .Y(_06238_));
 sky130_fd_sc_hd__a21o_2 _19174_ (.A1(\systolic_inst.B_outs[7][0] ),
    .A2(\systolic_inst.B_outs[7][1] ),
    .B1(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__and2b_2 _19175_ (.A_N(_06239_),
    .B(_06236_),
    .X(_06240_));
 sky130_fd_sc_hd__xnor2_2 _19176_ (.A(_06236_),
    .B(_06239_),
    .Y(_06241_));
 sky130_fd_sc_hd__xnor2_2 _19177_ (.A(_06235_),
    .B(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__and4_2 _19178_ (.A(\systolic_inst.B_outs[7][3] ),
    .B(\systolic_inst.B_outs[7][4] ),
    .C(\systolic_inst.A_outs[7][4] ),
    .D(\systolic_inst.A_outs[7][5] ),
    .X(_06243_));
 sky130_fd_sc_hd__a22oi_2 _19179_ (.A1(\systolic_inst.B_outs[7][4] ),
    .A2(\systolic_inst.A_outs[7][4] ),
    .B1(\systolic_inst.A_outs[7][5] ),
    .B2(\systolic_inst.B_outs[7][3] ),
    .Y(_06244_));
 sky130_fd_sc_hd__nor2_2 _19180_ (.A(_06243_),
    .B(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__nand2_2 _19181_ (.A(\systolic_inst.B_outs[7][2] ),
    .B(\systolic_inst.A_outs[7][6] ),
    .Y(_06246_));
 sky130_fd_sc_hd__xnor2_2 _19182_ (.A(_06245_),
    .B(_06246_),
    .Y(_06247_));
 sky130_fd_sc_hd__nand2_2 _19183_ (.A(\systolic_inst.A_outs[7][3] ),
    .B(\systolic_inst.B_outs[7][5] ),
    .Y(_06248_));
 sky130_fd_sc_hd__and4b_2 _19184_ (.A_N(\systolic_inst.A_outs[7][1] ),
    .B(\systolic_inst.A_outs[7][2] ),
    .C(\systolic_inst.B_outs[7][6] ),
    .D(\systolic_inst.B_outs[7][7] ),
    .X(_06249_));
 sky130_fd_sc_hd__o2bb2a_2 _19185_ (.A1_N(\systolic_inst.A_outs[7][2] ),
    .A2_N(\systolic_inst.B_outs[7][6] ),
    .B1(_11261_),
    .B2(\systolic_inst.A_outs[7][1] ),
    .X(_06250_));
 sky130_fd_sc_hd__nor2_2 _19186_ (.A(_06249_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__xnor2_2 _19187_ (.A(_06248_),
    .B(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__a31oi_2 _19188_ (.A1(\systolic_inst.A_outs[7][2] ),
    .A2(\systolic_inst.B_outs[7][5] ),
    .A3(_06216_),
    .B1(_06215_),
    .Y(_06253_));
 sky130_fd_sc_hd__nand2b_2 _19189_ (.A_N(_06253_),
    .B(_06252_),
    .Y(_06254_));
 sky130_fd_sc_hd__xnor2_2 _19190_ (.A(_06252_),
    .B(_06253_),
    .Y(_06255_));
 sky130_fd_sc_hd__nand2_2 _19191_ (.A(_06247_),
    .B(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__xnor2_2 _19192_ (.A(_06247_),
    .B(_06255_),
    .Y(_06257_));
 sky130_fd_sc_hd__a21oi_2 _19193_ (.A1(_06182_),
    .A2(_06217_),
    .B1(_06219_),
    .Y(_06258_));
 sky130_fd_sc_hd__xnor2_2 _19194_ (.A(_06257_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__or2_2 _19195_ (.A(_06242_),
    .B(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__xor2_2 _19196_ (.A(_06242_),
    .B(_06259_),
    .X(_06261_));
 sky130_fd_sc_hd__o21a_2 _19197_ (.A1(_06207_),
    .A2(_06222_),
    .B1(_06221_),
    .X(_06262_));
 sky130_fd_sc_hd__nand2b_2 _19198_ (.A_N(_06262_),
    .B(_06261_),
    .Y(_06263_));
 sky130_fd_sc_hd__xor2_2 _19199_ (.A(_06261_),
    .B(_06262_),
    .X(_06264_));
 sky130_fd_sc_hd__nand2b_2 _19200_ (.A_N(_06264_),
    .B(_06234_),
    .Y(_06265_));
 sky130_fd_sc_hd__xor2_2 _19201_ (.A(_06234_),
    .B(_06264_),
    .X(_06266_));
 sky130_fd_sc_hd__nor2_2 _19202_ (.A(_06226_),
    .B(_06228_),
    .Y(_06267_));
 sky130_fd_sc_hd__nor2_2 _19203_ (.A(_06266_),
    .B(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__xor2_2 _19204_ (.A(_06266_),
    .B(_06267_),
    .X(_06269_));
 sky130_fd_sc_hd__a21o_2 _19205_ (.A1(_06231_),
    .A2(_06232_),
    .B1(_06230_),
    .X(_06270_));
 sky130_fd_sc_hd__xor2_2 _19206_ (.A(_06269_),
    .B(_06270_),
    .X(_06271_));
 sky130_fd_sc_hd__mux2_1 _19207_ (.A0(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[8] ),
    .A1(_06271_),
    .S(\systolic_inst.ce_local ),
    .X(_01482_));
 sky130_fd_sc_hd__a21o_2 _19208_ (.A1(_06235_),
    .A2(_06241_),
    .B1(_06240_),
    .X(_06272_));
 sky130_fd_sc_hd__o21ba_2 _19209_ (.A1(_06244_),
    .A2(_06246_),
    .B1_N(_06243_),
    .X(_06273_));
 sky130_fd_sc_hd__nor2_2 _19210_ (.A(_06238_),
    .B(_06273_),
    .Y(_06274_));
 sky130_fd_sc_hd__and2_2 _19211_ (.A(_06238_),
    .B(_06273_),
    .X(_06275_));
 sky130_fd_sc_hd__or2_2 _19212_ (.A(_06274_),
    .B(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__nand2_2 _19213_ (.A(\systolic_inst.B_outs[7][2] ),
    .B(\systolic_inst.A_outs[7][7] ),
    .Y(_06277_));
 sky130_fd_sc_hd__a22oi_2 _19214_ (.A1(\systolic_inst.B_outs[7][4] ),
    .A2(\systolic_inst.A_outs[7][5] ),
    .B1(\systolic_inst.A_outs[7][6] ),
    .B2(\systolic_inst.B_outs[7][3] ),
    .Y(_06278_));
 sky130_fd_sc_hd__and4_2 _19215_ (.A(\systolic_inst.B_outs[7][3] ),
    .B(\systolic_inst.B_outs[7][4] ),
    .C(\systolic_inst.A_outs[7][5] ),
    .D(\systolic_inst.A_outs[7][6] ),
    .X(_06279_));
 sky130_fd_sc_hd__nor2_2 _19216_ (.A(_06278_),
    .B(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__xnor2_2 _19217_ (.A(_06277_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2_2 _19218_ (.A(\systolic_inst.A_outs[7][4] ),
    .B(\systolic_inst.B_outs[7][5] ),
    .Y(_06282_));
 sky130_fd_sc_hd__and4b_2 _19219_ (.A_N(\systolic_inst.A_outs[7][2] ),
    .B(\systolic_inst.A_outs[7][3] ),
    .C(\systolic_inst.B_outs[7][6] ),
    .D(\systolic_inst.B_outs[7][7] ),
    .X(_06283_));
 sky130_fd_sc_hd__o2bb2a_2 _19220_ (.A1_N(\systolic_inst.A_outs[7][3] ),
    .A2_N(\systolic_inst.B_outs[7][6] ),
    .B1(_11261_),
    .B2(\systolic_inst.A_outs[7][2] ),
    .X(_06284_));
 sky130_fd_sc_hd__nor2_2 _19221_ (.A(_06283_),
    .B(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__xnor2_2 _19222_ (.A(_06282_),
    .B(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__o21ba_2 _19223_ (.A1(_06248_),
    .A2(_06250_),
    .B1_N(_06249_),
    .X(_06287_));
 sky130_fd_sc_hd__nand2b_2 _19224_ (.A_N(_06287_),
    .B(_06286_),
    .Y(_06288_));
 sky130_fd_sc_hd__xnor2_2 _19225_ (.A(_06286_),
    .B(_06287_),
    .Y(_06289_));
 sky130_fd_sc_hd__xnor2_2 _19226_ (.A(_06281_),
    .B(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__a21o_2 _19227_ (.A1(_06254_),
    .A2(_06256_),
    .B1(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__nand3_2 _19228_ (.A(_06254_),
    .B(_06256_),
    .C(_06290_),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_2 _19229_ (.A(_06291_),
    .B(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__xor2_2 _19230_ (.A(_06276_),
    .B(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__o21a_2 _19231_ (.A1(_06257_),
    .A2(_06258_),
    .B1(_06260_),
    .X(_06295_));
 sky130_fd_sc_hd__nand2b_2 _19232_ (.A_N(_06295_),
    .B(_06294_),
    .Y(_06296_));
 sky130_fd_sc_hd__xnor2_2 _19233_ (.A(_06294_),
    .B(_06295_),
    .Y(_06297_));
 sky130_fd_sc_hd__xnor2_2 _19234_ (.A(_06272_),
    .B(_06297_),
    .Y(_06298_));
 sky130_fd_sc_hd__a21o_2 _19235_ (.A1(_06263_),
    .A2(_06265_),
    .B1(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__nand3_2 _19236_ (.A(_06263_),
    .B(_06265_),
    .C(_06298_),
    .Y(_06300_));
 sky130_fd_sc_hd__a21o_2 _19237_ (.A1(_06269_),
    .A2(_06270_),
    .B1(_06268_),
    .X(_06301_));
 sky130_fd_sc_hd__and3_2 _19238_ (.A(_06299_),
    .B(_06300_),
    .C(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__a21oi_2 _19239_ (.A1(_06299_),
    .A2(_06300_),
    .B1(_06301_),
    .Y(_06303_));
 sky130_fd_sc_hd__nor2_2 _19240_ (.A(_06302_),
    .B(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__mux2_1 _19241_ (.A0(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[9] ),
    .A1(_06304_),
    .S(\systolic_inst.ce_local ),
    .X(_01483_));
 sky130_fd_sc_hd__o21ba_2 _19242_ (.A1(_06277_),
    .A2(_06278_),
    .B1_N(_06279_),
    .X(_06305_));
 sky130_fd_sc_hd__nor2_2 _19243_ (.A(_06238_),
    .B(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__and2_2 _19244_ (.A(_06238_),
    .B(_06305_),
    .X(_06307_));
 sky130_fd_sc_hd__or2_2 _19245_ (.A(_06306_),
    .B(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__a22o_2 _19246_ (.A1(\systolic_inst.B_outs[7][4] ),
    .A2(\systolic_inst.A_outs[7][6] ),
    .B1(\systolic_inst.A_outs[7][7] ),
    .B2(\systolic_inst.B_outs[7][3] ),
    .X(_06309_));
 sky130_fd_sc_hd__and3_2 _19247_ (.A(\systolic_inst.B_outs[7][3] ),
    .B(\systolic_inst.B_outs[7][4] ),
    .C(\systolic_inst.A_outs[7][7] ),
    .X(_06310_));
 sky130_fd_sc_hd__a21bo_2 _19248_ (.A1(\systolic_inst.A_outs[7][6] ),
    .A2(_06310_),
    .B1_N(_06309_),
    .X(_06311_));
 sky130_fd_sc_hd__xor2_2 _19249_ (.A(_06277_),
    .B(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__nand2_2 _19250_ (.A(\systolic_inst.B_outs[7][5] ),
    .B(\systolic_inst.A_outs[7][5] ),
    .Y(_06313_));
 sky130_fd_sc_hd__and4b_2 _19251_ (.A_N(\systolic_inst.A_outs[7][3] ),
    .B(\systolic_inst.A_outs[7][4] ),
    .C(\systolic_inst.B_outs[7][6] ),
    .D(\systolic_inst.B_outs[7][7] ),
    .X(_06314_));
 sky130_fd_sc_hd__o2bb2a_2 _19252_ (.A1_N(\systolic_inst.A_outs[7][4] ),
    .A2_N(\systolic_inst.B_outs[7][6] ),
    .B1(_11261_),
    .B2(\systolic_inst.A_outs[7][3] ),
    .X(_06315_));
 sky130_fd_sc_hd__nor2_2 _19253_ (.A(_06314_),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__xnor2_2 _19254_ (.A(_06313_),
    .B(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__o21ba_2 _19255_ (.A1(_06282_),
    .A2(_06284_),
    .B1_N(_06283_),
    .X(_06318_));
 sky130_fd_sc_hd__nand2b_2 _19256_ (.A_N(_06318_),
    .B(_06317_),
    .Y(_06319_));
 sky130_fd_sc_hd__xnor2_2 _19257_ (.A(_06317_),
    .B(_06318_),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_2 _19258_ (.A(_06312_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__or2_2 _19259_ (.A(_06312_),
    .B(_06320_),
    .X(_06322_));
 sky130_fd_sc_hd__nand2_2 _19260_ (.A(_06321_),
    .B(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__a21bo_2 _19261_ (.A1(_06281_),
    .A2(_06289_),
    .B1_N(_06288_),
    .X(_06324_));
 sky130_fd_sc_hd__nand2b_2 _19262_ (.A_N(_06323_),
    .B(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__xor2_2 _19263_ (.A(_06323_),
    .B(_06324_),
    .X(_06326_));
 sky130_fd_sc_hd__xor2_2 _19264_ (.A(_06308_),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__o21a_2 _19265_ (.A1(_06276_),
    .A2(_06293_),
    .B1(_06291_),
    .X(_06328_));
 sky130_fd_sc_hd__nand2b_2 _19266_ (.A_N(_06328_),
    .B(_06327_),
    .Y(_06329_));
 sky130_fd_sc_hd__xnor2_2 _19267_ (.A(_06327_),
    .B(_06328_),
    .Y(_06330_));
 sky130_fd_sc_hd__nand2_2 _19268_ (.A(_06274_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__or2_2 _19269_ (.A(_06274_),
    .B(_06330_),
    .X(_06332_));
 sky130_fd_sc_hd__nand2_2 _19270_ (.A(_06331_),
    .B(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__a21boi_2 _19271_ (.A1(_06272_),
    .A2(_06297_),
    .B1_N(_06296_),
    .Y(_06334_));
 sky130_fd_sc_hd__nor2_2 _19272_ (.A(_06333_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__xnor2_2 _19273_ (.A(_06333_),
    .B(_06334_),
    .Y(_06336_));
 sky130_fd_sc_hd__nand2_2 _19274_ (.A(_06300_),
    .B(_06301_),
    .Y(_06337_));
 sky130_fd_sc_hd__and3_2 _19275_ (.A(_06299_),
    .B(_06336_),
    .C(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__a21oi_2 _19276_ (.A1(_06299_),
    .A2(_06337_),
    .B1(_06336_),
    .Y(_06339_));
 sky130_fd_sc_hd__or2_2 _19277_ (.A(_11258_),
    .B(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__a2bb2o_2 _19278_ (.A1_N(_06340_),
    .A2_N(_06338_),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[10] ),
    .B2(_11258_),
    .X(_01484_));
 sky130_fd_sc_hd__or2_2 _19279_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[11] ),
    .X(_06341_));
 sky130_fd_sc_hd__o2bb2a_2 _19280_ (.A1_N(\systolic_inst.A_outs[7][6] ),
    .A2_N(_06310_),
    .B1(_06311_),
    .B2(_06277_),
    .X(_06342_));
 sky130_fd_sc_hd__or2_2 _19281_ (.A(_06238_),
    .B(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__nand2_2 _19282_ (.A(_06238_),
    .B(_06342_),
    .Y(_06344_));
 sky130_fd_sc_hd__nand2_2 _19283_ (.A(_06343_),
    .B(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__or2_2 _19284_ (.A(\systolic_inst.B_outs[7][3] ),
    .B(\systolic_inst.B_outs[7][4] ),
    .X(_06346_));
 sky130_fd_sc_hd__and3b_2 _19285_ (.A_N(_06310_),
    .B(_06346_),
    .C(\systolic_inst.A_outs[7][7] ),
    .X(_06347_));
 sky130_fd_sc_hd__xnor2_2 _19286_ (.A(_06277_),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__nand2_2 _19287_ (.A(\systolic_inst.B_outs[7][5] ),
    .B(\systolic_inst.A_outs[7][6] ),
    .Y(_06349_));
 sky130_fd_sc_hd__and4b_2 _19288_ (.A_N(\systolic_inst.A_outs[7][4] ),
    .B(\systolic_inst.A_outs[7][5] ),
    .C(\systolic_inst.B_outs[7][6] ),
    .D(\systolic_inst.B_outs[7][7] ),
    .X(_06350_));
 sky130_fd_sc_hd__o2bb2a_2 _19289_ (.A1_N(\systolic_inst.A_outs[7][5] ),
    .A2_N(\systolic_inst.B_outs[7][6] ),
    .B1(_11261_),
    .B2(\systolic_inst.A_outs[7][4] ),
    .X(_06351_));
 sky130_fd_sc_hd__or2_2 _19290_ (.A(_06350_),
    .B(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__xor2_2 _19291_ (.A(_06349_),
    .B(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__o21ba_2 _19292_ (.A1(_06313_),
    .A2(_06315_),
    .B1_N(_06314_),
    .X(_06354_));
 sky130_fd_sc_hd__nand2b_2 _19293_ (.A_N(_06354_),
    .B(_06353_),
    .Y(_06355_));
 sky130_fd_sc_hd__xnor2_2 _19294_ (.A(_06353_),
    .B(_06354_),
    .Y(_06356_));
 sky130_fd_sc_hd__nand2_2 _19295_ (.A(_06348_),
    .B(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__xnor2_2 _19296_ (.A(_06348_),
    .B(_06356_),
    .Y(_06358_));
 sky130_fd_sc_hd__a21o_2 _19297_ (.A1(_06319_),
    .A2(_06321_),
    .B1(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__nand3_2 _19298_ (.A(_06319_),
    .B(_06321_),
    .C(_06358_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand2_2 _19299_ (.A(_06359_),
    .B(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__xor2_2 _19300_ (.A(_06345_),
    .B(_06361_),
    .X(_06362_));
 sky130_fd_sc_hd__o21a_2 _19301_ (.A1(_06308_),
    .A2(_06326_),
    .B1(_06325_),
    .X(_06363_));
 sky130_fd_sc_hd__and2b_2 _19302_ (.A_N(_06363_),
    .B(_06362_),
    .X(_06364_));
 sky130_fd_sc_hd__xnor2_2 _19303_ (.A(_06362_),
    .B(_06363_),
    .Y(_06365_));
 sky130_fd_sc_hd__xnor2_2 _19304_ (.A(_06306_),
    .B(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__and3_2 _19305_ (.A(_06329_),
    .B(_06331_),
    .C(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__inv_2 _19306_ (.A(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__a21oi_2 _19307_ (.A1(_06329_),
    .A2(_06331_),
    .B1(_06366_),
    .Y(_06369_));
 sky130_fd_sc_hd__nor4_2 _19308_ (.A(_06335_),
    .B(_06339_),
    .C(_06367_),
    .D(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__o22a_2 _19309_ (.A1(_06335_),
    .A2(_06339_),
    .B1(_06367_),
    .B2(_06369_),
    .X(_06371_));
 sky130_fd_sc_hd__o31a_2 _19310_ (.A1(_11258_),
    .A2(_06370_),
    .A3(_06371_),
    .B1(_06341_),
    .X(_01485_));
 sky130_fd_sc_hd__a31o_2 _19311_ (.A1(\systolic_inst.B_outs[7][2] ),
    .A2(\systolic_inst.A_outs[7][7] ),
    .A3(_06346_),
    .B1(_06310_),
    .X(_06372_));
 sky130_fd_sc_hd__or2_2 _19312_ (.A(_06237_),
    .B(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__nand2_2 _19313_ (.A(_06237_),
    .B(_06372_),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_2 _19314_ (.A(_06373_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__inv_2 _19315_ (.A(_06375_),
    .Y(_06376_));
 sky130_fd_sc_hd__o2bb2a_2 _19316_ (.A1_N(\systolic_inst.B_outs[7][6] ),
    .A2_N(\systolic_inst.A_outs[7][6] ),
    .B1(_11261_),
    .B2(\systolic_inst.A_outs[7][5] ),
    .X(_06377_));
 sky130_fd_sc_hd__and4b_2 _19317_ (.A_N(\systolic_inst.A_outs[7][5] ),
    .B(\systolic_inst.B_outs[7][6] ),
    .C(\systolic_inst.A_outs[7][6] ),
    .D(\systolic_inst.B_outs[7][7] ),
    .X(_06378_));
 sky130_fd_sc_hd__nor2_2 _19318_ (.A(_06377_),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__nand2_2 _19319_ (.A(\systolic_inst.B_outs[7][5] ),
    .B(\systolic_inst.A_outs[7][7] ),
    .Y(_06380_));
 sky130_fd_sc_hd__xnor2_2 _19320_ (.A(_06379_),
    .B(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__o21ba_2 _19321_ (.A1(_06349_),
    .A2(_06351_),
    .B1_N(_06350_),
    .X(_06382_));
 sky130_fd_sc_hd__nand2b_2 _19322_ (.A_N(_06382_),
    .B(_06381_),
    .Y(_06383_));
 sky130_fd_sc_hd__xnor2_2 _19323_ (.A(_06381_),
    .B(_06382_),
    .Y(_06384_));
 sky130_fd_sc_hd__xnor2_2 _19324_ (.A(_06348_),
    .B(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__a21o_2 _19325_ (.A1(_06355_),
    .A2(_06357_),
    .B1(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__nand3_2 _19326_ (.A(_06355_),
    .B(_06357_),
    .C(_06385_),
    .Y(_06387_));
 sky130_fd_sc_hd__nand2_2 _19327_ (.A(_06386_),
    .B(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__xnor2_2 _19328_ (.A(_06376_),
    .B(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__o21a_2 _19329_ (.A1(_06345_),
    .A2(_06361_),
    .B1(_06359_),
    .X(_06390_));
 sky130_fd_sc_hd__and2b_2 _19330_ (.A_N(_06390_),
    .B(_06389_),
    .X(_06391_));
 sky130_fd_sc_hd__xnor2_2 _19331_ (.A(_06389_),
    .B(_06390_),
    .Y(_06392_));
 sky130_fd_sc_hd__and2b_2 _19332_ (.A_N(_06343_),
    .B(_06392_),
    .X(_06393_));
 sky130_fd_sc_hd__xor2_2 _19333_ (.A(_06343_),
    .B(_06392_),
    .X(_06394_));
 sky130_fd_sc_hd__a21oi_2 _19334_ (.A1(_06306_),
    .A2(_06365_),
    .B1(_06364_),
    .Y(_06395_));
 sky130_fd_sc_hd__nor2_2 _19335_ (.A(_06394_),
    .B(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__and2_2 _19336_ (.A(_06394_),
    .B(_06395_),
    .X(_06397_));
 sky130_fd_sc_hd__or2_2 _19337_ (.A(_06396_),
    .B(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__inv_2 _19338_ (.A(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__o31a_2 _19339_ (.A1(_06335_),
    .A2(_06339_),
    .A3(_06369_),
    .B1(_06368_),
    .X(_06400_));
 sky130_fd_sc_hd__o311a_2 _19340_ (.A1(_06335_),
    .A2(_06339_),
    .A3(_06369_),
    .B1(_06399_),
    .C1(_06368_),
    .X(_06401_));
 sky130_fd_sc_hd__nor2_2 _19341_ (.A(_06399_),
    .B(_06400_),
    .Y(_06402_));
 sky130_fd_sc_hd__nor2_2 _19342_ (.A(_06401_),
    .B(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__mux2_1 _19343_ (.A0(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[12] ),
    .A1(_06403_),
    .S(\systolic_inst.ce_local ),
    .X(_01486_));
 sky130_fd_sc_hd__nand2_2 _19344_ (.A(\systolic_inst.B_outs[7][6] ),
    .B(\systolic_inst.A_outs[7][7] ),
    .Y(_06404_));
 sky130_fd_sc_hd__or2_2 _19345_ (.A(\systolic_inst.A_outs[7][6] ),
    .B(_11261_),
    .X(_06405_));
 sky130_fd_sc_hd__and2_2 _19346_ (.A(_06404_),
    .B(_06405_),
    .X(_06406_));
 sky130_fd_sc_hd__nor2_2 _19347_ (.A(_06404_),
    .B(_06405_),
    .Y(_06407_));
 sky130_fd_sc_hd__nor2_2 _19348_ (.A(_06406_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__xnor2_2 _19349_ (.A(_06380_),
    .B(_06408_),
    .Y(_06409_));
 sky130_fd_sc_hd__o21ba_2 _19350_ (.A1(_06377_),
    .A2(_06380_),
    .B1_N(_06378_),
    .X(_06410_));
 sky130_fd_sc_hd__nand2b_2 _19351_ (.A_N(_06410_),
    .B(_06409_),
    .Y(_06411_));
 sky130_fd_sc_hd__xnor2_2 _19352_ (.A(_06409_),
    .B(_06410_),
    .Y(_06412_));
 sky130_fd_sc_hd__nand2_2 _19353_ (.A(_06348_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__or2_2 _19354_ (.A(_06348_),
    .B(_06412_),
    .X(_06414_));
 sky130_fd_sc_hd__nand2_2 _19355_ (.A(_06413_),
    .B(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__a21bo_2 _19356_ (.A1(_06348_),
    .A2(_06384_),
    .B1_N(_06383_),
    .X(_06416_));
 sky130_fd_sc_hd__nand2b_2 _19357_ (.A_N(_06415_),
    .B(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__xor2_2 _19358_ (.A(_06415_),
    .B(_06416_),
    .X(_06418_));
 sky130_fd_sc_hd__xnor2_2 _19359_ (.A(_06376_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__o21a_2 _19360_ (.A1(_06375_),
    .A2(_06388_),
    .B1(_06386_),
    .X(_06420_));
 sky130_fd_sc_hd__and2b_2 _19361_ (.A_N(_06420_),
    .B(_06419_),
    .X(_06421_));
 sky130_fd_sc_hd__and2b_2 _19362_ (.A_N(_06419_),
    .B(_06420_),
    .X(_06422_));
 sky130_fd_sc_hd__nor2_2 _19363_ (.A(_06421_),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__xnor2_2 _19364_ (.A(_06374_),
    .B(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__nor3_2 _19365_ (.A(_06391_),
    .B(_06393_),
    .C(_06424_),
    .Y(_06425_));
 sky130_fd_sc_hd__o21a_2 _19366_ (.A1(_06391_),
    .A2(_06393_),
    .B1(_06424_),
    .X(_06426_));
 sky130_fd_sc_hd__nor2_2 _19367_ (.A(_06425_),
    .B(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__o21ai_2 _19368_ (.A1(_06396_),
    .A2(_06401_),
    .B1(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__o31a_2 _19369_ (.A1(_06396_),
    .A2(_06401_),
    .A3(_06427_),
    .B1(\systolic_inst.ce_local ),
    .X(_06429_));
 sky130_fd_sc_hd__a22o_2 _19370_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[13] ),
    .B1(_06428_),
    .B2(_06429_),
    .X(_01487_));
 sky130_fd_sc_hd__a31o_2 _19371_ (.A1(\systolic_inst.B_outs[7][5] ),
    .A2(\systolic_inst.A_outs[7][7] ),
    .A3(_06408_),
    .B1(_06407_),
    .X(_06430_));
 sky130_fd_sc_hd__nand3_2 _19372_ (.A(\systolic_inst.B_outs[7][5] ),
    .B(\systolic_inst.B_outs[7][6] ),
    .C(\systolic_inst.A_outs[7][7] ),
    .Y(_06431_));
 sky130_fd_sc_hd__o211a_2 _19373_ (.A1(_11261_),
    .A2(\systolic_inst.A_outs[7][7] ),
    .B1(_06380_),
    .C1(_06404_),
    .X(_06432_));
 sky130_fd_sc_hd__a21oi_2 _19374_ (.A1(_06430_),
    .A2(_06431_),
    .B1(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__or2_2 _19375_ (.A(_06348_),
    .B(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__nand2_2 _19376_ (.A(_06348_),
    .B(_06433_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2_2 _19377_ (.A(_06434_),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__a21oi_2 _19378_ (.A1(_06411_),
    .A2(_06413_),
    .B1(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__and3_2 _19379_ (.A(_06411_),
    .B(_06413_),
    .C(_06436_),
    .X(_06438_));
 sky130_fd_sc_hd__nor2_2 _19380_ (.A(_06437_),
    .B(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__xnor2_2 _19381_ (.A(_06375_),
    .B(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__o21a_2 _19382_ (.A1(_06375_),
    .A2(_06418_),
    .B1(_06417_),
    .X(_06441_));
 sky130_fd_sc_hd__and2b_2 _19383_ (.A_N(_06441_),
    .B(_06440_),
    .X(_06442_));
 sky130_fd_sc_hd__and2b_2 _19384_ (.A_N(_06440_),
    .B(_06441_),
    .X(_06443_));
 sky130_fd_sc_hd__nor2_2 _19385_ (.A(_06442_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__xnor2_2 _19386_ (.A(_06374_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__o21ba_2 _19387_ (.A1(_06374_),
    .A2(_06422_),
    .B1_N(_06421_),
    .X(_06446_));
 sky130_fd_sc_hd__nand2b_2 _19388_ (.A_N(_06446_),
    .B(_06445_),
    .Y(_06447_));
 sky130_fd_sc_hd__xnor2_2 _19389_ (.A(_06445_),
    .B(_06446_),
    .Y(_06448_));
 sky130_fd_sc_hd__nor2_2 _19390_ (.A(_06396_),
    .B(_06426_),
    .Y(_06449_));
 sky130_fd_sc_hd__a2bb2o_2 _19391_ (.A1_N(_06425_),
    .A2_N(_06449_),
    .B1(_06427_),
    .B2(_06401_),
    .X(_06450_));
 sky130_fd_sc_hd__nand2_2 _19392_ (.A(_06448_),
    .B(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__xor2_2 _19393_ (.A(_06448_),
    .B(_06450_),
    .X(_06452_));
 sky130_fd_sc_hd__mux2_1 _19394_ (.A0(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[14] ),
    .A1(_06452_),
    .S(\systolic_inst.ce_local ),
    .X(_01488_));
 sky130_fd_sc_hd__a31o_2 _19395_ (.A1(_06237_),
    .A2(_06372_),
    .A3(_06444_),
    .B1(_06442_),
    .X(_06453_));
 sky130_fd_sc_hd__a21oi_2 _19396_ (.A1(_06376_),
    .A2(_06439_),
    .B1(_06437_),
    .Y(_06454_));
 sky130_fd_sc_hd__xnor2_2 _19397_ (.A(_06373_),
    .B(_06434_),
    .Y(_06455_));
 sky130_fd_sc_hd__xnor2_2 _19398_ (.A(_06454_),
    .B(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__xnor2_2 _19399_ (.A(_06453_),
    .B(_06456_),
    .Y(_06457_));
 sky130_fd_sc_hd__and3_2 _19400_ (.A(\systolic_inst.ce_local ),
    .B(_06447_),
    .C(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__a22o_2 _19401_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B1(_06451_),
    .B2(_06458_),
    .X(_01489_));
 sky130_fd_sc_hd__a21o_2 _19402_ (.A1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[7][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_06459_));
 sky130_fd_sc_hd__a21oi_2 _19403_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[7][0] ),
    .Y(_06460_));
 sky130_fd_sc_hd__a21oi_2 _19404_ (.A1(\systolic_inst.ce_local ),
    .A2(_06459_),
    .B1(_06460_),
    .Y(_01490_));
 sky130_fd_sc_hd__and2_2 _19405_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[7][1] ),
    .X(_06461_));
 sky130_fd_sc_hd__nand2_2 _19406_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[7][1] ),
    .Y(_06462_));
 sky130_fd_sc_hd__or2_2 _19407_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[7][1] ),
    .X(_06463_));
 sky130_fd_sc_hd__and4_2 _19408_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[7][0] ),
    .C(_06462_),
    .D(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__inv_2 _19409_ (.A(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__a22o_2 _19410_ (.A1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[7][0] ),
    .B1(_06462_),
    .B2(_06463_),
    .X(_06466_));
 sky130_fd_sc_hd__a32o_2 _19411_ (.A1(_11712_),
    .A2(_06465_),
    .A3(_06466_),
    .B1(\systolic_inst.acc_wires[7][1] ),
    .B2(_11258_),
    .X(_01491_));
 sky130_fd_sc_hd__and2_2 _19412_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[7][2] ),
    .X(_06467_));
 sky130_fd_sc_hd__nand2_2 _19413_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[7][2] ),
    .Y(_06468_));
 sky130_fd_sc_hd__or2_2 _19414_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[7][2] ),
    .X(_06469_));
 sky130_fd_sc_hd__a211o_2 _19415_ (.A1(_06468_),
    .A2(_06469_),
    .B1(_06461_),
    .C1(_06464_),
    .X(_06470_));
 sky130_fd_sc_hd__o211a_2 _19416_ (.A1(_06461_),
    .A2(_06464_),
    .B1(_06468_),
    .C1(_06469_),
    .X(_06471_));
 sky130_fd_sc_hd__inv_2 _19417_ (.A(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__a32o_2 _19418_ (.A1(_11712_),
    .A2(_06470_),
    .A3(_06472_),
    .B1(\systolic_inst.acc_wires[7][2] ),
    .B2(_11258_),
    .X(_01492_));
 sky130_fd_sc_hd__and2_2 _19419_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[7][3] ),
    .X(_06473_));
 sky130_fd_sc_hd__nand2_2 _19420_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[7][3] ),
    .Y(_06474_));
 sky130_fd_sc_hd__or2_2 _19421_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[7][3] ),
    .X(_06475_));
 sky130_fd_sc_hd__a211o_2 _19422_ (.A1(_06474_),
    .A2(_06475_),
    .B1(_06467_),
    .C1(_06471_),
    .X(_06476_));
 sky130_fd_sc_hd__o211a_2 _19423_ (.A1(_06467_),
    .A2(_06471_),
    .B1(_06474_),
    .C1(_06475_),
    .X(_06477_));
 sky130_fd_sc_hd__inv_2 _19424_ (.A(_06477_),
    .Y(_06478_));
 sky130_fd_sc_hd__a32o_2 _19425_ (.A1(_11712_),
    .A2(_06476_),
    .A3(_06478_),
    .B1(\systolic_inst.acc_wires[7][3] ),
    .B2(_11258_),
    .X(_01493_));
 sky130_fd_sc_hd__and2_2 _19426_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[7][4] ),
    .X(_06479_));
 sky130_fd_sc_hd__nand2_2 _19427_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[7][4] ),
    .Y(_06480_));
 sky130_fd_sc_hd__or2_2 _19428_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[7][4] ),
    .X(_06481_));
 sky130_fd_sc_hd__a211o_2 _19429_ (.A1(_06480_),
    .A2(_06481_),
    .B1(_06473_),
    .C1(_06477_),
    .X(_06482_));
 sky130_fd_sc_hd__o211a_2 _19430_ (.A1(_06473_),
    .A2(_06477_),
    .B1(_06480_),
    .C1(_06481_),
    .X(_06483_));
 sky130_fd_sc_hd__inv_2 _19431_ (.A(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__a32o_2 _19432_ (.A1(_11712_),
    .A2(_06482_),
    .A3(_06484_),
    .B1(\systolic_inst.acc_wires[7][4] ),
    .B2(_11258_),
    .X(_01494_));
 sky130_fd_sc_hd__and2_2 _19433_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[7][5] ),
    .X(_06485_));
 sky130_fd_sc_hd__nand2_2 _19434_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[7][5] ),
    .Y(_06486_));
 sky130_fd_sc_hd__or2_2 _19435_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[7][5] ),
    .X(_06487_));
 sky130_fd_sc_hd__a211o_2 _19436_ (.A1(_06486_),
    .A2(_06487_),
    .B1(_06479_),
    .C1(_06483_),
    .X(_06488_));
 sky130_fd_sc_hd__o211a_2 _19437_ (.A1(_06479_),
    .A2(_06483_),
    .B1(_06486_),
    .C1(_06487_),
    .X(_06489_));
 sky130_fd_sc_hd__inv_2 _19438_ (.A(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__a32o_2 _19439_ (.A1(_11712_),
    .A2(_06488_),
    .A3(_06490_),
    .B1(\systolic_inst.acc_wires[7][5] ),
    .B2(_11258_),
    .X(_01495_));
 sky130_fd_sc_hd__and2_2 _19440_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[7][6] ),
    .X(_06491_));
 sky130_fd_sc_hd__nand2_2 _19441_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[7][6] ),
    .Y(_06492_));
 sky130_fd_sc_hd__or2_2 _19442_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[7][6] ),
    .X(_06493_));
 sky130_fd_sc_hd__a211o_2 _19443_ (.A1(_06492_),
    .A2(_06493_),
    .B1(_06485_),
    .C1(_06489_),
    .X(_06494_));
 sky130_fd_sc_hd__o211a_2 _19444_ (.A1(_06485_),
    .A2(_06489_),
    .B1(_06492_),
    .C1(_06493_),
    .X(_06495_));
 sky130_fd_sc_hd__inv_2 _19445_ (.A(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__a32o_2 _19446_ (.A1(_11712_),
    .A2(_06494_),
    .A3(_06496_),
    .B1(\systolic_inst.acc_wires[7][6] ),
    .B2(_11258_),
    .X(_01496_));
 sky130_fd_sc_hd__nand2_2 _19447_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[7][7] ),
    .Y(_06497_));
 sky130_fd_sc_hd__or2_2 _19448_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[7][7] ),
    .X(_06498_));
 sky130_fd_sc_hd__a211o_2 _19449_ (.A1(_06497_),
    .A2(_06498_),
    .B1(_06491_),
    .C1(_06495_),
    .X(_06499_));
 sky130_fd_sc_hd__o211ai_2 _19450_ (.A1(_06491_),
    .A2(_06495_),
    .B1(_06497_),
    .C1(_06498_),
    .Y(_06500_));
 sky130_fd_sc_hd__a32o_2 _19451_ (.A1(_11712_),
    .A2(_06499_),
    .A3(_06500_),
    .B1(\systolic_inst.acc_wires[7][7] ),
    .B2(_11258_),
    .X(_01497_));
 sky130_fd_sc_hd__and2_2 _19452_ (.A(_06497_),
    .B(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__nand2_2 _19453_ (.A(_06497_),
    .B(_06500_),
    .Y(_06502_));
 sky130_fd_sc_hd__nor2_2 _19454_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[7][8] ),
    .Y(_06503_));
 sky130_fd_sc_hd__and2_2 _19455_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[7][8] ),
    .X(_06504_));
 sky130_fd_sc_hd__nor2_2 _19456_ (.A(_06503_),
    .B(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__xnor2_2 _19457_ (.A(_06501_),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__a22o_2 _19458_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][8] ),
    .B1(_11712_),
    .B2(_06506_),
    .X(_01498_));
 sky130_fd_sc_hd__xor2_2 _19459_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[7][9] ),
    .X(_06507_));
 sky130_fd_sc_hd__a211o_2 _19460_ (.A1(_06502_),
    .A2(_06505_),
    .B1(_06507_),
    .C1(_06504_),
    .X(_06508_));
 sky130_fd_sc_hd__nand2_2 _19461_ (.A(_06505_),
    .B(_06507_),
    .Y(_06509_));
 sky130_fd_sc_hd__or2_2 _19462_ (.A(_06501_),
    .B(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__and2_2 _19463_ (.A(_06504_),
    .B(_06507_),
    .X(_06511_));
 sky130_fd_sc_hd__nor2_2 _19464_ (.A(_11713_),
    .B(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__a32o_2 _19465_ (.A1(_06508_),
    .A2(_06510_),
    .A3(_06512_),
    .B1(\systolic_inst.acc_wires[7][9] ),
    .B2(_11258_),
    .X(_01499_));
 sky130_fd_sc_hd__nand2_2 _19466_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[7][10] ),
    .Y(_06513_));
 sky130_fd_sc_hd__or2_2 _19467_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[7][10] ),
    .X(_06514_));
 sky130_fd_sc_hd__and2_2 _19468_ (.A(_06513_),
    .B(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__a21oi_2 _19469_ (.A1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[7][9] ),
    .B1(_06511_),
    .Y(_06516_));
 sky130_fd_sc_hd__nand2_2 _19470_ (.A(_06510_),
    .B(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__xor2_2 _19471_ (.A(_06515_),
    .B(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__a22o_2 _19472_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][10] ),
    .B1(_11712_),
    .B2(_06518_),
    .X(_01500_));
 sky130_fd_sc_hd__nor2_2 _19473_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[7][11] ),
    .Y(_06519_));
 sky130_fd_sc_hd__or2_2 _19474_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[7][11] ),
    .X(_06520_));
 sky130_fd_sc_hd__nand2_2 _19475_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[7][11] ),
    .Y(_06521_));
 sky130_fd_sc_hd__nand2_2 _19476_ (.A(_06520_),
    .B(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__a21bo_2 _19477_ (.A1(_06515_),
    .A2(_06517_),
    .B1_N(_06513_),
    .X(_06523_));
 sky130_fd_sc_hd__xnor2_2 _19478_ (.A(_06522_),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__a22o_2 _19479_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][11] ),
    .B1(_11712_),
    .B2(_06524_),
    .X(_01501_));
 sky130_fd_sc_hd__nand3_2 _19480_ (.A(_06515_),
    .B(_06520_),
    .C(_06521_),
    .Y(_06525_));
 sky130_fd_sc_hd__a211o_2 _19481_ (.A1(_06497_),
    .A2(_06500_),
    .B1(_06509_),
    .C1(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__o21a_2 _19482_ (.A1(_06513_),
    .A2(_06519_),
    .B1(_06521_),
    .X(_06527_));
 sky130_fd_sc_hd__o211a_2 _19483_ (.A1(_06516_),
    .A2(_06525_),
    .B1(_06526_),
    .C1(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__xnor2_2 _19484_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[7][12] ),
    .Y(_06529_));
 sky130_fd_sc_hd__inv_2 _19485_ (.A(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__nand2_2 _19486_ (.A(_06528_),
    .B(_06529_),
    .Y(_06531_));
 sky130_fd_sc_hd__nor2_2 _19487_ (.A(_06528_),
    .B(_06529_),
    .Y(_06532_));
 sky130_fd_sc_hd__nor2_2 _19488_ (.A(_11713_),
    .B(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__a22o_2 _19489_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][12] ),
    .B1(_06531_),
    .B2(_06533_),
    .X(_01502_));
 sky130_fd_sc_hd__xor2_2 _19490_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[7][13] ),
    .X(_06534_));
 sky130_fd_sc_hd__a211o_2 _19491_ (.A1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[7][12] ),
    .B1(_06532_),
    .C1(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__nand2_2 _19492_ (.A(_06530_),
    .B(_06534_),
    .Y(_06536_));
 sky130_fd_sc_hd__and3_2 _19493_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[7][12] ),
    .C(_06534_),
    .X(_06537_));
 sky130_fd_sc_hd__a21oi_2 _19494_ (.A1(_06532_),
    .A2(_06534_),
    .B1(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__a32o_2 _19495_ (.A1(_11712_),
    .A2(_06535_),
    .A3(_06538_),
    .B1(\systolic_inst.acc_wires[7][13] ),
    .B2(_11258_),
    .X(_01503_));
 sky130_fd_sc_hd__or2_2 _19496_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[7][14] ),
    .X(_06539_));
 sky130_fd_sc_hd__nand2_2 _19497_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[7][14] ),
    .Y(_06540_));
 sky130_fd_sc_hd__and2_2 _19498_ (.A(_06539_),
    .B(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__a21oi_2 _19499_ (.A1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[7][13] ),
    .B1(_06537_),
    .Y(_06542_));
 sky130_fd_sc_hd__o21ai_2 _19500_ (.A1(_06528_),
    .A2(_06536_),
    .B1(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__nand2_2 _19501_ (.A(_06541_),
    .B(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__or2_2 _19502_ (.A(_06541_),
    .B(_06543_),
    .X(_06545_));
 sky130_fd_sc_hd__a32o_2 _19503_ (.A1(_11712_),
    .A2(_06544_),
    .A3(_06545_),
    .B1(\systolic_inst.acc_wires[7][14] ),
    .B2(_11258_),
    .X(_01504_));
 sky130_fd_sc_hd__nor2_2 _19504_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][15] ),
    .Y(_06546_));
 sky130_fd_sc_hd__and2_2 _19505_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][15] ),
    .X(_06547_));
 sky130_fd_sc_hd__a211o_2 _19506_ (.A1(_06540_),
    .A2(_06544_),
    .B1(_06546_),
    .C1(_06547_),
    .X(_06548_));
 sky130_fd_sc_hd__o211ai_2 _19507_ (.A1(_06546_),
    .A2(_06547_),
    .B1(_06540_),
    .C1(_06544_),
    .Y(_06549_));
 sky130_fd_sc_hd__a32o_2 _19508_ (.A1(_11712_),
    .A2(_06548_),
    .A3(_06549_),
    .B1(\systolic_inst.acc_wires[7][15] ),
    .B2(_11258_),
    .X(_01505_));
 sky130_fd_sc_hd__or3b_2 _19509_ (.A(_06546_),
    .B(_06547_),
    .C_N(_06541_),
    .X(_06550_));
 sky130_fd_sc_hd__or2_2 _19510_ (.A(_06542_),
    .B(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__o31a_2 _19511_ (.A1(_06528_),
    .A2(_06536_),
    .A3(_06550_),
    .B1(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__o21ba_2 _19512_ (.A1(_06540_),
    .A2(_06546_),
    .B1_N(_06547_),
    .X(_06553_));
 sky130_fd_sc_hd__and2_2 _19513_ (.A(_06552_),
    .B(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__xnor2_2 _19514_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][16] ),
    .Y(_06555_));
 sky130_fd_sc_hd__nand2_2 _19515_ (.A(_06554_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__nor2_2 _19516_ (.A(_06554_),
    .B(_06555_),
    .Y(_06557_));
 sky130_fd_sc_hd__nor2_2 _19517_ (.A(_11713_),
    .B(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__a22o_2 _19518_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][16] ),
    .B1(_06556_),
    .B2(_06558_),
    .X(_01506_));
 sky130_fd_sc_hd__xor2_2 _19519_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][17] ),
    .X(_06559_));
 sky130_fd_sc_hd__inv_2 _19520_ (.A(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__a21oi_2 _19521_ (.A1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[7][16] ),
    .B1(_06557_),
    .Y(_06561_));
 sky130_fd_sc_hd__xnor2_2 _19522_ (.A(_06559_),
    .B(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__a22o_2 _19523_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][17] ),
    .B1(_11712_),
    .B2(_06562_),
    .X(_01507_));
 sky130_fd_sc_hd__or2_2 _19524_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][18] ),
    .X(_06563_));
 sky130_fd_sc_hd__nand2_2 _19525_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][18] ),
    .Y(_06564_));
 sky130_fd_sc_hd__nand2_2 _19526_ (.A(_06563_),
    .B(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__o21a_2 _19527_ (.A1(\systolic_inst.acc_wires[7][16] ),
    .A2(\systolic_inst.acc_wires[7][17] ),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .X(_06566_));
 sky130_fd_sc_hd__a21oi_2 _19528_ (.A1(_06557_),
    .A2(_06559_),
    .B1(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__xor2_2 _19529_ (.A(_06565_),
    .B(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__a22o_2 _19530_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][18] ),
    .B1(_11712_),
    .B2(_06568_),
    .X(_01508_));
 sky130_fd_sc_hd__xnor2_2 _19531_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][19] ),
    .Y(_06569_));
 sky130_fd_sc_hd__o21ai_2 _19532_ (.A1(_06565_),
    .A2(_06567_),
    .B1(_06564_),
    .Y(_06570_));
 sky130_fd_sc_hd__xnor2_2 _19533_ (.A(_06569_),
    .B(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__a22o_2 _19534_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][19] ),
    .B1(_11712_),
    .B2(_06571_),
    .X(_01509_));
 sky130_fd_sc_hd__or2_2 _19535_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][20] ),
    .X(_06572_));
 sky130_fd_sc_hd__nand2_2 _19536_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][20] ),
    .Y(_06573_));
 sky130_fd_sc_hd__and2_2 _19537_ (.A(_06572_),
    .B(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__or4_2 _19538_ (.A(_06555_),
    .B(_06560_),
    .C(_06565_),
    .D(_06569_),
    .X(_06575_));
 sky130_fd_sc_hd__nor2_2 _19539_ (.A(_06554_),
    .B(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__o41a_2 _19540_ (.A1(\systolic_inst.acc_wires[7][16] ),
    .A2(\systolic_inst.acc_wires[7][17] ),
    .A3(\systolic_inst.acc_wires[7][18] ),
    .A4(\systolic_inst.acc_wires[7][19] ),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .X(_06577_));
 sky130_fd_sc_hd__or3_2 _19541_ (.A(_06574_),
    .B(_06576_),
    .C(_06577_),
    .X(_06578_));
 sky130_fd_sc_hd__o21ai_2 _19542_ (.A1(_06576_),
    .A2(_06577_),
    .B1(_06574_),
    .Y(_06579_));
 sky130_fd_sc_hd__a32o_2 _19543_ (.A1(_11712_),
    .A2(_06578_),
    .A3(_06579_),
    .B1(\systolic_inst.acc_wires[7][20] ),
    .B2(_11258_),
    .X(_01510_));
 sky130_fd_sc_hd__xnor2_2 _19544_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][21] ),
    .Y(_06580_));
 sky130_fd_sc_hd__inv_2 _19545_ (.A(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__a21oi_2 _19546_ (.A1(_06573_),
    .A2(_06579_),
    .B1(_06580_),
    .Y(_06582_));
 sky130_fd_sc_hd__a31o_2 _19547_ (.A1(_06573_),
    .A2(_06579_),
    .A3(_06580_),
    .B1(_11713_),
    .X(_06583_));
 sky130_fd_sc_hd__a2bb2o_2 _19548_ (.A1_N(_06583_),
    .A2_N(_06582_),
    .B1(\systolic_inst.acc_wires[7][21] ),
    .B2(_11258_),
    .X(_01511_));
 sky130_fd_sc_hd__or2_2 _19549_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][22] ),
    .X(_06584_));
 sky130_fd_sc_hd__nand2_2 _19550_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][22] ),
    .Y(_06585_));
 sky130_fd_sc_hd__and2_2 _19551_ (.A(_06584_),
    .B(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__o21a_2 _19552_ (.A1(\systolic_inst.acc_wires[7][20] ),
    .A2(\systolic_inst.acc_wires[7][21] ),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .X(_06587_));
 sky130_fd_sc_hd__nor2_2 _19553_ (.A(_06579_),
    .B(_06580_),
    .Y(_06588_));
 sky130_fd_sc_hd__o21ai_2 _19554_ (.A1(_06587_),
    .A2(_06588_),
    .B1(_06586_),
    .Y(_06589_));
 sky130_fd_sc_hd__or3_2 _19555_ (.A(_06586_),
    .B(_06587_),
    .C(_06588_),
    .X(_06590_));
 sky130_fd_sc_hd__a32o_2 _19556_ (.A1(_11712_),
    .A2(_06589_),
    .A3(_06590_),
    .B1(\systolic_inst.acc_wires[7][22] ),
    .B2(_11258_),
    .X(_01512_));
 sky130_fd_sc_hd__xor2_2 _19557_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][23] ),
    .X(_06591_));
 sky130_fd_sc_hd__inv_2 _19558_ (.A(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__nand3_2 _19559_ (.A(_06585_),
    .B(_06589_),
    .C(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__a21o_2 _19560_ (.A1(_06585_),
    .A2(_06589_),
    .B1(_06592_),
    .X(_06594_));
 sky130_fd_sc_hd__a32o_2 _19561_ (.A1(_11712_),
    .A2(_06593_),
    .A3(_06594_),
    .B1(\systolic_inst.acc_wires[7][23] ),
    .B2(_11258_),
    .X(_01513_));
 sky130_fd_sc_hd__nand4_2 _19562_ (.A(_06574_),
    .B(_06581_),
    .C(_06586_),
    .D(_06591_),
    .Y(_06595_));
 sky130_fd_sc_hd__a211o_2 _19563_ (.A1(_06552_),
    .A2(_06553_),
    .B1(_06575_),
    .C1(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__o41a_2 _19564_ (.A1(\systolic_inst.acc_wires[7][20] ),
    .A2(\systolic_inst.acc_wires[7][21] ),
    .A3(\systolic_inst.acc_wires[7][22] ),
    .A4(\systolic_inst.acc_wires[7][23] ),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .X(_06597_));
 sky130_fd_sc_hd__nor2_2 _19565_ (.A(_06577_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__nor2_2 _19566_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][24] ),
    .Y(_06599_));
 sky130_fd_sc_hd__and2_2 _19567_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][24] ),
    .X(_06600_));
 sky130_fd_sc_hd__or2_2 _19568_ (.A(_06599_),
    .B(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__a21oi_2 _19569_ (.A1(_06596_),
    .A2(_06598_),
    .B1(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__a31o_2 _19570_ (.A1(_06596_),
    .A2(_06598_),
    .A3(_06601_),
    .B1(_11713_),
    .X(_06603_));
 sky130_fd_sc_hd__a2bb2o_2 _19571_ (.A1_N(_06603_),
    .A2_N(_06602_),
    .B1(\systolic_inst.acc_wires[7][24] ),
    .B2(_11258_),
    .X(_01514_));
 sky130_fd_sc_hd__xor2_2 _19572_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][25] ),
    .X(_06604_));
 sky130_fd_sc_hd__or3_2 _19573_ (.A(_06600_),
    .B(_06602_),
    .C(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__o21ai_2 _19574_ (.A1(_06600_),
    .A2(_06602_),
    .B1(_06604_),
    .Y(_06606_));
 sky130_fd_sc_hd__a32o_2 _19575_ (.A1(_11712_),
    .A2(_06605_),
    .A3(_06606_),
    .B1(\systolic_inst.acc_wires[7][25] ),
    .B2(_11258_),
    .X(_01515_));
 sky130_fd_sc_hd__or2_2 _19576_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][26] ),
    .X(_06607_));
 sky130_fd_sc_hd__nand2_2 _19577_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][26] ),
    .Y(_06608_));
 sky130_fd_sc_hd__nand2_2 _19578_ (.A(_06607_),
    .B(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__o21a_2 _19579_ (.A1(\systolic_inst.acc_wires[7][24] ),
    .A2(\systolic_inst.acc_wires[7][25] ),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .X(_06610_));
 sky130_fd_sc_hd__a21o_2 _19580_ (.A1(_06602_),
    .A2(_06604_),
    .B1(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__xnor2_2 _19581_ (.A(_06609_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__a22o_2 _19582_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][26] ),
    .B1(_11712_),
    .B2(_06612_),
    .X(_01516_));
 sky130_fd_sc_hd__xnor2_2 _19583_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][27] ),
    .Y(_06613_));
 sky130_fd_sc_hd__a21bo_2 _19584_ (.A1(_06607_),
    .A2(_06611_),
    .B1_N(_06608_),
    .X(_06614_));
 sky130_fd_sc_hd__xnor2_2 _19585_ (.A(_06613_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__a22o_2 _19586_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][27] ),
    .B1(_11712_),
    .B2(_06615_),
    .X(_01517_));
 sky130_fd_sc_hd__nor2_2 _19587_ (.A(_06609_),
    .B(_06613_),
    .Y(_06616_));
 sky130_fd_sc_hd__o21a_2 _19588_ (.A1(\systolic_inst.acc_wires[7][26] ),
    .A2(\systolic_inst.acc_wires[7][27] ),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .X(_06617_));
 sky130_fd_sc_hd__a311oi_2 _19589_ (.A1(_06602_),
    .A2(_06604_),
    .A3(_06616_),
    .B1(_06617_),
    .C1(_06610_),
    .Y(_06618_));
 sky130_fd_sc_hd__or2_2 _19590_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][28] ),
    .X(_06619_));
 sky130_fd_sc_hd__nand2_2 _19591_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][28] ),
    .Y(_06620_));
 sky130_fd_sc_hd__nand2_2 _19592_ (.A(_06619_),
    .B(_06620_),
    .Y(_06621_));
 sky130_fd_sc_hd__xor2_2 _19593_ (.A(_06618_),
    .B(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__a22o_2 _19594_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][28] ),
    .B1(_11712_),
    .B2(_06622_),
    .X(_01518_));
 sky130_fd_sc_hd__xor2_2 _19595_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][29] ),
    .X(_06623_));
 sky130_fd_sc_hd__inv_2 _19596_ (.A(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__o21a_2 _19597_ (.A1(_06618_),
    .A2(_06621_),
    .B1(_06620_),
    .X(_06625_));
 sky130_fd_sc_hd__xnor2_2 _19598_ (.A(_06623_),
    .B(_06625_),
    .Y(_06626_));
 sky130_fd_sc_hd__a22o_2 _19599_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[7][29] ),
    .B1(_11712_),
    .B2(_06626_),
    .X(_01519_));
 sky130_fd_sc_hd__o21ai_2 _19600_ (.A1(\systolic_inst.acc_wires[7][28] ),
    .A2(\systolic_inst.acc_wires[7][29] ),
    .B1(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .Y(_06627_));
 sky130_fd_sc_hd__o31a_2 _19601_ (.A1(_06618_),
    .A2(_06621_),
    .A3(_06624_),
    .B1(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__nand2_2 _19602_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][30] ),
    .Y(_06629_));
 sky130_fd_sc_hd__or2_2 _19603_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][30] ),
    .X(_06630_));
 sky130_fd_sc_hd__nand2_2 _19604_ (.A(_06629_),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_2 _19605_ (.A(_06628_),
    .B(_06631_),
    .Y(_06632_));
 sky130_fd_sc_hd__or2_2 _19606_ (.A(_06628_),
    .B(_06631_),
    .X(_06633_));
 sky130_fd_sc_hd__a32o_2 _19607_ (.A1(_11712_),
    .A2(_06632_),
    .A3(_06633_),
    .B1(\systolic_inst.acc_wires[7][30] ),
    .B2(_11258_),
    .X(_01520_));
 sky130_fd_sc_hd__xnor2_2 _19608_ (.A(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[7][31] ),
    .Y(_06634_));
 sky130_fd_sc_hd__a21oi_2 _19609_ (.A1(_06629_),
    .A2(_06633_),
    .B1(_06634_),
    .Y(_06635_));
 sky130_fd_sc_hd__a31o_2 _19610_ (.A1(_06629_),
    .A2(_06633_),
    .A3(_06634_),
    .B1(_11713_),
    .X(_06636_));
 sky130_fd_sc_hd__a2bb2o_2 _19611_ (.A1_N(_06636_),
    .A2_N(_06635_),
    .B1(\systolic_inst.acc_wires[7][31] ),
    .B2(_11258_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _19612_ (.A0(\systolic_inst.A_outs[6][0] ),
    .A1(\systolic_inst.A_outs[5][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _19613_ (.A0(\systolic_inst.A_outs[6][1] ),
    .A1(\systolic_inst.A_outs[5][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _19614_ (.A0(\systolic_inst.A_outs[6][2] ),
    .A1(\systolic_inst.A_outs[5][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _19615_ (.A0(\systolic_inst.A_outs[6][3] ),
    .A1(\systolic_inst.A_outs[5][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _19616_ (.A0(\systolic_inst.A_outs[6][4] ),
    .A1(\systolic_inst.A_outs[5][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _19617_ (.A0(\systolic_inst.A_outs[6][5] ),
    .A1(\systolic_inst.A_outs[5][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _19618_ (.A0(\systolic_inst.A_outs[6][6] ),
    .A1(\systolic_inst.A_outs[5][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _19619_ (.A0(\systolic_inst.A_outs[6][7] ),
    .A1(\systolic_inst.A_outs[5][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _19620_ (.A0(\systolic_inst.B_outs[5][0] ),
    .A1(\systolic_inst.B_outs[1][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _19621_ (.A0(\systolic_inst.B_outs[5][1] ),
    .A1(\systolic_inst.B_outs[1][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _19622_ (.A0(\systolic_inst.B_outs[5][2] ),
    .A1(\systolic_inst.B_outs[1][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _19623_ (.A0(\systolic_inst.B_outs[5][3] ),
    .A1(\systolic_inst.B_outs[1][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _19624_ (.A0(\systolic_inst.B_outs[5][4] ),
    .A1(\systolic_inst.B_outs[1][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _19625_ (.A0(\systolic_inst.B_outs[5][5] ),
    .A1(\systolic_inst.B_outs[1][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _19626_ (.A0(\systolic_inst.B_outs[5][6] ),
    .A1(\systolic_inst.B_outs[1][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _19627_ (.A0(\systolic_inst.B_outs[5][7] ),
    .A1(\systolic_inst.B_outs[1][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01537_));
 sky130_fd_sc_hd__and3_2 _19628_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[6][0] ),
    .C(\systolic_inst.A_outs[6][0] ),
    .X(_06637_));
 sky130_fd_sc_hd__a21o_2 _19629_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[0] ),
    .B1(_06637_),
    .X(_01538_));
 sky130_fd_sc_hd__and4_2 _19630_ (.A(\systolic_inst.B_outs[6][0] ),
    .B(\systolic_inst.A_outs[6][0] ),
    .C(\systolic_inst.B_outs[6][1] ),
    .D(\systolic_inst.A_outs[6][1] ),
    .X(_06638_));
 sky130_fd_sc_hd__a22o_2 _19631_ (.A1(\systolic_inst.A_outs[6][0] ),
    .A2(\systolic_inst.B_outs[6][1] ),
    .B1(\systolic_inst.A_outs[6][1] ),
    .B2(\systolic_inst.B_outs[6][0] ),
    .X(_06639_));
 sky130_fd_sc_hd__nand2_2 _19632_ (.A(\systolic_inst.ce_local ),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__a2bb2o_2 _19633_ (.A1_N(_06640_),
    .A2_N(_06638_),
    .B1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01539_));
 sky130_fd_sc_hd__nand2_2 _19634_ (.A(\systolic_inst.B_outs[6][1] ),
    .B(\systolic_inst.A_outs[6][1] ),
    .Y(_06641_));
 sky130_fd_sc_hd__nand2_2 _19635_ (.A(\systolic_inst.B_outs[6][0] ),
    .B(\systolic_inst.A_outs[6][2] ),
    .Y(_06642_));
 sky130_fd_sc_hd__and4_2 _19636_ (.A(\systolic_inst.B_outs[6][0] ),
    .B(\systolic_inst.B_outs[6][1] ),
    .C(\systolic_inst.A_outs[6][1] ),
    .D(\systolic_inst.A_outs[6][2] ),
    .X(_06643_));
 sky130_fd_sc_hd__a21o_2 _19637_ (.A1(_06641_),
    .A2(_06642_),
    .B1(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__inv_2 _19638_ (.A(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__xnor2_2 _19639_ (.A(_06638_),
    .B(_06644_),
    .Y(_06646_));
 sky130_fd_sc_hd__nand3_2 _19640_ (.A(\systolic_inst.A_outs[6][0] ),
    .B(\systolic_inst.B_outs[6][2] ),
    .C(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__a21o_2 _19641_ (.A1(\systolic_inst.A_outs[6][0] ),
    .A2(\systolic_inst.B_outs[6][2] ),
    .B1(_06646_),
    .X(_06648_));
 sky130_fd_sc_hd__and2_2 _19642_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[2] ),
    .X(_06649_));
 sky130_fd_sc_hd__a31o_2 _19643_ (.A1(\systolic_inst.ce_local ),
    .A2(_06647_),
    .A3(_06648_),
    .B1(_06649_),
    .X(_01540_));
 sky130_fd_sc_hd__a22oi_2 _19644_ (.A1(\systolic_inst.A_outs[6][1] ),
    .A2(\systolic_inst.B_outs[6][2] ),
    .B1(\systolic_inst.B_outs[6][3] ),
    .B2(\systolic_inst.A_outs[6][0] ),
    .Y(_06650_));
 sky130_fd_sc_hd__and4_2 _19645_ (.A(\systolic_inst.A_outs[6][0] ),
    .B(\systolic_inst.A_outs[6][1] ),
    .C(\systolic_inst.B_outs[6][2] ),
    .D(\systolic_inst.B_outs[6][3] ),
    .X(_06651_));
 sky130_fd_sc_hd__or2_2 _19646_ (.A(_06650_),
    .B(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__nand2_2 _19647_ (.A(\systolic_inst.B_outs[6][1] ),
    .B(\systolic_inst.A_outs[6][3] ),
    .Y(_06653_));
 sky130_fd_sc_hd__or2_2 _19648_ (.A(_06642_),
    .B(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__a22o_2 _19649_ (.A1(\systolic_inst.B_outs[6][1] ),
    .A2(\systolic_inst.A_outs[6][2] ),
    .B1(\systolic_inst.A_outs[6][3] ),
    .B2(\systolic_inst.B_outs[6][0] ),
    .X(_06655_));
 sky130_fd_sc_hd__nand3_2 _19650_ (.A(_06643_),
    .B(_06654_),
    .C(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__a21o_2 _19651_ (.A1(_06654_),
    .A2(_06655_),
    .B1(_06643_),
    .X(_06657_));
 sky130_fd_sc_hd__nand2_2 _19652_ (.A(_06656_),
    .B(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__xnor2_2 _19653_ (.A(_06652_),
    .B(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__a21bo_2 _19654_ (.A1(_06638_),
    .A2(_06645_),
    .B1_N(_06647_),
    .X(_06660_));
 sky130_fd_sc_hd__and2b_2 _19655_ (.A_N(_06659_),
    .B(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__xnor2_2 _19656_ (.A(_06659_),
    .B(_06660_),
    .Y(_06662_));
 sky130_fd_sc_hd__mux2_1 _19657_ (.A0(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[3] ),
    .A1(_06662_),
    .S(\systolic_inst.ce_local ),
    .X(_01541_));
 sky130_fd_sc_hd__and2_2 _19658_ (.A(\systolic_inst.B_outs[6][2] ),
    .B(\systolic_inst.A_outs[6][2] ),
    .X(_06663_));
 sky130_fd_sc_hd__nand4_2 _19659_ (.A(\systolic_inst.A_outs[6][0] ),
    .B(\systolic_inst.A_outs[6][1] ),
    .C(\systolic_inst.B_outs[6][3] ),
    .D(\systolic_inst.B_outs[6][4] ),
    .Y(_06664_));
 sky130_fd_sc_hd__a22o_2 _19660_ (.A1(\systolic_inst.A_outs[6][1] ),
    .A2(\systolic_inst.B_outs[6][3] ),
    .B1(\systolic_inst.B_outs[6][4] ),
    .B2(\systolic_inst.A_outs[6][0] ),
    .X(_06665_));
 sky130_fd_sc_hd__nand2_2 _19661_ (.A(_06664_),
    .B(_06665_),
    .Y(_06666_));
 sky130_fd_sc_hd__xnor2_2 _19662_ (.A(_06663_),
    .B(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__inv_2 _19663_ (.A(_06667_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_2 _19664_ (.A(\systolic_inst.B_outs[6][0] ),
    .B(\systolic_inst.A_outs[6][4] ),
    .Y(_06669_));
 sky130_fd_sc_hd__and4_2 _19665_ (.A(\systolic_inst.B_outs[6][0] ),
    .B(\systolic_inst.B_outs[6][1] ),
    .C(\systolic_inst.A_outs[6][3] ),
    .D(\systolic_inst.A_outs[6][4] ),
    .X(_06670_));
 sky130_fd_sc_hd__a21oi_2 _19666_ (.A1(_06653_),
    .A2(_06669_),
    .B1(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__xnor2_2 _19667_ (.A(_06651_),
    .B(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__nor2_2 _19668_ (.A(_06654_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__xnor2_2 _19669_ (.A(_06654_),
    .B(_06672_),
    .Y(_06674_));
 sky130_fd_sc_hd__nor2_2 _19670_ (.A(_06668_),
    .B(_06674_),
    .Y(_06675_));
 sky130_fd_sc_hd__and2_2 _19671_ (.A(_06668_),
    .B(_06674_),
    .X(_06676_));
 sky130_fd_sc_hd__or2_2 _19672_ (.A(_06675_),
    .B(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__o21ai_2 _19673_ (.A1(_06652_),
    .A2(_06658_),
    .B1(_06656_),
    .Y(_06678_));
 sky130_fd_sc_hd__nand2b_2 _19674_ (.A_N(_06677_),
    .B(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__xnor2_2 _19675_ (.A(_06677_),
    .B(_06678_),
    .Y(_06680_));
 sky130_fd_sc_hd__or2_2 _19676_ (.A(_06661_),
    .B(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__nand2_2 _19677_ (.A(_06661_),
    .B(_06680_),
    .Y(_06682_));
 sky130_fd_sc_hd__and2_2 _19678_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[4] ),
    .X(_06683_));
 sky130_fd_sc_hd__a31o_2 _19679_ (.A1(\systolic_inst.ce_local ),
    .A2(_06681_),
    .A3(_06682_),
    .B1(_06683_),
    .X(_01542_));
 sky130_fd_sc_hd__a21oi_2 _19680_ (.A1(_06651_),
    .A2(_06671_),
    .B1(_06673_),
    .Y(_06684_));
 sky130_fd_sc_hd__a21bo_2 _19681_ (.A1(_06663_),
    .A2(_06665_),
    .B1_N(_06664_),
    .X(_06685_));
 sky130_fd_sc_hd__a22oi_2 _19682_ (.A1(\systolic_inst.B_outs[6][1] ),
    .A2(\systolic_inst.A_outs[6][4] ),
    .B1(\systolic_inst.A_outs[6][5] ),
    .B2(\systolic_inst.B_outs[6][0] ),
    .Y(_06686_));
 sky130_fd_sc_hd__and4_2 _19683_ (.A(\systolic_inst.B_outs[6][0] ),
    .B(\systolic_inst.B_outs[6][1] ),
    .C(\systolic_inst.A_outs[6][4] ),
    .D(\systolic_inst.A_outs[6][5] ),
    .X(_06687_));
 sky130_fd_sc_hd__or2_2 _19684_ (.A(_06686_),
    .B(_06687_),
    .X(_06688_));
 sky130_fd_sc_hd__nand2b_2 _19685_ (.A_N(_06688_),
    .B(_06685_),
    .Y(_06689_));
 sky130_fd_sc_hd__xnor2_2 _19686_ (.A(_06685_),
    .B(_06688_),
    .Y(_06690_));
 sky130_fd_sc_hd__nand2_2 _19687_ (.A(_06670_),
    .B(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__xnor2_2 _19688_ (.A(_06670_),
    .B(_06690_),
    .Y(_06692_));
 sky130_fd_sc_hd__nand2_2 _19689_ (.A(\systolic_inst.A_outs[6][0] ),
    .B(\systolic_inst.B_outs[6][5] ),
    .Y(_06693_));
 sky130_fd_sc_hd__nand2_2 _19690_ (.A(\systolic_inst.B_outs[6][2] ),
    .B(\systolic_inst.A_outs[6][3] ),
    .Y(_06694_));
 sky130_fd_sc_hd__and4_2 _19691_ (.A(\systolic_inst.A_outs[6][1] ),
    .B(\systolic_inst.A_outs[6][2] ),
    .C(\systolic_inst.B_outs[6][3] ),
    .D(\systolic_inst.B_outs[6][4] ),
    .X(_06695_));
 sky130_fd_sc_hd__a22o_2 _19692_ (.A1(\systolic_inst.A_outs[6][2] ),
    .A2(\systolic_inst.B_outs[6][3] ),
    .B1(\systolic_inst.B_outs[6][4] ),
    .B2(\systolic_inst.A_outs[6][1] ),
    .X(_06696_));
 sky130_fd_sc_hd__and2b_2 _19693_ (.A_N(_06695_),
    .B(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__xnor2_2 _19694_ (.A(_06694_),
    .B(_06697_),
    .Y(_06698_));
 sky130_fd_sc_hd__nand2b_2 _19695_ (.A_N(_06693_),
    .B(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__xor2_2 _19696_ (.A(_06693_),
    .B(_06698_),
    .X(_06700_));
 sky130_fd_sc_hd__nor2_2 _19697_ (.A(_06692_),
    .B(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__inv_2 _19698_ (.A(_06701_),
    .Y(_06702_));
 sky130_fd_sc_hd__xor2_2 _19699_ (.A(_06692_),
    .B(_06700_),
    .X(_06703_));
 sky130_fd_sc_hd__nand2_2 _19700_ (.A(_06675_),
    .B(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__or2_2 _19701_ (.A(_06675_),
    .B(_06703_),
    .X(_06705_));
 sky130_fd_sc_hd__and2_2 _19702_ (.A(_06704_),
    .B(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__nand2b_2 _19703_ (.A_N(_06684_),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__xnor2_2 _19704_ (.A(_06684_),
    .B(_06706_),
    .Y(_06708_));
 sky130_fd_sc_hd__a21bo_2 _19705_ (.A1(_06661_),
    .A2(_06680_),
    .B1_N(_06679_),
    .X(_06709_));
 sky130_fd_sc_hd__nand2_2 _19706_ (.A(_06708_),
    .B(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__o21a_2 _19707_ (.A1(_06708_),
    .A2(_06709_),
    .B1(\systolic_inst.ce_local ),
    .X(_06711_));
 sky130_fd_sc_hd__a22o_2 _19708_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[5] ),
    .B1(_06710_),
    .B2(_06711_),
    .X(_01543_));
 sky130_fd_sc_hd__a31o_2 _19709_ (.A1(\systolic_inst.B_outs[6][2] ),
    .A2(\systolic_inst.A_outs[6][3] ),
    .A3(_06696_),
    .B1(_06695_),
    .X(_06712_));
 sky130_fd_sc_hd__a22oi_2 _19710_ (.A1(\systolic_inst.B_outs[6][1] ),
    .A2(\systolic_inst.A_outs[6][5] ),
    .B1(\systolic_inst.A_outs[6][6] ),
    .B2(\systolic_inst.B_outs[6][0] ),
    .Y(_06713_));
 sky130_fd_sc_hd__and4_2 _19711_ (.A(\systolic_inst.B_outs[6][0] ),
    .B(\systolic_inst.B_outs[6][1] ),
    .C(\systolic_inst.A_outs[6][5] ),
    .D(\systolic_inst.A_outs[6][6] ),
    .X(_06714_));
 sky130_fd_sc_hd__nor2_2 _19712_ (.A(_06713_),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__xor2_2 _19713_ (.A(_06712_),
    .B(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__and2_2 _19714_ (.A(_06687_),
    .B(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__nor2_2 _19715_ (.A(_06687_),
    .B(_06716_),
    .Y(_06718_));
 sky130_fd_sc_hd__or2_2 _19716_ (.A(_06717_),
    .B(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__nand2_2 _19717_ (.A(\systolic_inst.B_outs[6][2] ),
    .B(\systolic_inst.A_outs[6][4] ),
    .Y(_06720_));
 sky130_fd_sc_hd__and4_2 _19718_ (.A(\systolic_inst.A_outs[6][2] ),
    .B(\systolic_inst.B_outs[6][3] ),
    .C(\systolic_inst.A_outs[6][3] ),
    .D(\systolic_inst.B_outs[6][4] ),
    .X(_06721_));
 sky130_fd_sc_hd__a22oi_2 _19719_ (.A1(\systolic_inst.B_outs[6][3] ),
    .A2(\systolic_inst.A_outs[6][3] ),
    .B1(\systolic_inst.B_outs[6][4] ),
    .B2(\systolic_inst.A_outs[6][2] ),
    .Y(_06722_));
 sky130_fd_sc_hd__or2_2 _19720_ (.A(_06721_),
    .B(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__xnor2_2 _19721_ (.A(_06720_),
    .B(_06723_),
    .Y(_06724_));
 sky130_fd_sc_hd__a22oi_2 _19722_ (.A1(\systolic_inst.A_outs[6][1] ),
    .A2(\systolic_inst.B_outs[6][5] ),
    .B1(\systolic_inst.B_outs[6][6] ),
    .B2(\systolic_inst.A_outs[6][0] ),
    .Y(_06725_));
 sky130_fd_sc_hd__nand2_2 _19723_ (.A(\systolic_inst.A_outs[6][1] ),
    .B(\systolic_inst.B_outs[6][6] ),
    .Y(_06726_));
 sky130_fd_sc_hd__nor2_2 _19724_ (.A(_06693_),
    .B(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__nor2_2 _19725_ (.A(_06725_),
    .B(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__or3_2 _19726_ (.A(_06724_),
    .B(_06725_),
    .C(_06727_),
    .X(_06729_));
 sky130_fd_sc_hd__xor2_2 _19727_ (.A(_06724_),
    .B(_06728_),
    .X(_06730_));
 sky130_fd_sc_hd__xnor2_2 _19728_ (.A(_06699_),
    .B(_06730_),
    .Y(_06731_));
 sky130_fd_sc_hd__xnor2_2 _19729_ (.A(_06719_),
    .B(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__xnor2_2 _19730_ (.A(_06702_),
    .B(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__a21oi_2 _19731_ (.A1(_06689_),
    .A2(_06691_),
    .B1(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__and3_2 _19732_ (.A(_06689_),
    .B(_06691_),
    .C(_06733_),
    .X(_06735_));
 sky130_fd_sc_hd__a211oi_2 _19733_ (.A1(_06704_),
    .A2(_06707_),
    .B1(_06734_),
    .C1(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__o211a_2 _19734_ (.A1(_06734_),
    .A2(_06735_),
    .B1(_06704_),
    .C1(_06707_),
    .X(_06737_));
 sky130_fd_sc_hd__o21ai_2 _19735_ (.A1(_06736_),
    .A2(_06737_),
    .B1(_06710_),
    .Y(_06738_));
 sky130_fd_sc_hd__nor3_2 _19736_ (.A(_06710_),
    .B(_06736_),
    .C(_06737_),
    .Y(_06739_));
 sky130_fd_sc_hd__nor2_2 _19737_ (.A(_11258_),
    .B(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__a22o_2 _19738_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[6] ),
    .B1(_06738_),
    .B2(_06740_),
    .X(_01544_));
 sky130_fd_sc_hd__o21ba_2 _19739_ (.A1(_06702_),
    .A2(_06732_),
    .B1_N(_06734_),
    .X(_06741_));
 sky130_fd_sc_hd__a21oi_2 _19740_ (.A1(_06712_),
    .A2(_06715_),
    .B1(_06717_),
    .Y(_06742_));
 sky130_fd_sc_hd__o21ba_2 _19741_ (.A1(_06720_),
    .A2(_06722_),
    .B1_N(_06721_),
    .X(_06743_));
 sky130_fd_sc_hd__a22o_2 _19742_ (.A1(\systolic_inst.B_outs[6][1] ),
    .A2(\systolic_inst.A_outs[6][6] ),
    .B1(\systolic_inst.A_outs[6][7] ),
    .B2(\systolic_inst.B_outs[6][0] ),
    .X(_06744_));
 sky130_fd_sc_hd__nand4_2 _19743_ (.A(\systolic_inst.B_outs[6][0] ),
    .B(\systolic_inst.B_outs[6][1] ),
    .C(\systolic_inst.A_outs[6][6] ),
    .D(\systolic_inst.A_outs[6][7] ),
    .Y(_06745_));
 sky130_fd_sc_hd__nand2_2 _19744_ (.A(_06744_),
    .B(_06745_),
    .Y(_06746_));
 sky130_fd_sc_hd__xnor2_2 _19745_ (.A(_11278_),
    .B(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__nor2_2 _19746_ (.A(_06743_),
    .B(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__and2_2 _19747_ (.A(_06743_),
    .B(_06747_),
    .X(_06749_));
 sky130_fd_sc_hd__nor2_2 _19748_ (.A(_06748_),
    .B(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__xnor2_2 _19749_ (.A(_06714_),
    .B(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__nand2_2 _19750_ (.A(\systolic_inst.B_outs[6][2] ),
    .B(\systolic_inst.A_outs[6][5] ),
    .Y(_06752_));
 sky130_fd_sc_hd__and4_2 _19751_ (.A(\systolic_inst.B_outs[6][3] ),
    .B(\systolic_inst.A_outs[6][3] ),
    .C(\systolic_inst.B_outs[6][4] ),
    .D(\systolic_inst.A_outs[6][4] ),
    .X(_06753_));
 sky130_fd_sc_hd__a22oi_2 _19752_ (.A1(\systolic_inst.A_outs[6][3] ),
    .A2(\systolic_inst.B_outs[6][4] ),
    .B1(\systolic_inst.A_outs[6][4] ),
    .B2(\systolic_inst.B_outs[6][3] ),
    .Y(_06754_));
 sky130_fd_sc_hd__or2_2 _19753_ (.A(_06753_),
    .B(_06754_),
    .X(_06755_));
 sky130_fd_sc_hd__xnor2_2 _19754_ (.A(_06752_),
    .B(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__nand2_2 _19755_ (.A(\systolic_inst.A_outs[6][2] ),
    .B(\systolic_inst.B_outs[6][5] ),
    .Y(_06757_));
 sky130_fd_sc_hd__and2b_2 _19756_ (.A_N(\systolic_inst.A_outs[6][0] ),
    .B(\systolic_inst.B_outs[6][7] ),
    .X(_06758_));
 sky130_fd_sc_hd__and3_2 _19757_ (.A(\systolic_inst.A_outs[6][1] ),
    .B(\systolic_inst.B_outs[6][6] ),
    .C(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__xnor2_2 _19758_ (.A(_06726_),
    .B(_06758_),
    .Y(_06760_));
 sky130_fd_sc_hd__xnor2_2 _19759_ (.A(_06757_),
    .B(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__xnor2_2 _19760_ (.A(_06727_),
    .B(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__nor2_2 _19761_ (.A(_06756_),
    .B(_06762_),
    .Y(_06763_));
 sky130_fd_sc_hd__xnor2_2 _19762_ (.A(_06756_),
    .B(_06762_),
    .Y(_06764_));
 sky130_fd_sc_hd__or2_2 _19763_ (.A(_06729_),
    .B(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__and2_2 _19764_ (.A(_06729_),
    .B(_06764_),
    .X(_06766_));
 sky130_fd_sc_hd__xor2_2 _19765_ (.A(_06729_),
    .B(_06764_),
    .X(_06767_));
 sky130_fd_sc_hd__xnor2_2 _19766_ (.A(_06751_),
    .B(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__o32a_2 _19767_ (.A1(_06717_),
    .A2(_06718_),
    .A3(_06731_),
    .B1(_06730_),
    .B2(_06699_),
    .X(_06769_));
 sky130_fd_sc_hd__nand2b_2 _19768_ (.A_N(_06769_),
    .B(_06768_),
    .Y(_06770_));
 sky130_fd_sc_hd__xnor2_2 _19769_ (.A(_06768_),
    .B(_06769_),
    .Y(_06771_));
 sky130_fd_sc_hd__nand2b_2 _19770_ (.A_N(_06742_),
    .B(_06771_),
    .Y(_06772_));
 sky130_fd_sc_hd__xnor2_2 _19771_ (.A(_06742_),
    .B(_06771_),
    .Y(_06773_));
 sky130_fd_sc_hd__and2b_2 _19772_ (.A_N(_06741_),
    .B(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__xnor2_2 _19773_ (.A(_06741_),
    .B(_06773_),
    .Y(_06775_));
 sky130_fd_sc_hd__nor3_2 _19774_ (.A(_06736_),
    .B(_06739_),
    .C(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__o21a_2 _19775_ (.A1(_06736_),
    .A2(_06739_),
    .B1(_06775_),
    .X(_06777_));
 sky130_fd_sc_hd__nand2_2 _19776_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[7] ),
    .Y(_06778_));
 sky130_fd_sc_hd__o31ai_2 _19777_ (.A1(_11258_),
    .A2(_06776_),
    .A3(_06777_),
    .B1(_06778_),
    .Y(_01545_));
 sky130_fd_sc_hd__a21o_2 _19778_ (.A1(_06714_),
    .A2(_06750_),
    .B1(_06748_),
    .X(_06779_));
 sky130_fd_sc_hd__a21bo_2 _19779_ (.A1(\systolic_inst.B_outs[6][7] ),
    .A2(_06744_),
    .B1_N(_06745_),
    .X(_06780_));
 sky130_fd_sc_hd__o21bai_2 _19780_ (.A1(_06752_),
    .A2(_06754_),
    .B1_N(_06753_),
    .Y(_06781_));
 sky130_fd_sc_hd__o21a_2 _19781_ (.A1(\systolic_inst.B_outs[6][0] ),
    .A2(\systolic_inst.B_outs[6][1] ),
    .B1(\systolic_inst.A_outs[6][7] ),
    .X(_06782_));
 sky130_fd_sc_hd__o21ai_2 _19782_ (.A1(\systolic_inst.B_outs[6][0] ),
    .A2(\systolic_inst.B_outs[6][1] ),
    .B1(\systolic_inst.A_outs[6][7] ),
    .Y(_06783_));
 sky130_fd_sc_hd__a21o_2 _19783_ (.A1(\systolic_inst.B_outs[6][0] ),
    .A2(\systolic_inst.B_outs[6][1] ),
    .B1(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__and2b_2 _19784_ (.A_N(_06784_),
    .B(_06781_),
    .X(_06785_));
 sky130_fd_sc_hd__xnor2_2 _19785_ (.A(_06781_),
    .B(_06784_),
    .Y(_06786_));
 sky130_fd_sc_hd__xnor2_2 _19786_ (.A(_06780_),
    .B(_06786_),
    .Y(_06787_));
 sky130_fd_sc_hd__and4_2 _19787_ (.A(\systolic_inst.B_outs[6][3] ),
    .B(\systolic_inst.B_outs[6][4] ),
    .C(\systolic_inst.A_outs[6][4] ),
    .D(\systolic_inst.A_outs[6][5] ),
    .X(_06788_));
 sky130_fd_sc_hd__a22oi_2 _19788_ (.A1(\systolic_inst.B_outs[6][4] ),
    .A2(\systolic_inst.A_outs[6][4] ),
    .B1(\systolic_inst.A_outs[6][5] ),
    .B2(\systolic_inst.B_outs[6][3] ),
    .Y(_06789_));
 sky130_fd_sc_hd__nor2_2 _19789_ (.A(_06788_),
    .B(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__nand2_2 _19790_ (.A(\systolic_inst.B_outs[6][2] ),
    .B(\systolic_inst.A_outs[6][6] ),
    .Y(_06791_));
 sky130_fd_sc_hd__xnor2_2 _19791_ (.A(_06790_),
    .B(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__nand2_2 _19792_ (.A(\systolic_inst.A_outs[6][3] ),
    .B(\systolic_inst.B_outs[6][5] ),
    .Y(_06793_));
 sky130_fd_sc_hd__and4b_2 _19793_ (.A_N(\systolic_inst.A_outs[6][1] ),
    .B(\systolic_inst.A_outs[6][2] ),
    .C(\systolic_inst.B_outs[6][6] ),
    .D(\systolic_inst.B_outs[6][7] ),
    .X(_06794_));
 sky130_fd_sc_hd__o2bb2a_2 _19794_ (.A1_N(\systolic_inst.A_outs[6][2] ),
    .A2_N(\systolic_inst.B_outs[6][6] ),
    .B1(_11278_),
    .B2(\systolic_inst.A_outs[6][1] ),
    .X(_06795_));
 sky130_fd_sc_hd__nor2_2 _19795_ (.A(_06794_),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__xnor2_2 _19796_ (.A(_06793_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__a31oi_2 _19797_ (.A1(\systolic_inst.A_outs[6][2] ),
    .A2(\systolic_inst.B_outs[6][5] ),
    .A3(_06760_),
    .B1(_06759_),
    .Y(_06798_));
 sky130_fd_sc_hd__nand2b_2 _19798_ (.A_N(_06798_),
    .B(_06797_),
    .Y(_06799_));
 sky130_fd_sc_hd__xnor2_2 _19799_ (.A(_06797_),
    .B(_06798_),
    .Y(_06800_));
 sky130_fd_sc_hd__nand2_2 _19800_ (.A(_06792_),
    .B(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__xnor2_2 _19801_ (.A(_06792_),
    .B(_06800_),
    .Y(_06802_));
 sky130_fd_sc_hd__a21oi_2 _19802_ (.A1(_06727_),
    .A2(_06761_),
    .B1(_06763_),
    .Y(_06803_));
 sky130_fd_sc_hd__xnor2_2 _19803_ (.A(_06802_),
    .B(_06803_),
    .Y(_06804_));
 sky130_fd_sc_hd__or2_2 _19804_ (.A(_06787_),
    .B(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__xor2_2 _19805_ (.A(_06787_),
    .B(_06804_),
    .X(_06806_));
 sky130_fd_sc_hd__o21a_2 _19806_ (.A1(_06751_),
    .A2(_06766_),
    .B1(_06765_),
    .X(_06807_));
 sky130_fd_sc_hd__nand2b_2 _19807_ (.A_N(_06807_),
    .B(_06806_),
    .Y(_06808_));
 sky130_fd_sc_hd__xor2_2 _19808_ (.A(_06806_),
    .B(_06807_),
    .X(_06809_));
 sky130_fd_sc_hd__nand2b_2 _19809_ (.A_N(_06809_),
    .B(_06779_),
    .Y(_06810_));
 sky130_fd_sc_hd__xor2_2 _19810_ (.A(_06779_),
    .B(_06809_),
    .X(_06811_));
 sky130_fd_sc_hd__and2_2 _19811_ (.A(_06770_),
    .B(_06772_),
    .X(_06812_));
 sky130_fd_sc_hd__nor2_2 _19812_ (.A(_06811_),
    .B(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__and2_2 _19813_ (.A(_06811_),
    .B(_06812_),
    .X(_06814_));
 sky130_fd_sc_hd__nor2_2 _19814_ (.A(_06813_),
    .B(_06814_),
    .Y(_06815_));
 sky130_fd_sc_hd__nor2_2 _19815_ (.A(_06774_),
    .B(_06777_),
    .Y(_06816_));
 sky130_fd_sc_hd__or3_2 _19816_ (.A(_06774_),
    .B(_06777_),
    .C(_06815_),
    .X(_06817_));
 sky130_fd_sc_hd__and2b_2 _19817_ (.A_N(_06816_),
    .B(_06815_),
    .X(_06818_));
 sky130_fd_sc_hd__nor2_2 _19818_ (.A(_11258_),
    .B(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__a22o_2 _19819_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[8] ),
    .B1(_06817_),
    .B2(_06819_),
    .X(_01546_));
 sky130_fd_sc_hd__a21o_2 _19820_ (.A1(_06780_),
    .A2(_06786_),
    .B1(_06785_),
    .X(_06820_));
 sky130_fd_sc_hd__o21ba_2 _19821_ (.A1(_06789_),
    .A2(_06791_),
    .B1_N(_06788_),
    .X(_06821_));
 sky130_fd_sc_hd__nor2_2 _19822_ (.A(_06783_),
    .B(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__and2_2 _19823_ (.A(_06783_),
    .B(_06821_),
    .X(_06823_));
 sky130_fd_sc_hd__or2_2 _19824_ (.A(_06822_),
    .B(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__nand2_2 _19825_ (.A(\systolic_inst.B_outs[6][2] ),
    .B(\systolic_inst.A_outs[6][7] ),
    .Y(_06825_));
 sky130_fd_sc_hd__a22oi_2 _19826_ (.A1(\systolic_inst.B_outs[6][4] ),
    .A2(\systolic_inst.A_outs[6][5] ),
    .B1(\systolic_inst.A_outs[6][6] ),
    .B2(\systolic_inst.B_outs[6][3] ),
    .Y(_06826_));
 sky130_fd_sc_hd__and4_2 _19827_ (.A(\systolic_inst.B_outs[6][3] ),
    .B(\systolic_inst.B_outs[6][4] ),
    .C(\systolic_inst.A_outs[6][5] ),
    .D(\systolic_inst.A_outs[6][6] ),
    .X(_06827_));
 sky130_fd_sc_hd__nor2_2 _19828_ (.A(_06826_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__xnor2_2 _19829_ (.A(_06825_),
    .B(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__nand2_2 _19830_ (.A(\systolic_inst.A_outs[6][4] ),
    .B(\systolic_inst.B_outs[6][5] ),
    .Y(_06830_));
 sky130_fd_sc_hd__and4b_2 _19831_ (.A_N(\systolic_inst.A_outs[6][2] ),
    .B(\systolic_inst.A_outs[6][3] ),
    .C(\systolic_inst.B_outs[6][6] ),
    .D(\systolic_inst.B_outs[6][7] ),
    .X(_06831_));
 sky130_fd_sc_hd__o2bb2a_2 _19832_ (.A1_N(\systolic_inst.A_outs[6][3] ),
    .A2_N(\systolic_inst.B_outs[6][6] ),
    .B1(_11278_),
    .B2(\systolic_inst.A_outs[6][2] ),
    .X(_06832_));
 sky130_fd_sc_hd__nor2_2 _19833_ (.A(_06831_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__xnor2_2 _19834_ (.A(_06830_),
    .B(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__o21ba_2 _19835_ (.A1(_06793_),
    .A2(_06795_),
    .B1_N(_06794_),
    .X(_06835_));
 sky130_fd_sc_hd__nand2b_2 _19836_ (.A_N(_06835_),
    .B(_06834_),
    .Y(_06836_));
 sky130_fd_sc_hd__xnor2_2 _19837_ (.A(_06834_),
    .B(_06835_),
    .Y(_06837_));
 sky130_fd_sc_hd__xnor2_2 _19838_ (.A(_06829_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__a21o_2 _19839_ (.A1(_06799_),
    .A2(_06801_),
    .B1(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__nand3_2 _19840_ (.A(_06799_),
    .B(_06801_),
    .C(_06838_),
    .Y(_06840_));
 sky130_fd_sc_hd__nand2_2 _19841_ (.A(_06839_),
    .B(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__xor2_2 _19842_ (.A(_06824_),
    .B(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__o21a_2 _19843_ (.A1(_06802_),
    .A2(_06803_),
    .B1(_06805_),
    .X(_06843_));
 sky130_fd_sc_hd__nand2b_2 _19844_ (.A_N(_06843_),
    .B(_06842_),
    .Y(_06844_));
 sky130_fd_sc_hd__xnor2_2 _19845_ (.A(_06842_),
    .B(_06843_),
    .Y(_06845_));
 sky130_fd_sc_hd__xnor2_2 _19846_ (.A(_06820_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__a21oi_2 _19847_ (.A1(_06808_),
    .A2(_06810_),
    .B1(_06846_),
    .Y(_06847_));
 sky130_fd_sc_hd__and3_2 _19848_ (.A(_06808_),
    .B(_06810_),
    .C(_06846_),
    .X(_06848_));
 sky130_fd_sc_hd__nor2_2 _19849_ (.A(_06847_),
    .B(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__nor2_2 _19850_ (.A(_06813_),
    .B(_06818_),
    .Y(_06850_));
 sky130_fd_sc_hd__xnor2_2 _19851_ (.A(_06849_),
    .B(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__mux2_1 _19852_ (.A0(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[9] ),
    .A1(_06851_),
    .S(\systolic_inst.ce_local ),
    .X(_01547_));
 sky130_fd_sc_hd__and2_2 _19853_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[10] ),
    .X(_06852_));
 sky130_fd_sc_hd__o21ba_2 _19854_ (.A1(_06825_),
    .A2(_06826_),
    .B1_N(_06827_),
    .X(_06853_));
 sky130_fd_sc_hd__nor2_2 _19855_ (.A(_06783_),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__and2_2 _19856_ (.A(_06783_),
    .B(_06853_),
    .X(_06855_));
 sky130_fd_sc_hd__or2_2 _19857_ (.A(_06854_),
    .B(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__a22o_2 _19858_ (.A1(\systolic_inst.B_outs[6][4] ),
    .A2(\systolic_inst.A_outs[6][6] ),
    .B1(\systolic_inst.A_outs[6][7] ),
    .B2(\systolic_inst.B_outs[6][3] ),
    .X(_06857_));
 sky130_fd_sc_hd__and3_2 _19859_ (.A(\systolic_inst.B_outs[6][3] ),
    .B(\systolic_inst.B_outs[6][4] ),
    .C(\systolic_inst.A_outs[6][7] ),
    .X(_06858_));
 sky130_fd_sc_hd__a21bo_2 _19860_ (.A1(\systolic_inst.A_outs[6][6] ),
    .A2(_06858_),
    .B1_N(_06857_),
    .X(_06859_));
 sky130_fd_sc_hd__xor2_2 _19861_ (.A(_06825_),
    .B(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__nand2_2 _19862_ (.A(\systolic_inst.B_outs[6][5] ),
    .B(\systolic_inst.A_outs[6][5] ),
    .Y(_06861_));
 sky130_fd_sc_hd__and4b_2 _19863_ (.A_N(\systolic_inst.A_outs[6][3] ),
    .B(\systolic_inst.A_outs[6][4] ),
    .C(\systolic_inst.B_outs[6][6] ),
    .D(\systolic_inst.B_outs[6][7] ),
    .X(_06862_));
 sky130_fd_sc_hd__o2bb2a_2 _19864_ (.A1_N(\systolic_inst.A_outs[6][4] ),
    .A2_N(\systolic_inst.B_outs[6][6] ),
    .B1(_11278_),
    .B2(\systolic_inst.A_outs[6][3] ),
    .X(_06863_));
 sky130_fd_sc_hd__nor2_2 _19865_ (.A(_06862_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__xnor2_2 _19866_ (.A(_06861_),
    .B(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__o21ba_2 _19867_ (.A1(_06830_),
    .A2(_06832_),
    .B1_N(_06831_),
    .X(_06866_));
 sky130_fd_sc_hd__nand2b_2 _19868_ (.A_N(_06866_),
    .B(_06865_),
    .Y(_06867_));
 sky130_fd_sc_hd__xnor2_2 _19869_ (.A(_06865_),
    .B(_06866_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand2_2 _19870_ (.A(_06860_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__or2_2 _19871_ (.A(_06860_),
    .B(_06868_),
    .X(_06870_));
 sky130_fd_sc_hd__nand2_2 _19872_ (.A(_06869_),
    .B(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__a21bo_2 _19873_ (.A1(_06829_),
    .A2(_06837_),
    .B1_N(_06836_),
    .X(_06872_));
 sky130_fd_sc_hd__nand2b_2 _19874_ (.A_N(_06871_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__xor2_2 _19875_ (.A(_06871_),
    .B(_06872_),
    .X(_06874_));
 sky130_fd_sc_hd__xor2_2 _19876_ (.A(_06856_),
    .B(_06874_),
    .X(_06875_));
 sky130_fd_sc_hd__o21a_2 _19877_ (.A1(_06824_),
    .A2(_06841_),
    .B1(_06839_),
    .X(_06876_));
 sky130_fd_sc_hd__nand2b_2 _19878_ (.A_N(_06876_),
    .B(_06875_),
    .Y(_06877_));
 sky130_fd_sc_hd__xnor2_2 _19879_ (.A(_06875_),
    .B(_06876_),
    .Y(_06878_));
 sky130_fd_sc_hd__nand2_2 _19880_ (.A(_06822_),
    .B(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__or2_2 _19881_ (.A(_06822_),
    .B(_06878_),
    .X(_06880_));
 sky130_fd_sc_hd__nand2_2 _19882_ (.A(_06879_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__a21boi_2 _19883_ (.A1(_06820_),
    .A2(_06845_),
    .B1_N(_06844_),
    .Y(_06882_));
 sky130_fd_sc_hd__or2_2 _19884_ (.A(_06881_),
    .B(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__xor2_2 _19885_ (.A(_06881_),
    .B(_06882_),
    .X(_06884_));
 sky130_fd_sc_hd__nor4b_2 _19886_ (.A(_06816_),
    .B(_06847_),
    .C(_06848_),
    .D_N(_06815_),
    .Y(_06885_));
 sky130_fd_sc_hd__o21ba_2 _19887_ (.A1(_06813_),
    .A2(_06847_),
    .B1_N(_06848_),
    .X(_06886_));
 sky130_fd_sc_hd__or3_2 _19888_ (.A(_06884_),
    .B(_06885_),
    .C(_06886_),
    .X(_06887_));
 sky130_fd_sc_hd__o21ai_2 _19889_ (.A1(_06885_),
    .A2(_06886_),
    .B1(_06884_),
    .Y(_06888_));
 sky130_fd_sc_hd__a31o_2 _19890_ (.A1(\systolic_inst.ce_local ),
    .A2(_06887_),
    .A3(_06888_),
    .B1(_06852_),
    .X(_01548_));
 sky130_fd_sc_hd__o2bb2a_2 _19891_ (.A1_N(\systolic_inst.A_outs[6][6] ),
    .A2_N(_06858_),
    .B1(_06859_),
    .B2(_06825_),
    .X(_06889_));
 sky130_fd_sc_hd__or2_2 _19892_ (.A(_06783_),
    .B(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__nand2_2 _19893_ (.A(_06783_),
    .B(_06889_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand2_2 _19894_ (.A(_06890_),
    .B(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__or2_2 _19895_ (.A(\systolic_inst.B_outs[6][3] ),
    .B(\systolic_inst.B_outs[6][4] ),
    .X(_06893_));
 sky130_fd_sc_hd__and3b_2 _19896_ (.A_N(_06858_),
    .B(_06893_),
    .C(\systolic_inst.A_outs[6][7] ),
    .X(_06894_));
 sky130_fd_sc_hd__xnor2_2 _19897_ (.A(_06825_),
    .B(_06894_),
    .Y(_06895_));
 sky130_fd_sc_hd__nand2_2 _19898_ (.A(\systolic_inst.B_outs[6][5] ),
    .B(\systolic_inst.A_outs[6][6] ),
    .Y(_06896_));
 sky130_fd_sc_hd__and4b_2 _19899_ (.A_N(\systolic_inst.A_outs[6][4] ),
    .B(\systolic_inst.A_outs[6][5] ),
    .C(\systolic_inst.B_outs[6][6] ),
    .D(\systolic_inst.B_outs[6][7] ),
    .X(_06897_));
 sky130_fd_sc_hd__o2bb2a_2 _19900_ (.A1_N(\systolic_inst.A_outs[6][5] ),
    .A2_N(\systolic_inst.B_outs[6][6] ),
    .B1(_11278_),
    .B2(\systolic_inst.A_outs[6][4] ),
    .X(_06898_));
 sky130_fd_sc_hd__nor2_2 _19901_ (.A(_06897_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__xnor2_2 _19902_ (.A(_06896_),
    .B(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__o21ba_2 _19903_ (.A1(_06861_),
    .A2(_06863_),
    .B1_N(_06862_),
    .X(_06901_));
 sky130_fd_sc_hd__nand2b_2 _19904_ (.A_N(_06901_),
    .B(_06900_),
    .Y(_06902_));
 sky130_fd_sc_hd__xnor2_2 _19905_ (.A(_06900_),
    .B(_06901_),
    .Y(_06903_));
 sky130_fd_sc_hd__nand2_2 _19906_ (.A(_06895_),
    .B(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__xnor2_2 _19907_ (.A(_06895_),
    .B(_06903_),
    .Y(_06905_));
 sky130_fd_sc_hd__a21o_2 _19908_ (.A1(_06867_),
    .A2(_06869_),
    .B1(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__nand3_2 _19909_ (.A(_06867_),
    .B(_06869_),
    .C(_06905_),
    .Y(_06907_));
 sky130_fd_sc_hd__nand2_2 _19910_ (.A(_06906_),
    .B(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__xor2_2 _19911_ (.A(_06892_),
    .B(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__o21a_2 _19912_ (.A1(_06856_),
    .A2(_06874_),
    .B1(_06873_),
    .X(_06910_));
 sky130_fd_sc_hd__and2b_2 _19913_ (.A_N(_06910_),
    .B(_06909_),
    .X(_06911_));
 sky130_fd_sc_hd__xnor2_2 _19914_ (.A(_06909_),
    .B(_06910_),
    .Y(_06912_));
 sky130_fd_sc_hd__xnor2_2 _19915_ (.A(_06854_),
    .B(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__and3_2 _19916_ (.A(_06877_),
    .B(_06879_),
    .C(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__a21oi_2 _19917_ (.A1(_06877_),
    .A2(_06879_),
    .B1(_06913_),
    .Y(_06915_));
 sky130_fd_sc_hd__inv_2 _19918_ (.A(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__o211a_2 _19919_ (.A1(_06914_),
    .A2(_06915_),
    .B1(_06883_),
    .C1(_06888_),
    .X(_06917_));
 sky130_fd_sc_hd__a211o_2 _19920_ (.A1(_06883_),
    .A2(_06888_),
    .B1(_06914_),
    .C1(_06915_),
    .X(_06918_));
 sky130_fd_sc_hd__and2b_2 _19921_ (.A_N(_06917_),
    .B(_06918_),
    .X(_06919_));
 sky130_fd_sc_hd__mux2_1 _19922_ (.A0(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[11] ),
    .A1(_06919_),
    .S(\systolic_inst.ce_local ),
    .X(_01549_));
 sky130_fd_sc_hd__a31o_2 _19923_ (.A1(\systolic_inst.B_outs[6][2] ),
    .A2(\systolic_inst.A_outs[6][7] ),
    .A3(_06893_),
    .B1(_06858_),
    .X(_06920_));
 sky130_fd_sc_hd__or2_2 _19924_ (.A(_06782_),
    .B(_06920_),
    .X(_06921_));
 sky130_fd_sc_hd__nand2_2 _19925_ (.A(_06782_),
    .B(_06920_),
    .Y(_06922_));
 sky130_fd_sc_hd__nand2_2 _19926_ (.A(_06921_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__inv_2 _19927_ (.A(_06923_),
    .Y(_06924_));
 sky130_fd_sc_hd__o2bb2a_2 _19928_ (.A1_N(\systolic_inst.B_outs[6][6] ),
    .A2_N(\systolic_inst.A_outs[6][6] ),
    .B1(_11278_),
    .B2(\systolic_inst.A_outs[6][5] ),
    .X(_06925_));
 sky130_fd_sc_hd__and4b_2 _19929_ (.A_N(\systolic_inst.A_outs[6][5] ),
    .B(\systolic_inst.B_outs[6][6] ),
    .C(\systolic_inst.A_outs[6][6] ),
    .D(\systolic_inst.B_outs[6][7] ),
    .X(_06926_));
 sky130_fd_sc_hd__nor2_2 _19930_ (.A(_06925_),
    .B(_06926_),
    .Y(_06927_));
 sky130_fd_sc_hd__nand2_2 _19931_ (.A(\systolic_inst.B_outs[6][5] ),
    .B(\systolic_inst.A_outs[6][7] ),
    .Y(_06928_));
 sky130_fd_sc_hd__xnor2_2 _19932_ (.A(_06927_),
    .B(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__o21ba_2 _19933_ (.A1(_06896_),
    .A2(_06898_),
    .B1_N(_06897_),
    .X(_06930_));
 sky130_fd_sc_hd__nand2b_2 _19934_ (.A_N(_06930_),
    .B(_06929_),
    .Y(_06931_));
 sky130_fd_sc_hd__xnor2_2 _19935_ (.A(_06929_),
    .B(_06930_),
    .Y(_06932_));
 sky130_fd_sc_hd__xnor2_2 _19936_ (.A(_06895_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__a21o_2 _19937_ (.A1(_06902_),
    .A2(_06904_),
    .B1(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__nand3_2 _19938_ (.A(_06902_),
    .B(_06904_),
    .C(_06933_),
    .Y(_06935_));
 sky130_fd_sc_hd__nand2_2 _19939_ (.A(_06934_),
    .B(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__xnor2_2 _19940_ (.A(_06924_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__o21a_2 _19941_ (.A1(_06892_),
    .A2(_06908_),
    .B1(_06906_),
    .X(_06938_));
 sky130_fd_sc_hd__and2b_2 _19942_ (.A_N(_06938_),
    .B(_06937_),
    .X(_06939_));
 sky130_fd_sc_hd__xnor2_2 _19943_ (.A(_06937_),
    .B(_06938_),
    .Y(_06940_));
 sky130_fd_sc_hd__and2b_2 _19944_ (.A_N(_06890_),
    .B(_06940_),
    .X(_06941_));
 sky130_fd_sc_hd__xor2_2 _19945_ (.A(_06890_),
    .B(_06940_),
    .X(_06942_));
 sky130_fd_sc_hd__a21oi_2 _19946_ (.A1(_06854_),
    .A2(_06912_),
    .B1(_06911_),
    .Y(_06943_));
 sky130_fd_sc_hd__or2_2 _19947_ (.A(_06942_),
    .B(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__nand2_2 _19948_ (.A(_06942_),
    .B(_06943_),
    .Y(_06945_));
 sky130_fd_sc_hd__and2_2 _19949_ (.A(_06944_),
    .B(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__inv_2 _19950_ (.A(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__a31o_2 _19951_ (.A1(_06883_),
    .A2(_06888_),
    .A3(_06916_),
    .B1(_06914_),
    .X(_06948_));
 sky130_fd_sc_hd__a311o_2 _19952_ (.A1(_06883_),
    .A2(_06888_),
    .A3(_06916_),
    .B1(_06947_),
    .C1(_06914_),
    .X(_06949_));
 sky130_fd_sc_hd__xnor2_2 _19953_ (.A(_06946_),
    .B(_06948_),
    .Y(_06950_));
 sky130_fd_sc_hd__mux2_1 _19954_ (.A0(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[12] ),
    .A1(_06950_),
    .S(\systolic_inst.ce_local ),
    .X(_01550_));
 sky130_fd_sc_hd__nand2_2 _19955_ (.A(\systolic_inst.B_outs[6][6] ),
    .B(\systolic_inst.A_outs[6][7] ),
    .Y(_06951_));
 sky130_fd_sc_hd__or2_2 _19956_ (.A(\systolic_inst.A_outs[6][6] ),
    .B(_11278_),
    .X(_06952_));
 sky130_fd_sc_hd__and2_2 _19957_ (.A(_06951_),
    .B(_06952_),
    .X(_06953_));
 sky130_fd_sc_hd__nor2_2 _19958_ (.A(_06951_),
    .B(_06952_),
    .Y(_06954_));
 sky130_fd_sc_hd__nor2_2 _19959_ (.A(_06953_),
    .B(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__xnor2_2 _19960_ (.A(_06928_),
    .B(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__o21ba_2 _19961_ (.A1(_06925_),
    .A2(_06928_),
    .B1_N(_06926_),
    .X(_06957_));
 sky130_fd_sc_hd__nand2b_2 _19962_ (.A_N(_06957_),
    .B(_06956_),
    .Y(_06958_));
 sky130_fd_sc_hd__xnor2_2 _19963_ (.A(_06956_),
    .B(_06957_),
    .Y(_06959_));
 sky130_fd_sc_hd__nand2_2 _19964_ (.A(_06895_),
    .B(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__or2_2 _19965_ (.A(_06895_),
    .B(_06959_),
    .X(_06961_));
 sky130_fd_sc_hd__nand2_2 _19966_ (.A(_06960_),
    .B(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__a21bo_2 _19967_ (.A1(_06895_),
    .A2(_06932_),
    .B1_N(_06931_),
    .X(_06963_));
 sky130_fd_sc_hd__nand2b_2 _19968_ (.A_N(_06962_),
    .B(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__xor2_2 _19969_ (.A(_06962_),
    .B(_06963_),
    .X(_06965_));
 sky130_fd_sc_hd__xnor2_2 _19970_ (.A(_06924_),
    .B(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__o21a_2 _19971_ (.A1(_06923_),
    .A2(_06936_),
    .B1(_06934_),
    .X(_06967_));
 sky130_fd_sc_hd__and2b_2 _19972_ (.A_N(_06967_),
    .B(_06966_),
    .X(_06968_));
 sky130_fd_sc_hd__and2b_2 _19973_ (.A_N(_06966_),
    .B(_06967_),
    .X(_06969_));
 sky130_fd_sc_hd__nor2_2 _19974_ (.A(_06968_),
    .B(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__xnor2_2 _19975_ (.A(_06922_),
    .B(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__nor3_2 _19976_ (.A(_06939_),
    .B(_06941_),
    .C(_06971_),
    .Y(_06972_));
 sky130_fd_sc_hd__o21ai_2 _19977_ (.A1(_06939_),
    .A2(_06941_),
    .B1(_06971_),
    .Y(_06973_));
 sky130_fd_sc_hd__and2b_2 _19978_ (.A_N(_06972_),
    .B(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__and2_2 _19979_ (.A(_06944_),
    .B(_06949_),
    .X(_06975_));
 sky130_fd_sc_hd__xnor2_2 _19980_ (.A(_06974_),
    .B(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__mux2_1 _19981_ (.A0(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[13] ),
    .A1(_06976_),
    .S(\systolic_inst.ce_local ),
    .X(_01551_));
 sky130_fd_sc_hd__a31o_2 _19982_ (.A1(\systolic_inst.B_outs[6][5] ),
    .A2(\systolic_inst.A_outs[6][7] ),
    .A3(_06955_),
    .B1(_06954_),
    .X(_06977_));
 sky130_fd_sc_hd__nand3_2 _19983_ (.A(\systolic_inst.B_outs[6][5] ),
    .B(\systolic_inst.B_outs[6][6] ),
    .C(\systolic_inst.A_outs[6][7] ),
    .Y(_06978_));
 sky130_fd_sc_hd__o211a_2 _19984_ (.A1(_11278_),
    .A2(\systolic_inst.A_outs[6][7] ),
    .B1(_06928_),
    .C1(_06951_),
    .X(_06979_));
 sky130_fd_sc_hd__a21oi_2 _19985_ (.A1(_06977_),
    .A2(_06978_),
    .B1(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__or2_2 _19986_ (.A(_06895_),
    .B(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__nand2_2 _19987_ (.A(_06895_),
    .B(_06980_),
    .Y(_06982_));
 sky130_fd_sc_hd__nand2_2 _19988_ (.A(_06981_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__a21oi_2 _19989_ (.A1(_06958_),
    .A2(_06960_),
    .B1(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__and3_2 _19990_ (.A(_06958_),
    .B(_06960_),
    .C(_06983_),
    .X(_06985_));
 sky130_fd_sc_hd__nor2_2 _19991_ (.A(_06984_),
    .B(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__xnor2_2 _19992_ (.A(_06923_),
    .B(_06986_),
    .Y(_06987_));
 sky130_fd_sc_hd__o21a_2 _19993_ (.A1(_06923_),
    .A2(_06965_),
    .B1(_06964_),
    .X(_06988_));
 sky130_fd_sc_hd__and2b_2 _19994_ (.A_N(_06988_),
    .B(_06987_),
    .X(_06989_));
 sky130_fd_sc_hd__and2b_2 _19995_ (.A_N(_06987_),
    .B(_06988_),
    .X(_06990_));
 sky130_fd_sc_hd__nor2_2 _19996_ (.A(_06989_),
    .B(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__xnor2_2 _19997_ (.A(_06922_),
    .B(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__o21ba_2 _19998_ (.A1(_06922_),
    .A2(_06969_),
    .B1_N(_06968_),
    .X(_06993_));
 sky130_fd_sc_hd__nand2b_2 _19999_ (.A_N(_06993_),
    .B(_06992_),
    .Y(_06994_));
 sky130_fd_sc_hd__xnor2_2 _20000_ (.A(_06992_),
    .B(_06993_),
    .Y(_06995_));
 sky130_fd_sc_hd__or2_2 _20001_ (.A(_06944_),
    .B(_06972_),
    .X(_06996_));
 sky130_fd_sc_hd__o211ai_2 _20002_ (.A1(_06949_),
    .A2(_06972_),
    .B1(_06973_),
    .C1(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__nand2_2 _20003_ (.A(_06995_),
    .B(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__xor2_2 _20004_ (.A(_06995_),
    .B(_06997_),
    .X(_06999_));
 sky130_fd_sc_hd__mux2_1 _20005_ (.A0(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[14] ),
    .A1(_06999_),
    .S(\systolic_inst.ce_local ),
    .X(_01552_));
 sky130_fd_sc_hd__a31o_2 _20006_ (.A1(_06782_),
    .A2(_06920_),
    .A3(_06991_),
    .B1(_06989_),
    .X(_07000_));
 sky130_fd_sc_hd__a21oi_2 _20007_ (.A1(_06924_),
    .A2(_06986_),
    .B1(_06984_),
    .Y(_07001_));
 sky130_fd_sc_hd__xnor2_2 _20008_ (.A(_06921_),
    .B(_06981_),
    .Y(_07002_));
 sky130_fd_sc_hd__xnor2_2 _20009_ (.A(_07001_),
    .B(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__xnor2_2 _20010_ (.A(_07000_),
    .B(_07003_),
    .Y(_07004_));
 sky130_fd_sc_hd__and3_2 _20011_ (.A(\systolic_inst.ce_local ),
    .B(_06994_),
    .C(_07004_),
    .X(_07005_));
 sky130_fd_sc_hd__a22o_2 _20012_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B1(_06998_),
    .B2(_07005_),
    .X(_01553_));
 sky130_fd_sc_hd__a21o_2 _20013_ (.A1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[6][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_07006_));
 sky130_fd_sc_hd__a21oi_2 _20014_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[6][0] ),
    .Y(_07007_));
 sky130_fd_sc_hd__a21oi_2 _20015_ (.A1(\systolic_inst.ce_local ),
    .A2(_07006_),
    .B1(_07007_),
    .Y(_01554_));
 sky130_fd_sc_hd__and2_2 _20016_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[6][1] ),
    .X(_07008_));
 sky130_fd_sc_hd__nand2_2 _20017_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[6][1] ),
    .Y(_07009_));
 sky130_fd_sc_hd__or2_2 _20018_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[6][1] ),
    .X(_07010_));
 sky130_fd_sc_hd__and4_2 _20019_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[6][0] ),
    .C(_07009_),
    .D(_07010_),
    .X(_07011_));
 sky130_fd_sc_hd__inv_2 _20020_ (.A(_07011_),
    .Y(_07012_));
 sky130_fd_sc_hd__a22o_2 _20021_ (.A1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[6][0] ),
    .B1(_07009_),
    .B2(_07010_),
    .X(_07013_));
 sky130_fd_sc_hd__a32o_2 _20022_ (.A1(_11712_),
    .A2(_07012_),
    .A3(_07013_),
    .B1(\systolic_inst.acc_wires[6][1] ),
    .B2(_11258_),
    .X(_01555_));
 sky130_fd_sc_hd__nand2_2 _20023_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[6][2] ),
    .Y(_07014_));
 sky130_fd_sc_hd__or2_2 _20024_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[6][2] ),
    .X(_07015_));
 sky130_fd_sc_hd__a31o_2 _20025_ (.A1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[6][0] ),
    .A3(_07010_),
    .B1(_07008_),
    .X(_07016_));
 sky130_fd_sc_hd__a21o_2 _20026_ (.A1(_07014_),
    .A2(_07015_),
    .B1(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__and3_2 _20027_ (.A(_07014_),
    .B(_07015_),
    .C(_07016_),
    .X(_07018_));
 sky130_fd_sc_hd__inv_2 _20028_ (.A(_07018_),
    .Y(_07019_));
 sky130_fd_sc_hd__a32o_2 _20029_ (.A1(_11712_),
    .A2(_07017_),
    .A3(_07019_),
    .B1(\systolic_inst.acc_wires[6][2] ),
    .B2(_11258_),
    .X(_01556_));
 sky130_fd_sc_hd__nand2_2 _20030_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[6][3] ),
    .Y(_07020_));
 sky130_fd_sc_hd__or2_2 _20031_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[6][3] ),
    .X(_07021_));
 sky130_fd_sc_hd__a21bo_2 _20032_ (.A1(_07015_),
    .A2(_07016_),
    .B1_N(_07014_),
    .X(_07022_));
 sky130_fd_sc_hd__a21o_2 _20033_ (.A1(_07020_),
    .A2(_07021_),
    .B1(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__and3_2 _20034_ (.A(_07020_),
    .B(_07021_),
    .C(_07022_),
    .X(_07024_));
 sky130_fd_sc_hd__inv_2 _20035_ (.A(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__a32o_2 _20036_ (.A1(_11712_),
    .A2(_07023_),
    .A3(_07025_),
    .B1(\systolic_inst.acc_wires[6][3] ),
    .B2(_11258_),
    .X(_01557_));
 sky130_fd_sc_hd__nand2_2 _20037_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[6][4] ),
    .Y(_07026_));
 sky130_fd_sc_hd__or2_2 _20038_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[6][4] ),
    .X(_07027_));
 sky130_fd_sc_hd__a21bo_2 _20039_ (.A1(_07021_),
    .A2(_07022_),
    .B1_N(_07020_),
    .X(_07028_));
 sky130_fd_sc_hd__a21o_2 _20040_ (.A1(_07026_),
    .A2(_07027_),
    .B1(_07028_),
    .X(_07029_));
 sky130_fd_sc_hd__and3_2 _20041_ (.A(_07026_),
    .B(_07027_),
    .C(_07028_),
    .X(_07030_));
 sky130_fd_sc_hd__inv_2 _20042_ (.A(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__a32o_2 _20043_ (.A1(_11712_),
    .A2(_07029_),
    .A3(_07031_),
    .B1(\systolic_inst.acc_wires[6][4] ),
    .B2(_11258_),
    .X(_01558_));
 sky130_fd_sc_hd__nand2_2 _20044_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[6][5] ),
    .Y(_07032_));
 sky130_fd_sc_hd__or2_2 _20045_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[6][5] ),
    .X(_07033_));
 sky130_fd_sc_hd__a21bo_2 _20046_ (.A1(_07027_),
    .A2(_07028_),
    .B1_N(_07026_),
    .X(_07034_));
 sky130_fd_sc_hd__a21o_2 _20047_ (.A1(_07032_),
    .A2(_07033_),
    .B1(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__and3_2 _20048_ (.A(_07032_),
    .B(_07033_),
    .C(_07034_),
    .X(_07036_));
 sky130_fd_sc_hd__inv_2 _20049_ (.A(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__a32o_2 _20050_ (.A1(_11712_),
    .A2(_07035_),
    .A3(_07037_),
    .B1(\systolic_inst.acc_wires[6][5] ),
    .B2(_11258_),
    .X(_01559_));
 sky130_fd_sc_hd__nand2_2 _20051_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[6][6] ),
    .Y(_07038_));
 sky130_fd_sc_hd__or2_2 _20052_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[6][6] ),
    .X(_07039_));
 sky130_fd_sc_hd__a21bo_2 _20053_ (.A1(_07033_),
    .A2(_07034_),
    .B1_N(_07032_),
    .X(_07040_));
 sky130_fd_sc_hd__a21o_2 _20054_ (.A1(_07038_),
    .A2(_07039_),
    .B1(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__and3_2 _20055_ (.A(_07038_),
    .B(_07039_),
    .C(_07040_),
    .X(_07042_));
 sky130_fd_sc_hd__inv_2 _20056_ (.A(_07042_),
    .Y(_07043_));
 sky130_fd_sc_hd__a32o_2 _20057_ (.A1(_11712_),
    .A2(_07041_),
    .A3(_07043_),
    .B1(\systolic_inst.acc_wires[6][6] ),
    .B2(_11258_),
    .X(_01560_));
 sky130_fd_sc_hd__nand2_2 _20058_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[6][7] ),
    .Y(_07044_));
 sky130_fd_sc_hd__or2_2 _20059_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[6][7] ),
    .X(_07045_));
 sky130_fd_sc_hd__a21bo_2 _20060_ (.A1(_07039_),
    .A2(_07040_),
    .B1_N(_07038_),
    .X(_07046_));
 sky130_fd_sc_hd__a21o_2 _20061_ (.A1(_07044_),
    .A2(_07045_),
    .B1(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__nand3_2 _20062_ (.A(_07044_),
    .B(_07045_),
    .C(_07046_),
    .Y(_07048_));
 sky130_fd_sc_hd__a32o_2 _20063_ (.A1(_11712_),
    .A2(_07047_),
    .A3(_07048_),
    .B1(\systolic_inst.acc_wires[6][7] ),
    .B2(_11258_),
    .X(_01561_));
 sky130_fd_sc_hd__a21bo_2 _20064_ (.A1(_07045_),
    .A2(_07046_),
    .B1_N(_07044_),
    .X(_07049_));
 sky130_fd_sc_hd__xor2_2 _20065_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[6][8] ),
    .X(_07050_));
 sky130_fd_sc_hd__and2_2 _20066_ (.A(_07049_),
    .B(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__o21ai_2 _20067_ (.A1(_07049_),
    .A2(_07050_),
    .B1(_11712_),
    .Y(_07052_));
 sky130_fd_sc_hd__a2bb2o_2 _20068_ (.A1_N(_07052_),
    .A2_N(_07051_),
    .B1(\systolic_inst.acc_wires[6][8] ),
    .B2(_11258_),
    .X(_01562_));
 sky130_fd_sc_hd__xor2_2 _20069_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[6][9] ),
    .X(_07053_));
 sky130_fd_sc_hd__a211o_2 _20070_ (.A1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[6][8] ),
    .B1(_07051_),
    .C1(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__nand2_2 _20071_ (.A(_07050_),
    .B(_07053_),
    .Y(_07055_));
 sky130_fd_sc_hd__nand2_2 _20072_ (.A(_07051_),
    .B(_07053_),
    .Y(_07056_));
 sky130_fd_sc_hd__and3_2 _20073_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[6][8] ),
    .C(_07053_),
    .X(_07057_));
 sky130_fd_sc_hd__nor2_2 _20074_ (.A(_11713_),
    .B(_07057_),
    .Y(_07058_));
 sky130_fd_sc_hd__a32o_2 _20075_ (.A1(_07054_),
    .A2(_07056_),
    .A3(_07058_),
    .B1(\systolic_inst.acc_wires[6][9] ),
    .B2(_11258_),
    .X(_01563_));
 sky130_fd_sc_hd__nand2_2 _20076_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[6][10] ),
    .Y(_07059_));
 sky130_fd_sc_hd__or2_2 _20077_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[6][10] ),
    .X(_07060_));
 sky130_fd_sc_hd__and2_2 _20078_ (.A(_07059_),
    .B(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__a21oi_2 _20079_ (.A1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[6][9] ),
    .B1(_07057_),
    .Y(_07062_));
 sky130_fd_sc_hd__nand2_2 _20080_ (.A(_07056_),
    .B(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__xor2_2 _20081_ (.A(_07061_),
    .B(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__a22o_2 _20082_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][10] ),
    .B1(_11712_),
    .B2(_07064_),
    .X(_01564_));
 sky130_fd_sc_hd__nor2_2 _20083_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[6][11] ),
    .Y(_07065_));
 sky130_fd_sc_hd__or2_2 _20084_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[6][11] ),
    .X(_07066_));
 sky130_fd_sc_hd__nand2_2 _20085_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[6][11] ),
    .Y(_07067_));
 sky130_fd_sc_hd__nand2_2 _20086_ (.A(_07066_),
    .B(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__a21bo_2 _20087_ (.A1(_07061_),
    .A2(_07063_),
    .B1_N(_07059_),
    .X(_07069_));
 sky130_fd_sc_hd__xnor2_2 _20088_ (.A(_07068_),
    .B(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__a22o_2 _20089_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][11] ),
    .B1(_11712_),
    .B2(_07070_),
    .X(_01565_));
 sky130_fd_sc_hd__nand3_2 _20090_ (.A(_07061_),
    .B(_07066_),
    .C(_07067_),
    .Y(_07071_));
 sky130_fd_sc_hd__nor2_2 _20091_ (.A(_07055_),
    .B(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__o2bb2a_2 _20092_ (.A1_N(_07049_),
    .A2_N(_07072_),
    .B1(_07062_),
    .B2(_07071_),
    .X(_07073_));
 sky130_fd_sc_hd__o21a_2 _20093_ (.A1(_07059_),
    .A2(_07065_),
    .B1(_07067_),
    .X(_07074_));
 sky130_fd_sc_hd__xnor2_2 _20094_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[6][12] ),
    .Y(_07075_));
 sky130_fd_sc_hd__and3_2 _20095_ (.A(_07073_),
    .B(_07074_),
    .C(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__a21oi_2 _20096_ (.A1(_07073_),
    .A2(_07074_),
    .B1(_07075_),
    .Y(_07077_));
 sky130_fd_sc_hd__nor2_2 _20097_ (.A(_07076_),
    .B(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__a22o_2 _20098_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][12] ),
    .B1(_11712_),
    .B2(_07078_),
    .X(_01566_));
 sky130_fd_sc_hd__xor2_2 _20099_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[6][13] ),
    .X(_07079_));
 sky130_fd_sc_hd__a211o_2 _20100_ (.A1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[6][12] ),
    .B1(_07077_),
    .C1(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__nand2b_2 _20101_ (.A_N(_07075_),
    .B(_07079_),
    .Y(_07081_));
 sky130_fd_sc_hd__a21o_2 _20102_ (.A1(_07073_),
    .A2(_07074_),
    .B1(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__and3_2 _20103_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[6][12] ),
    .C(_07079_),
    .X(_07083_));
 sky130_fd_sc_hd__nor2_2 _20104_ (.A(_11713_),
    .B(_07083_),
    .Y(_07084_));
 sky130_fd_sc_hd__a32o_2 _20105_ (.A1(_07080_),
    .A2(_07082_),
    .A3(_07084_),
    .B1(\systolic_inst.acc_wires[6][13] ),
    .B2(_11258_),
    .X(_01567_));
 sky130_fd_sc_hd__or2_2 _20106_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[6][14] ),
    .X(_07085_));
 sky130_fd_sc_hd__nand2_2 _20107_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[6][14] ),
    .Y(_07086_));
 sky130_fd_sc_hd__and2_2 _20108_ (.A(_07085_),
    .B(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__nand2_2 _20109_ (.A(_07085_),
    .B(_07086_),
    .Y(_07088_));
 sky130_fd_sc_hd__a21oi_2 _20110_ (.A1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[6][13] ),
    .B1(_07083_),
    .Y(_07089_));
 sky130_fd_sc_hd__nand2_2 _20111_ (.A(_07082_),
    .B(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__nand2_2 _20112_ (.A(_07087_),
    .B(_07090_),
    .Y(_07091_));
 sky130_fd_sc_hd__or2_2 _20113_ (.A(_07087_),
    .B(_07090_),
    .X(_07092_));
 sky130_fd_sc_hd__a32o_2 _20114_ (.A1(_11712_),
    .A2(_07091_),
    .A3(_07092_),
    .B1(\systolic_inst.acc_wires[6][14] ),
    .B2(_11258_),
    .X(_01568_));
 sky130_fd_sc_hd__nor2_2 _20115_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][15] ),
    .Y(_07093_));
 sky130_fd_sc_hd__and2_2 _20116_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][15] ),
    .X(_07094_));
 sky130_fd_sc_hd__or2_2 _20117_ (.A(_07093_),
    .B(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__a21oi_2 _20118_ (.A1(_07086_),
    .A2(_07091_),
    .B1(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__a31o_2 _20119_ (.A1(_07086_),
    .A2(_07091_),
    .A3(_07095_),
    .B1(_11713_),
    .X(_07097_));
 sky130_fd_sc_hd__a2bb2o_2 _20120_ (.A1_N(_07097_),
    .A2_N(_07096_),
    .B1(\systolic_inst.acc_wires[6][15] ),
    .B2(_11258_),
    .X(_01569_));
 sky130_fd_sc_hd__a211o_2 _20121_ (.A1(_07082_),
    .A2(_07089_),
    .B1(_07095_),
    .C1(_07088_),
    .X(_07098_));
 sky130_fd_sc_hd__o21ba_2 _20122_ (.A1(_07086_),
    .A2(_07093_),
    .B1_N(_07094_),
    .X(_07099_));
 sky130_fd_sc_hd__and2_2 _20123_ (.A(_07098_),
    .B(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__xnor2_2 _20124_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][16] ),
    .Y(_07101_));
 sky130_fd_sc_hd__nand2_2 _20125_ (.A(_07100_),
    .B(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__nor2_2 _20126_ (.A(_07100_),
    .B(_07101_),
    .Y(_07103_));
 sky130_fd_sc_hd__nor2_2 _20127_ (.A(_11713_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__a22o_2 _20128_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][16] ),
    .B1(_07102_),
    .B2(_07104_),
    .X(_01570_));
 sky130_fd_sc_hd__xor2_2 _20129_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][17] ),
    .X(_07105_));
 sky130_fd_sc_hd__inv_2 _20130_ (.A(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__a21oi_2 _20131_ (.A1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[6][16] ),
    .B1(_07103_),
    .Y(_07107_));
 sky130_fd_sc_hd__xnor2_2 _20132_ (.A(_07105_),
    .B(_07107_),
    .Y(_07108_));
 sky130_fd_sc_hd__a22o_2 _20133_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][17] ),
    .B1(_11712_),
    .B2(_07108_),
    .X(_01571_));
 sky130_fd_sc_hd__or2_2 _20134_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][18] ),
    .X(_07109_));
 sky130_fd_sc_hd__nand2_2 _20135_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][18] ),
    .Y(_07110_));
 sky130_fd_sc_hd__nand2_2 _20136_ (.A(_07109_),
    .B(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__o21a_2 _20137_ (.A1(\systolic_inst.acc_wires[6][16] ),
    .A2(\systolic_inst.acc_wires[6][17] ),
    .B1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .X(_07112_));
 sky130_fd_sc_hd__a21oi_2 _20138_ (.A1(_07103_),
    .A2(_07105_),
    .B1(_07112_),
    .Y(_07113_));
 sky130_fd_sc_hd__xor2_2 _20139_ (.A(_07111_),
    .B(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__a22o_2 _20140_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][18] ),
    .B1(_11712_),
    .B2(_07114_),
    .X(_01572_));
 sky130_fd_sc_hd__xnor2_2 _20141_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][19] ),
    .Y(_07115_));
 sky130_fd_sc_hd__o21ai_2 _20142_ (.A1(_07111_),
    .A2(_07113_),
    .B1(_07110_),
    .Y(_07116_));
 sky130_fd_sc_hd__xnor2_2 _20143_ (.A(_07115_),
    .B(_07116_),
    .Y(_07117_));
 sky130_fd_sc_hd__a22o_2 _20144_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][19] ),
    .B1(_11712_),
    .B2(_07117_),
    .X(_01573_));
 sky130_fd_sc_hd__or2_2 _20145_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][20] ),
    .X(_07118_));
 sky130_fd_sc_hd__nand2_2 _20146_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][20] ),
    .Y(_07119_));
 sky130_fd_sc_hd__and2_2 _20147_ (.A(_07118_),
    .B(_07119_),
    .X(_07120_));
 sky130_fd_sc_hd__or4_2 _20148_ (.A(_07101_),
    .B(_07106_),
    .C(_07111_),
    .D(_07115_),
    .X(_07121_));
 sky130_fd_sc_hd__nor2_2 _20149_ (.A(_07100_),
    .B(_07121_),
    .Y(_07122_));
 sky130_fd_sc_hd__o41a_2 _20150_ (.A1(\systolic_inst.acc_wires[6][16] ),
    .A2(\systolic_inst.acc_wires[6][17] ),
    .A3(\systolic_inst.acc_wires[6][18] ),
    .A4(\systolic_inst.acc_wires[6][19] ),
    .B1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .X(_07123_));
 sky130_fd_sc_hd__or3_2 _20151_ (.A(_07120_),
    .B(_07122_),
    .C(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__o21ai_2 _20152_ (.A1(_07122_),
    .A2(_07123_),
    .B1(_07120_),
    .Y(_07125_));
 sky130_fd_sc_hd__a32o_2 _20153_ (.A1(_11712_),
    .A2(_07124_),
    .A3(_07125_),
    .B1(\systolic_inst.acc_wires[6][20] ),
    .B2(_11258_),
    .X(_01574_));
 sky130_fd_sc_hd__xnor2_2 _20154_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][21] ),
    .Y(_07126_));
 sky130_fd_sc_hd__inv_2 _20155_ (.A(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__a21oi_2 _20156_ (.A1(_07119_),
    .A2(_07125_),
    .B1(_07126_),
    .Y(_07128_));
 sky130_fd_sc_hd__a31o_2 _20157_ (.A1(_07119_),
    .A2(_07125_),
    .A3(_07126_),
    .B1(_11713_),
    .X(_07129_));
 sky130_fd_sc_hd__a2bb2o_2 _20158_ (.A1_N(_07129_),
    .A2_N(_07128_),
    .B1(\systolic_inst.acc_wires[6][21] ),
    .B2(_11258_),
    .X(_01575_));
 sky130_fd_sc_hd__or2_2 _20159_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][22] ),
    .X(_07130_));
 sky130_fd_sc_hd__nand2_2 _20160_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][22] ),
    .Y(_07131_));
 sky130_fd_sc_hd__and2_2 _20161_ (.A(_07130_),
    .B(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__o21a_2 _20162_ (.A1(\systolic_inst.acc_wires[6][20] ),
    .A2(\systolic_inst.acc_wires[6][21] ),
    .B1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .X(_07133_));
 sky130_fd_sc_hd__nor2_2 _20163_ (.A(_07125_),
    .B(_07126_),
    .Y(_07134_));
 sky130_fd_sc_hd__o21ai_2 _20164_ (.A1(_07133_),
    .A2(_07134_),
    .B1(_07132_),
    .Y(_07135_));
 sky130_fd_sc_hd__or3_2 _20165_ (.A(_07132_),
    .B(_07133_),
    .C(_07134_),
    .X(_07136_));
 sky130_fd_sc_hd__a32o_2 _20166_ (.A1(_11712_),
    .A2(_07135_),
    .A3(_07136_),
    .B1(\systolic_inst.acc_wires[6][22] ),
    .B2(_11258_),
    .X(_01576_));
 sky130_fd_sc_hd__xor2_2 _20167_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][23] ),
    .X(_07137_));
 sky130_fd_sc_hd__inv_2 _20168_ (.A(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__nand3_2 _20169_ (.A(_07131_),
    .B(_07135_),
    .C(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__a21o_2 _20170_ (.A1(_07131_),
    .A2(_07135_),
    .B1(_07138_),
    .X(_07140_));
 sky130_fd_sc_hd__a32o_2 _20171_ (.A1(_11712_),
    .A2(_07139_),
    .A3(_07140_),
    .B1(\systolic_inst.acc_wires[6][23] ),
    .B2(_11258_),
    .X(_01577_));
 sky130_fd_sc_hd__nand4_2 _20172_ (.A(_07120_),
    .B(_07127_),
    .C(_07132_),
    .D(_07137_),
    .Y(_07141_));
 sky130_fd_sc_hd__a211o_2 _20173_ (.A1(_07098_),
    .A2(_07099_),
    .B1(_07121_),
    .C1(_07141_),
    .X(_07142_));
 sky130_fd_sc_hd__o41a_2 _20174_ (.A1(\systolic_inst.acc_wires[6][20] ),
    .A2(\systolic_inst.acc_wires[6][21] ),
    .A3(\systolic_inst.acc_wires[6][22] ),
    .A4(\systolic_inst.acc_wires[6][23] ),
    .B1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .X(_07143_));
 sky130_fd_sc_hd__nor2_2 _20175_ (.A(_07123_),
    .B(_07143_),
    .Y(_07144_));
 sky130_fd_sc_hd__nor2_2 _20176_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][24] ),
    .Y(_07145_));
 sky130_fd_sc_hd__and2_2 _20177_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][24] ),
    .X(_07146_));
 sky130_fd_sc_hd__or2_2 _20178_ (.A(_07145_),
    .B(_07146_),
    .X(_07147_));
 sky130_fd_sc_hd__and3_2 _20179_ (.A(_07142_),
    .B(_07144_),
    .C(_07147_),
    .X(_07148_));
 sky130_fd_sc_hd__a21oi_2 _20180_ (.A1(_07142_),
    .A2(_07144_),
    .B1(_07147_),
    .Y(_07149_));
 sky130_fd_sc_hd__nor2_2 _20181_ (.A(_07148_),
    .B(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__a22o_2 _20182_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][24] ),
    .B1(_11712_),
    .B2(_07150_),
    .X(_01578_));
 sky130_fd_sc_hd__xor2_2 _20183_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][25] ),
    .X(_07151_));
 sky130_fd_sc_hd__or3_2 _20184_ (.A(_07146_),
    .B(_07149_),
    .C(_07151_),
    .X(_07152_));
 sky130_fd_sc_hd__o21ai_2 _20185_ (.A1(_07146_),
    .A2(_07149_),
    .B1(_07151_),
    .Y(_07153_));
 sky130_fd_sc_hd__a32o_2 _20186_ (.A1(_11712_),
    .A2(_07152_),
    .A3(_07153_),
    .B1(\systolic_inst.acc_wires[6][25] ),
    .B2(_11258_),
    .X(_01579_));
 sky130_fd_sc_hd__or2_2 _20187_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][26] ),
    .X(_07154_));
 sky130_fd_sc_hd__nand2_2 _20188_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][26] ),
    .Y(_07155_));
 sky130_fd_sc_hd__nand2_2 _20189_ (.A(_07154_),
    .B(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__o21a_2 _20190_ (.A1(\systolic_inst.acc_wires[6][24] ),
    .A2(\systolic_inst.acc_wires[6][25] ),
    .B1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .X(_07157_));
 sky130_fd_sc_hd__a21o_2 _20191_ (.A1(_07149_),
    .A2(_07151_),
    .B1(_07157_),
    .X(_07158_));
 sky130_fd_sc_hd__xnor2_2 _20192_ (.A(_07156_),
    .B(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__a22o_2 _20193_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][26] ),
    .B1(_11712_),
    .B2(_07159_),
    .X(_01580_));
 sky130_fd_sc_hd__xnor2_2 _20194_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][27] ),
    .Y(_07160_));
 sky130_fd_sc_hd__a21bo_2 _20195_ (.A1(_07154_),
    .A2(_07158_),
    .B1_N(_07155_),
    .X(_07161_));
 sky130_fd_sc_hd__xnor2_2 _20196_ (.A(_07160_),
    .B(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__a22o_2 _20197_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][27] ),
    .B1(_11712_),
    .B2(_07162_),
    .X(_01581_));
 sky130_fd_sc_hd__nor2_2 _20198_ (.A(_07156_),
    .B(_07160_),
    .Y(_07163_));
 sky130_fd_sc_hd__o21a_2 _20199_ (.A1(\systolic_inst.acc_wires[6][26] ),
    .A2(\systolic_inst.acc_wires[6][27] ),
    .B1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .X(_07164_));
 sky130_fd_sc_hd__a311oi_2 _20200_ (.A1(_07149_),
    .A2(_07151_),
    .A3(_07163_),
    .B1(_07164_),
    .C1(_07157_),
    .Y(_07165_));
 sky130_fd_sc_hd__or2_2 _20201_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][28] ),
    .X(_07166_));
 sky130_fd_sc_hd__nand2_2 _20202_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][28] ),
    .Y(_07167_));
 sky130_fd_sc_hd__nand2_2 _20203_ (.A(_07166_),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__xor2_2 _20204_ (.A(_07165_),
    .B(_07168_),
    .X(_07169_));
 sky130_fd_sc_hd__a22o_2 _20205_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][28] ),
    .B1(_11712_),
    .B2(_07169_),
    .X(_01582_));
 sky130_fd_sc_hd__xor2_2 _20206_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][29] ),
    .X(_07170_));
 sky130_fd_sc_hd__inv_2 _20207_ (.A(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__o21a_2 _20208_ (.A1(_07165_),
    .A2(_07168_),
    .B1(_07167_),
    .X(_07172_));
 sky130_fd_sc_hd__xnor2_2 _20209_ (.A(_07170_),
    .B(_07172_),
    .Y(_07173_));
 sky130_fd_sc_hd__a22o_2 _20210_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[6][29] ),
    .B1(_11712_),
    .B2(_07173_),
    .X(_01583_));
 sky130_fd_sc_hd__o21ai_2 _20211_ (.A1(\systolic_inst.acc_wires[6][28] ),
    .A2(\systolic_inst.acc_wires[6][29] ),
    .B1(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .Y(_07174_));
 sky130_fd_sc_hd__o31a_2 _20212_ (.A1(_07165_),
    .A2(_07168_),
    .A3(_07171_),
    .B1(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__nand2_2 _20213_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][30] ),
    .Y(_07176_));
 sky130_fd_sc_hd__or2_2 _20214_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][30] ),
    .X(_07177_));
 sky130_fd_sc_hd__nand2_2 _20215_ (.A(_07176_),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2_2 _20216_ (.A(_07175_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__or2_2 _20217_ (.A(_07175_),
    .B(_07178_),
    .X(_07180_));
 sky130_fd_sc_hd__a32o_2 _20218_ (.A1(_11712_),
    .A2(_07179_),
    .A3(_07180_),
    .B1(\systolic_inst.acc_wires[6][30] ),
    .B2(_11258_),
    .X(_01584_));
 sky130_fd_sc_hd__xnor2_2 _20219_ (.A(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[6][31] ),
    .Y(_07181_));
 sky130_fd_sc_hd__a21oi_2 _20220_ (.A1(_07176_),
    .A2(_07180_),
    .B1(_07181_),
    .Y(_07182_));
 sky130_fd_sc_hd__a31o_2 _20221_ (.A1(_07176_),
    .A2(_07180_),
    .A3(_07181_),
    .B1(_11713_),
    .X(_07183_));
 sky130_fd_sc_hd__a2bb2o_2 _20222_ (.A1_N(_07183_),
    .A2_N(_07182_),
    .B1(\systolic_inst.acc_wires[6][31] ),
    .B2(_11258_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _20223_ (.A0(\systolic_inst.A_outs[5][0] ),
    .A1(\systolic_inst.A_outs[4][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _20224_ (.A0(\systolic_inst.A_outs[5][1] ),
    .A1(\systolic_inst.A_outs[4][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _20225_ (.A0(\systolic_inst.A_outs[5][2] ),
    .A1(\systolic_inst.A_outs[4][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _20226_ (.A0(\systolic_inst.A_outs[5][3] ),
    .A1(\systolic_inst.A_outs[4][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _20227_ (.A0(\systolic_inst.A_outs[5][4] ),
    .A1(\systolic_inst.A_outs[4][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _20228_ (.A0(\systolic_inst.A_outs[5][5] ),
    .A1(\systolic_inst.A_outs[4][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _20229_ (.A0(\systolic_inst.A_outs[5][6] ),
    .A1(\systolic_inst.A_outs[4][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _20230_ (.A0(\systolic_inst.A_outs[5][7] ),
    .A1(\systolic_inst.A_outs[4][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _20231_ (.A0(\systolic_inst.B_outs[4][0] ),
    .A1(\systolic_inst.B_outs[0][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _20232_ (.A0(\systolic_inst.B_outs[4][1] ),
    .A1(\systolic_inst.B_outs[0][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _20233_ (.A0(\systolic_inst.B_outs[4][2] ),
    .A1(\systolic_inst.B_outs[0][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _20234_ (.A0(\systolic_inst.B_outs[4][3] ),
    .A1(\systolic_inst.B_outs[0][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _20235_ (.A0(\systolic_inst.B_outs[4][4] ),
    .A1(\systolic_inst.B_outs[0][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _20236_ (.A0(\systolic_inst.B_outs[4][5] ),
    .A1(\systolic_inst.B_outs[0][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _20237_ (.A0(\systolic_inst.B_outs[4][6] ),
    .A1(\systolic_inst.B_outs[0][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_1 _20238_ (.A0(\systolic_inst.B_outs[4][7] ),
    .A1(\systolic_inst.B_outs[0][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01601_));
 sky130_fd_sc_hd__and3_2 _20239_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[5][0] ),
    .C(\systolic_inst.A_outs[5][0] ),
    .X(_07184_));
 sky130_fd_sc_hd__a21o_2 _20240_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[0] ),
    .B1(_07184_),
    .X(_01602_));
 sky130_fd_sc_hd__and4_2 _20241_ (.A(\systolic_inst.B_outs[5][0] ),
    .B(\systolic_inst.A_outs[5][0] ),
    .C(\systolic_inst.B_outs[5][1] ),
    .D(\systolic_inst.A_outs[5][1] ),
    .X(_07185_));
 sky130_fd_sc_hd__a22o_2 _20242_ (.A1(\systolic_inst.A_outs[5][0] ),
    .A2(\systolic_inst.B_outs[5][1] ),
    .B1(\systolic_inst.A_outs[5][1] ),
    .B2(\systolic_inst.B_outs[5][0] ),
    .X(_07186_));
 sky130_fd_sc_hd__nand2_2 _20243_ (.A(\systolic_inst.ce_local ),
    .B(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__a2bb2o_2 _20244_ (.A1_N(_07187_),
    .A2_N(_07185_),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01603_));
 sky130_fd_sc_hd__and2_2 _20245_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[2] ),
    .X(_07188_));
 sky130_fd_sc_hd__a22oi_2 _20246_ (.A1(\systolic_inst.B_outs[5][1] ),
    .A2(\systolic_inst.A_outs[5][1] ),
    .B1(\systolic_inst.A_outs[5][2] ),
    .B2(\systolic_inst.B_outs[5][0] ),
    .Y(_07189_));
 sky130_fd_sc_hd__and4_2 _20247_ (.A(\systolic_inst.B_outs[5][0] ),
    .B(\systolic_inst.B_outs[5][1] ),
    .C(\systolic_inst.A_outs[5][1] ),
    .D(\systolic_inst.A_outs[5][2] ),
    .X(_07190_));
 sky130_fd_sc_hd__or2_2 _20248_ (.A(_07189_),
    .B(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__or3b_2 _20249_ (.A(_07189_),
    .B(_07190_),
    .C_N(_07185_),
    .X(_07192_));
 sky130_fd_sc_hd__xnor2_2 _20250_ (.A(_07185_),
    .B(_07191_),
    .Y(_07193_));
 sky130_fd_sc_hd__nand3_2 _20251_ (.A(\systolic_inst.A_outs[5][0] ),
    .B(\systolic_inst.B_outs[5][2] ),
    .C(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__a21o_2 _20252_ (.A1(\systolic_inst.A_outs[5][0] ),
    .A2(\systolic_inst.B_outs[5][2] ),
    .B1(_07193_),
    .X(_07195_));
 sky130_fd_sc_hd__a31o_2 _20253_ (.A1(\systolic_inst.ce_local ),
    .A2(_07194_),
    .A3(_07195_),
    .B1(_07188_),
    .X(_01604_));
 sky130_fd_sc_hd__a22oi_2 _20254_ (.A1(\systolic_inst.A_outs[5][1] ),
    .A2(\systolic_inst.B_outs[5][2] ),
    .B1(\systolic_inst.B_outs[5][3] ),
    .B2(\systolic_inst.A_outs[5][0] ),
    .Y(_07196_));
 sky130_fd_sc_hd__and4_2 _20255_ (.A(\systolic_inst.A_outs[5][0] ),
    .B(\systolic_inst.A_outs[5][1] ),
    .C(\systolic_inst.B_outs[5][2] ),
    .D(\systolic_inst.B_outs[5][3] ),
    .X(_07197_));
 sky130_fd_sc_hd__nor2_2 _20256_ (.A(_07196_),
    .B(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__nand4_2 _20257_ (.A(\systolic_inst.B_outs[5][0] ),
    .B(\systolic_inst.B_outs[5][1] ),
    .C(\systolic_inst.A_outs[5][2] ),
    .D(\systolic_inst.A_outs[5][3] ),
    .Y(_07199_));
 sky130_fd_sc_hd__a22o_2 _20258_ (.A1(\systolic_inst.B_outs[5][1] ),
    .A2(\systolic_inst.A_outs[5][2] ),
    .B1(\systolic_inst.A_outs[5][3] ),
    .B2(\systolic_inst.B_outs[5][0] ),
    .X(_07200_));
 sky130_fd_sc_hd__nand3_2 _20259_ (.A(_07190_),
    .B(_07199_),
    .C(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__a21o_2 _20260_ (.A1(_07199_),
    .A2(_07200_),
    .B1(_07190_),
    .X(_07202_));
 sky130_fd_sc_hd__and2_2 _20261_ (.A(_07201_),
    .B(_07202_),
    .X(_07203_));
 sky130_fd_sc_hd__nand2_2 _20262_ (.A(_07198_),
    .B(_07203_),
    .Y(_07204_));
 sky130_fd_sc_hd__xnor2_2 _20263_ (.A(_07198_),
    .B(_07203_),
    .Y(_07205_));
 sky130_fd_sc_hd__and3_2 _20264_ (.A(_07192_),
    .B(_07194_),
    .C(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__a21oi_2 _20265_ (.A1(_07192_),
    .A2(_07194_),
    .B1(_07205_),
    .Y(_07207_));
 sky130_fd_sc_hd__nand2_2 _20266_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[3] ),
    .Y(_07208_));
 sky130_fd_sc_hd__o31ai_2 _20267_ (.A1(_11258_),
    .A2(_07206_),
    .A3(_07207_),
    .B1(_07208_),
    .Y(_01605_));
 sky130_fd_sc_hd__and2_2 _20268_ (.A(\systolic_inst.B_outs[5][2] ),
    .B(\systolic_inst.A_outs[5][2] ),
    .X(_07209_));
 sky130_fd_sc_hd__nand4_2 _20269_ (.A(\systolic_inst.A_outs[5][0] ),
    .B(\systolic_inst.A_outs[5][1] ),
    .C(\systolic_inst.B_outs[5][3] ),
    .D(\systolic_inst.B_outs[5][4] ),
    .Y(_07210_));
 sky130_fd_sc_hd__a22o_2 _20270_ (.A1(\systolic_inst.A_outs[5][1] ),
    .A2(\systolic_inst.B_outs[5][3] ),
    .B1(\systolic_inst.B_outs[5][4] ),
    .B2(\systolic_inst.A_outs[5][0] ),
    .X(_07211_));
 sky130_fd_sc_hd__nand2_2 _20271_ (.A(_07210_),
    .B(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__xnor2_2 _20272_ (.A(_07209_),
    .B(_07212_),
    .Y(_07213_));
 sky130_fd_sc_hd__a22o_2 _20273_ (.A1(\systolic_inst.B_outs[5][1] ),
    .A2(\systolic_inst.A_outs[5][3] ),
    .B1(\systolic_inst.A_outs[5][4] ),
    .B2(\systolic_inst.B_outs[5][0] ),
    .X(_07214_));
 sky130_fd_sc_hd__and3_2 _20274_ (.A(\systolic_inst.B_outs[5][0] ),
    .B(\systolic_inst.B_outs[5][1] ),
    .C(\systolic_inst.A_outs[5][3] ),
    .X(_07215_));
 sky130_fd_sc_hd__nand2_2 _20275_ (.A(\systolic_inst.A_outs[5][4] ),
    .B(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__and3_2 _20276_ (.A(_07197_),
    .B(_07214_),
    .C(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__a21oi_2 _20277_ (.A1(_07214_),
    .A2(_07216_),
    .B1(_07197_),
    .Y(_07218_));
 sky130_fd_sc_hd__o21ai_2 _20278_ (.A1(_07217_),
    .A2(_07218_),
    .B1(_07199_),
    .Y(_07219_));
 sky130_fd_sc_hd__nor3_2 _20279_ (.A(_07199_),
    .B(_07217_),
    .C(_07218_),
    .Y(_07220_));
 sky130_fd_sc_hd__or3_2 _20280_ (.A(_07199_),
    .B(_07217_),
    .C(_07218_),
    .X(_07221_));
 sky130_fd_sc_hd__and3_2 _20281_ (.A(_07213_),
    .B(_07219_),
    .C(_07221_),
    .X(_07222_));
 sky130_fd_sc_hd__a21oi_2 _20282_ (.A1(_07219_),
    .A2(_07221_),
    .B1(_07213_),
    .Y(_07223_));
 sky130_fd_sc_hd__a211o_2 _20283_ (.A1(_07201_),
    .A2(_07204_),
    .B1(_07222_),
    .C1(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__o211ai_2 _20284_ (.A1(_07222_),
    .A2(_07223_),
    .B1(_07201_),
    .C1(_07204_),
    .Y(_07225_));
 sky130_fd_sc_hd__a21oi_2 _20285_ (.A1(_07224_),
    .A2(_07225_),
    .B1(_07207_),
    .Y(_07226_));
 sky130_fd_sc_hd__a31o_2 _20286_ (.A1(_07207_),
    .A2(_07224_),
    .A3(_07225_),
    .B1(_11258_),
    .X(_07227_));
 sky130_fd_sc_hd__a2bb2o_2 _20287_ (.A1_N(_07227_),
    .A2_N(_07226_),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[4] ),
    .B2(_11258_),
    .X(_01606_));
 sky130_fd_sc_hd__a21bo_2 _20288_ (.A1(_07209_),
    .A2(_07211_),
    .B1_N(_07210_),
    .X(_07228_));
 sky130_fd_sc_hd__a22oi_2 _20289_ (.A1(\systolic_inst.B_outs[5][1] ),
    .A2(\systolic_inst.A_outs[5][4] ),
    .B1(\systolic_inst.A_outs[5][5] ),
    .B2(\systolic_inst.B_outs[5][0] ),
    .Y(_07229_));
 sky130_fd_sc_hd__and4_2 _20290_ (.A(\systolic_inst.B_outs[5][0] ),
    .B(\systolic_inst.B_outs[5][1] ),
    .C(\systolic_inst.A_outs[5][4] ),
    .D(\systolic_inst.A_outs[5][5] ),
    .X(_07230_));
 sky130_fd_sc_hd__nor2_2 _20291_ (.A(_07229_),
    .B(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__xor2_2 _20292_ (.A(_07228_),
    .B(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__xor2_2 _20293_ (.A(_07216_),
    .B(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__and2_2 _20294_ (.A(\systolic_inst.A_outs[5][0] ),
    .B(\systolic_inst.B_outs[5][5] ),
    .X(_07234_));
 sky130_fd_sc_hd__nand2_2 _20295_ (.A(\systolic_inst.A_outs[5][0] ),
    .B(\systolic_inst.B_outs[5][5] ),
    .Y(_07235_));
 sky130_fd_sc_hd__nand2_2 _20296_ (.A(\systolic_inst.B_outs[5][2] ),
    .B(\systolic_inst.A_outs[5][3] ),
    .Y(_07236_));
 sky130_fd_sc_hd__and4_2 _20297_ (.A(\systolic_inst.A_outs[5][1] ),
    .B(\systolic_inst.A_outs[5][2] ),
    .C(\systolic_inst.B_outs[5][3] ),
    .D(\systolic_inst.B_outs[5][4] ),
    .X(_07237_));
 sky130_fd_sc_hd__a22oi_2 _20298_ (.A1(\systolic_inst.A_outs[5][2] ),
    .A2(\systolic_inst.B_outs[5][3] ),
    .B1(\systolic_inst.B_outs[5][4] ),
    .B2(\systolic_inst.A_outs[5][1] ),
    .Y(_07238_));
 sky130_fd_sc_hd__or3_2 _20299_ (.A(_07236_),
    .B(_07237_),
    .C(_07238_),
    .X(_07239_));
 sky130_fd_sc_hd__o21ai_2 _20300_ (.A1(_07237_),
    .A2(_07238_),
    .B1(_07236_),
    .Y(_07240_));
 sky130_fd_sc_hd__and3_2 _20301_ (.A(_07234_),
    .B(_07239_),
    .C(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__a21oi_2 _20302_ (.A1(_07239_),
    .A2(_07240_),
    .B1(_07234_),
    .Y(_07242_));
 sky130_fd_sc_hd__or2_2 _20303_ (.A(_07241_),
    .B(_07242_),
    .X(_07243_));
 sky130_fd_sc_hd__nor2_2 _20304_ (.A(_07233_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__xor2_2 _20305_ (.A(_07233_),
    .B(_07243_),
    .X(_07245_));
 sky130_fd_sc_hd__and2_2 _20306_ (.A(_07222_),
    .B(_07245_),
    .X(_07246_));
 sky130_fd_sc_hd__xor2_2 _20307_ (.A(_07222_),
    .B(_07245_),
    .X(_07247_));
 sky130_fd_sc_hd__o21a_2 _20308_ (.A1(_07217_),
    .A2(_07220_),
    .B1(_07247_),
    .X(_07248_));
 sky130_fd_sc_hd__nor3_2 _20309_ (.A(_07217_),
    .B(_07220_),
    .C(_07247_),
    .Y(_07249_));
 sky130_fd_sc_hd__nor2_2 _20310_ (.A(_07248_),
    .B(_07249_),
    .Y(_07250_));
 sky130_fd_sc_hd__a21bo_2 _20311_ (.A1(_07207_),
    .A2(_07225_),
    .B1_N(_07224_),
    .X(_07251_));
 sky130_fd_sc_hd__nand2_2 _20312_ (.A(_07250_),
    .B(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__o21a_2 _20313_ (.A1(_07250_),
    .A2(_07251_),
    .B1(\systolic_inst.ce_local ),
    .X(_07253_));
 sky130_fd_sc_hd__a22o_2 _20314_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[5] ),
    .B1(_07252_),
    .B2(_07253_),
    .X(_01607_));
 sky130_fd_sc_hd__a32o_2 _20315_ (.A1(\systolic_inst.A_outs[5][4] ),
    .A2(_07215_),
    .A3(_07232_),
    .B1(_07231_),
    .B2(_07228_),
    .X(_07254_));
 sky130_fd_sc_hd__o21bai_2 _20316_ (.A1(_07236_),
    .A2(_07238_),
    .B1_N(_07237_),
    .Y(_07255_));
 sky130_fd_sc_hd__a22oi_2 _20317_ (.A1(\systolic_inst.B_outs[5][1] ),
    .A2(\systolic_inst.A_outs[5][5] ),
    .B1(\systolic_inst.A_outs[5][6] ),
    .B2(\systolic_inst.B_outs[5][0] ),
    .Y(_07256_));
 sky130_fd_sc_hd__and4_2 _20318_ (.A(\systolic_inst.B_outs[5][0] ),
    .B(\systolic_inst.B_outs[5][1] ),
    .C(\systolic_inst.A_outs[5][5] ),
    .D(\systolic_inst.A_outs[5][6] ),
    .X(_07257_));
 sky130_fd_sc_hd__or2_2 _20319_ (.A(_07256_),
    .B(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__nand2b_2 _20320_ (.A_N(_07258_),
    .B(_07255_),
    .Y(_07259_));
 sky130_fd_sc_hd__xnor2_2 _20321_ (.A(_07255_),
    .B(_07258_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_2 _20322_ (.A(_07230_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__xor2_2 _20323_ (.A(_07230_),
    .B(_07260_),
    .X(_07262_));
 sky130_fd_sc_hd__nand4_2 _20324_ (.A(\systolic_inst.A_outs[5][2] ),
    .B(\systolic_inst.B_outs[5][3] ),
    .C(\systolic_inst.A_outs[5][3] ),
    .D(\systolic_inst.B_outs[5][4] ),
    .Y(_07263_));
 sky130_fd_sc_hd__a22o_2 _20325_ (.A1(\systolic_inst.B_outs[5][3] ),
    .A2(\systolic_inst.A_outs[5][3] ),
    .B1(\systolic_inst.B_outs[5][4] ),
    .B2(\systolic_inst.A_outs[5][2] ),
    .X(_07264_));
 sky130_fd_sc_hd__nand4_2 _20326_ (.A(\systolic_inst.B_outs[5][2] ),
    .B(\systolic_inst.A_outs[5][4] ),
    .C(_07263_),
    .D(_07264_),
    .Y(_07265_));
 sky130_fd_sc_hd__a22o_2 _20327_ (.A1(\systolic_inst.B_outs[5][2] ),
    .A2(\systolic_inst.A_outs[5][4] ),
    .B1(_07263_),
    .B2(_07264_),
    .X(_07266_));
 sky130_fd_sc_hd__nand2_2 _20328_ (.A(\systolic_inst.A_outs[5][1] ),
    .B(\systolic_inst.B_outs[5][6] ),
    .Y(_07267_));
 sky130_fd_sc_hd__a22o_2 _20329_ (.A1(\systolic_inst.A_outs[5][1] ),
    .A2(\systolic_inst.B_outs[5][5] ),
    .B1(\systolic_inst.B_outs[5][6] ),
    .B2(\systolic_inst.A_outs[5][0] ),
    .X(_07268_));
 sky130_fd_sc_hd__o21a_2 _20330_ (.A1(_07235_),
    .A2(_07267_),
    .B1(_07268_),
    .X(_07269_));
 sky130_fd_sc_hd__and3_2 _20331_ (.A(_07265_),
    .B(_07266_),
    .C(_07269_),
    .X(_07270_));
 sky130_fd_sc_hd__nand3_2 _20332_ (.A(_07265_),
    .B(_07266_),
    .C(_07269_),
    .Y(_07271_));
 sky130_fd_sc_hd__a21o_2 _20333_ (.A1(_07265_),
    .A2(_07266_),
    .B1(_07269_),
    .X(_07272_));
 sky130_fd_sc_hd__nand3_2 _20334_ (.A(_07241_),
    .B(_07271_),
    .C(_07272_),
    .Y(_07273_));
 sky130_fd_sc_hd__a21o_2 _20335_ (.A1(_07271_),
    .A2(_07272_),
    .B1(_07241_),
    .X(_07274_));
 sky130_fd_sc_hd__nand3_2 _20336_ (.A(_07262_),
    .B(_07273_),
    .C(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__a21o_2 _20337_ (.A1(_07273_),
    .A2(_07274_),
    .B1(_07262_),
    .X(_07276_));
 sky130_fd_sc_hd__nand3_2 _20338_ (.A(_07244_),
    .B(_07275_),
    .C(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__a21o_2 _20339_ (.A1(_07275_),
    .A2(_07276_),
    .B1(_07244_),
    .X(_07278_));
 sky130_fd_sc_hd__nand3_2 _20340_ (.A(_07254_),
    .B(_07277_),
    .C(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__a21o_2 _20341_ (.A1(_07277_),
    .A2(_07278_),
    .B1(_07254_),
    .X(_07280_));
 sky130_fd_sc_hd__o211a_2 _20342_ (.A1(_07246_),
    .A2(_07248_),
    .B1(_07279_),
    .C1(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__a211o_2 _20343_ (.A1(_07279_),
    .A2(_07280_),
    .B1(_07246_),
    .C1(_07248_),
    .X(_07282_));
 sky130_fd_sc_hd__and2b_2 _20344_ (.A_N(_07281_),
    .B(_07282_),
    .X(_07283_));
 sky130_fd_sc_hd__xnor2_2 _20345_ (.A(_07252_),
    .B(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__mux2_1 _20346_ (.A0(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[6] ),
    .A1(_07284_),
    .S(\systolic_inst.ce_local ),
    .X(_01608_));
 sky130_fd_sc_hd__nand2_2 _20347_ (.A(_07263_),
    .B(_07265_),
    .Y(_07285_));
 sky130_fd_sc_hd__nand2_2 _20348_ (.A(\systolic_inst.B_outs[5][0] ),
    .B(\systolic_inst.A_outs[5][7] ),
    .Y(_07286_));
 sky130_fd_sc_hd__nand2_2 _20349_ (.A(\systolic_inst.B_outs[5][2] ),
    .B(\systolic_inst.A_outs[5][6] ),
    .Y(_07287_));
 sky130_fd_sc_hd__and4_2 _20350_ (.A(\systolic_inst.B_outs[5][1] ),
    .B(\systolic_inst.B_outs[5][2] ),
    .C(\systolic_inst.A_outs[5][5] ),
    .D(\systolic_inst.A_outs[5][6] ),
    .X(_07288_));
 sky130_fd_sc_hd__a22o_2 _20351_ (.A1(\systolic_inst.B_outs[5][2] ),
    .A2(\systolic_inst.A_outs[5][5] ),
    .B1(\systolic_inst.A_outs[5][6] ),
    .B2(\systolic_inst.B_outs[5][1] ),
    .X(_07289_));
 sky130_fd_sc_hd__and2b_2 _20352_ (.A_N(_07288_),
    .B(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__xnor2_2 _20353_ (.A(_07286_),
    .B(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__xor2_2 _20354_ (.A(_07285_),
    .B(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__and2_2 _20355_ (.A(_07257_),
    .B(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__xnor2_2 _20356_ (.A(_07257_),
    .B(_07292_),
    .Y(_07294_));
 sky130_fd_sc_hd__nand2_2 _20357_ (.A(\systolic_inst.B_outs[5][3] ),
    .B(\systolic_inst.A_outs[5][4] ),
    .Y(_07295_));
 sky130_fd_sc_hd__nand2_2 _20358_ (.A(\systolic_inst.A_outs[5][3] ),
    .B(\systolic_inst.B_outs[5][5] ),
    .Y(_07296_));
 sky130_fd_sc_hd__and4_2 _20359_ (.A(\systolic_inst.A_outs[5][2] ),
    .B(\systolic_inst.A_outs[5][3] ),
    .C(\systolic_inst.B_outs[5][4] ),
    .D(\systolic_inst.B_outs[5][5] ),
    .X(_07297_));
 sky130_fd_sc_hd__a22o_2 _20360_ (.A1(\systolic_inst.A_outs[5][3] ),
    .A2(\systolic_inst.B_outs[5][4] ),
    .B1(\systolic_inst.B_outs[5][5] ),
    .B2(\systolic_inst.A_outs[5][2] ),
    .X(_07298_));
 sky130_fd_sc_hd__and2b_2 _20361_ (.A_N(_07297_),
    .B(_07298_),
    .X(_07299_));
 sky130_fd_sc_hd__xnor2_2 _20362_ (.A(_07295_),
    .B(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__o211ai_2 _20363_ (.A1(\systolic_inst.B_outs[5][5] ),
    .A2(_07267_),
    .B1(\systolic_inst.B_outs[5][7] ),
    .C1(\systolic_inst.A_outs[5][0] ),
    .Y(_07301_));
 sky130_fd_sc_hd__a211o_2 _20364_ (.A1(\systolic_inst.A_outs[5][0] ),
    .A2(\systolic_inst.B_outs[5][7] ),
    .B1(_07234_),
    .C1(_07267_),
    .X(_07302_));
 sky130_fd_sc_hd__nand2_2 _20365_ (.A(_07301_),
    .B(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand2_2 _20366_ (.A(_07300_),
    .B(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__xor2_2 _20367_ (.A(_07300_),
    .B(_07303_),
    .X(_07305_));
 sky130_fd_sc_hd__xnor2_2 _20368_ (.A(_07270_),
    .B(_07305_),
    .Y(_07306_));
 sky130_fd_sc_hd__or2_2 _20369_ (.A(_07294_),
    .B(_07306_),
    .X(_07307_));
 sky130_fd_sc_hd__nand2_2 _20370_ (.A(_07294_),
    .B(_07306_),
    .Y(_07308_));
 sky130_fd_sc_hd__nand2_2 _20371_ (.A(_07273_),
    .B(_07275_),
    .Y(_07309_));
 sky130_fd_sc_hd__and3_2 _20372_ (.A(_07307_),
    .B(_07308_),
    .C(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__a21oi_2 _20373_ (.A1(_07307_),
    .A2(_07308_),
    .B1(_07309_),
    .Y(_07311_));
 sky130_fd_sc_hd__a211oi_2 _20374_ (.A1(_07259_),
    .A2(_07261_),
    .B1(_07310_),
    .C1(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__o211a_2 _20375_ (.A1(_07310_),
    .A2(_07311_),
    .B1(_07259_),
    .C1(_07261_),
    .X(_07313_));
 sky130_fd_sc_hd__a211oi_2 _20376_ (.A1(_07277_),
    .A2(_07279_),
    .B1(_07312_),
    .C1(_07313_),
    .Y(_07314_));
 sky130_fd_sc_hd__o211ai_2 _20377_ (.A1(_07312_),
    .A2(_07313_),
    .B1(_07277_),
    .C1(_07279_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand2b_2 _20378_ (.A_N(_07314_),
    .B(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__a31o_2 _20379_ (.A1(_07250_),
    .A2(_07251_),
    .A3(_07282_),
    .B1(_07281_),
    .X(_07317_));
 sky130_fd_sc_hd__xnor2_2 _20380_ (.A(_07316_),
    .B(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__mux2_1 _20381_ (.A0(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[7] ),
    .A1(_07318_),
    .S(\systolic_inst.ce_local ),
    .X(_01609_));
 sky130_fd_sc_hd__a21oi_2 _20382_ (.A1(_07285_),
    .A2(_07291_),
    .B1(_07293_),
    .Y(_07319_));
 sky130_fd_sc_hd__a31o_2 _20383_ (.A1(\systolic_inst.B_outs[5][0] ),
    .A2(\systolic_inst.A_outs[5][7] ),
    .A3(_07289_),
    .B1(_07288_),
    .X(_07320_));
 sky130_fd_sc_hd__a31o_2 _20384_ (.A1(\systolic_inst.B_outs[5][3] ),
    .A2(\systolic_inst.A_outs[5][4] ),
    .A3(_07298_),
    .B1(_07297_),
    .X(_07321_));
 sky130_fd_sc_hd__o21ai_2 _20385_ (.A1(\systolic_inst.B_outs[5][0] ),
    .A2(\systolic_inst.B_outs[5][1] ),
    .B1(\systolic_inst.A_outs[5][7] ),
    .Y(_07322_));
 sky130_fd_sc_hd__o21a_2 _20386_ (.A1(\systolic_inst.B_outs[5][0] ),
    .A2(\systolic_inst.B_outs[5][1] ),
    .B1(\systolic_inst.A_outs[5][7] ),
    .X(_07323_));
 sky130_fd_sc_hd__a21o_2 _20387_ (.A1(\systolic_inst.B_outs[5][0] ),
    .A2(\systolic_inst.B_outs[5][1] ),
    .B1(_07322_),
    .X(_07324_));
 sky130_fd_sc_hd__and2b_2 _20388_ (.A_N(_07324_),
    .B(_07321_),
    .X(_07325_));
 sky130_fd_sc_hd__xnor2_2 _20389_ (.A(_07321_),
    .B(_07324_),
    .Y(_07326_));
 sky130_fd_sc_hd__xnor2_2 _20390_ (.A(_07320_),
    .B(_07326_),
    .Y(_07327_));
 sky130_fd_sc_hd__and4_2 _20391_ (.A(\systolic_inst.B_outs[5][3] ),
    .B(\systolic_inst.B_outs[5][4] ),
    .C(\systolic_inst.A_outs[5][4] ),
    .D(\systolic_inst.A_outs[5][5] ),
    .X(_07328_));
 sky130_fd_sc_hd__a22oi_2 _20392_ (.A1(\systolic_inst.B_outs[5][4] ),
    .A2(\systolic_inst.A_outs[5][4] ),
    .B1(\systolic_inst.A_outs[5][5] ),
    .B2(\systolic_inst.B_outs[5][3] ),
    .Y(_07329_));
 sky130_fd_sc_hd__nor2_2 _20393_ (.A(_07328_),
    .B(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__xnor2_2 _20394_ (.A(_07287_),
    .B(_07330_),
    .Y(_07331_));
 sky130_fd_sc_hd__inv_2 _20395_ (.A(_07331_),
    .Y(_07332_));
 sky130_fd_sc_hd__and2b_2 _20396_ (.A_N(\systolic_inst.A_outs[5][1] ),
    .B(\systolic_inst.B_outs[5][7] ),
    .X(_07333_));
 sky130_fd_sc_hd__nand2_2 _20397_ (.A(\systolic_inst.A_outs[5][2] ),
    .B(\systolic_inst.B_outs[5][6] ),
    .Y(_07334_));
 sky130_fd_sc_hd__and3_2 _20398_ (.A(\systolic_inst.A_outs[5][2] ),
    .B(\systolic_inst.B_outs[5][6] ),
    .C(_07333_),
    .X(_07335_));
 sky130_fd_sc_hd__xnor2_2 _20399_ (.A(_07333_),
    .B(_07334_),
    .Y(_07336_));
 sky130_fd_sc_hd__xnor2_2 _20400_ (.A(_07296_),
    .B(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__nand2_2 _20401_ (.A(\systolic_inst.A_outs[5][0] ),
    .B(_07267_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand2_2 _20402_ (.A(\systolic_inst.B_outs[5][7] ),
    .B(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__and3_2 _20403_ (.A(\systolic_inst.B_outs[5][7] ),
    .B(_07337_),
    .C(_07338_),
    .X(_07340_));
 sky130_fd_sc_hd__xor2_2 _20404_ (.A(_07337_),
    .B(_07339_),
    .X(_07341_));
 sky130_fd_sc_hd__xnor2_2 _20405_ (.A(_07332_),
    .B(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__o31a_2 _20406_ (.A1(\systolic_inst.B_outs[5][7] ),
    .A2(_07235_),
    .A3(_07267_),
    .B1(_07304_),
    .X(_07343_));
 sky130_fd_sc_hd__or2_2 _20407_ (.A(_07342_),
    .B(_07343_),
    .X(_07344_));
 sky130_fd_sc_hd__xnor2_2 _20408_ (.A(_07342_),
    .B(_07343_),
    .Y(_07345_));
 sky130_fd_sc_hd__xnor2_2 _20409_ (.A(_07327_),
    .B(_07345_),
    .Y(_07346_));
 sky130_fd_sc_hd__a21bo_2 _20410_ (.A1(_07270_),
    .A2(_07305_),
    .B1_N(_07307_),
    .X(_07347_));
 sky130_fd_sc_hd__nand2b_2 _20411_ (.A_N(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__xnor2_2 _20412_ (.A(_07346_),
    .B(_07347_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand2b_2 _20413_ (.A_N(_07319_),
    .B(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__xnor2_2 _20414_ (.A(_07319_),
    .B(_07349_),
    .Y(_07351_));
 sky130_fd_sc_hd__nor2_2 _20415_ (.A(_07310_),
    .B(_07312_),
    .Y(_07352_));
 sky130_fd_sc_hd__nand2b_2 _20416_ (.A_N(_07352_),
    .B(_07351_),
    .Y(_07353_));
 sky130_fd_sc_hd__xnor2_2 _20417_ (.A(_07351_),
    .B(_07352_),
    .Y(_07354_));
 sky130_fd_sc_hd__a21oi_2 _20418_ (.A1(_07315_),
    .A2(_07317_),
    .B1(_07314_),
    .Y(_07355_));
 sky130_fd_sc_hd__nand2b_2 _20419_ (.A_N(_07355_),
    .B(_07354_),
    .Y(_07356_));
 sky130_fd_sc_hd__nand2b_2 _20420_ (.A_N(_07354_),
    .B(_07355_),
    .Y(_07357_));
 sky130_fd_sc_hd__and2_2 _20421_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[8] ),
    .X(_07358_));
 sky130_fd_sc_hd__a31o_2 _20422_ (.A1(\systolic_inst.ce_local ),
    .A2(_07356_),
    .A3(_07357_),
    .B1(_07358_),
    .X(_01610_));
 sky130_fd_sc_hd__a21o_2 _20423_ (.A1(_07320_),
    .A2(_07326_),
    .B1(_07325_),
    .X(_07359_));
 sky130_fd_sc_hd__o21ba_2 _20424_ (.A1(_07287_),
    .A2(_07329_),
    .B1_N(_07328_),
    .X(_07360_));
 sky130_fd_sc_hd__nor2_2 _20425_ (.A(_07322_),
    .B(_07360_),
    .Y(_07361_));
 sky130_fd_sc_hd__and2_2 _20426_ (.A(_07322_),
    .B(_07360_),
    .X(_07362_));
 sky130_fd_sc_hd__or2_2 _20427_ (.A(_07361_),
    .B(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__nand2_2 _20428_ (.A(\systolic_inst.B_outs[5][2] ),
    .B(\systolic_inst.A_outs[5][7] ),
    .Y(_07364_));
 sky130_fd_sc_hd__a22oi_2 _20429_ (.A1(\systolic_inst.B_outs[5][4] ),
    .A2(\systolic_inst.A_outs[5][5] ),
    .B1(\systolic_inst.A_outs[5][6] ),
    .B2(\systolic_inst.B_outs[5][3] ),
    .Y(_07365_));
 sky130_fd_sc_hd__and4_2 _20430_ (.A(\systolic_inst.B_outs[5][3] ),
    .B(\systolic_inst.B_outs[5][4] ),
    .C(\systolic_inst.A_outs[5][5] ),
    .D(\systolic_inst.A_outs[5][6] ),
    .X(_07366_));
 sky130_fd_sc_hd__nor2_2 _20431_ (.A(_07365_),
    .B(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__xnor2_2 _20432_ (.A(_07364_),
    .B(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__nand2_2 _20433_ (.A(\systolic_inst.A_outs[5][4] ),
    .B(\systolic_inst.B_outs[5][5] ),
    .Y(_07369_));
 sky130_fd_sc_hd__and4b_2 _20434_ (.A_N(\systolic_inst.A_outs[5][2] ),
    .B(\systolic_inst.A_outs[5][3] ),
    .C(\systolic_inst.B_outs[5][6] ),
    .D(\systolic_inst.B_outs[5][7] ),
    .X(_07370_));
 sky130_fd_sc_hd__o2bb2a_2 _20435_ (.A1_N(\systolic_inst.A_outs[5][3] ),
    .A2_N(\systolic_inst.B_outs[5][6] ),
    .B1(_11276_),
    .B2(\systolic_inst.A_outs[5][2] ),
    .X(_07371_));
 sky130_fd_sc_hd__nor2_2 _20436_ (.A(_07370_),
    .B(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__xnor2_2 _20437_ (.A(_07369_),
    .B(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__a31oi_2 _20438_ (.A1(\systolic_inst.A_outs[5][3] ),
    .A2(\systolic_inst.B_outs[5][5] ),
    .A3(_07336_),
    .B1(_07335_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand2b_2 _20439_ (.A_N(_07374_),
    .B(_07373_),
    .Y(_07375_));
 sky130_fd_sc_hd__xnor2_2 _20440_ (.A(_07373_),
    .B(_07374_),
    .Y(_07376_));
 sky130_fd_sc_hd__xnor2_2 _20441_ (.A(_07368_),
    .B(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__o21ba_2 _20442_ (.A1(_07332_),
    .A2(_07341_),
    .B1_N(_07340_),
    .X(_07378_));
 sky130_fd_sc_hd__xnor2_2 _20443_ (.A(_07377_),
    .B(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__or2_2 _20444_ (.A(_07363_),
    .B(_07379_),
    .X(_07380_));
 sky130_fd_sc_hd__nand2_2 _20445_ (.A(_07363_),
    .B(_07379_),
    .Y(_07381_));
 sky130_fd_sc_hd__and2_2 _20446_ (.A(_07380_),
    .B(_07381_),
    .X(_07382_));
 sky130_fd_sc_hd__o21a_2 _20447_ (.A1(_07327_),
    .A2(_07345_),
    .B1(_07344_),
    .X(_07383_));
 sky130_fd_sc_hd__nand2b_2 _20448_ (.A_N(_07383_),
    .B(_07382_),
    .Y(_07384_));
 sky130_fd_sc_hd__xnor2_2 _20449_ (.A(_07382_),
    .B(_07383_),
    .Y(_07385_));
 sky130_fd_sc_hd__xnor2_2 _20450_ (.A(_07359_),
    .B(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__a21o_2 _20451_ (.A1(_07348_),
    .A2(_07350_),
    .B1(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__nand3_2 _20452_ (.A(_07348_),
    .B(_07350_),
    .C(_07386_),
    .Y(_07388_));
 sky130_fd_sc_hd__nand2_2 _20453_ (.A(_07353_),
    .B(_07356_),
    .Y(_07389_));
 sky130_fd_sc_hd__and3_2 _20454_ (.A(_07387_),
    .B(_07388_),
    .C(_07389_),
    .X(_07390_));
 sky130_fd_sc_hd__a21oi_2 _20455_ (.A1(_07387_),
    .A2(_07388_),
    .B1(_07389_),
    .Y(_07391_));
 sky130_fd_sc_hd__nor2_2 _20456_ (.A(_07390_),
    .B(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__mux2_1 _20457_ (.A0(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[9] ),
    .A1(_07392_),
    .S(\systolic_inst.ce_local ),
    .X(_01611_));
 sky130_fd_sc_hd__o21ba_2 _20458_ (.A1(_07364_),
    .A2(_07365_),
    .B1_N(_07366_),
    .X(_07393_));
 sky130_fd_sc_hd__nor2_2 _20459_ (.A(_07322_),
    .B(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__and2_2 _20460_ (.A(_07322_),
    .B(_07393_),
    .X(_07395_));
 sky130_fd_sc_hd__or2_2 _20461_ (.A(_07394_),
    .B(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__a22o_2 _20462_ (.A1(\systolic_inst.B_outs[5][4] ),
    .A2(\systolic_inst.A_outs[5][6] ),
    .B1(\systolic_inst.A_outs[5][7] ),
    .B2(\systolic_inst.B_outs[5][3] ),
    .X(_07397_));
 sky130_fd_sc_hd__and3_2 _20463_ (.A(\systolic_inst.B_outs[5][3] ),
    .B(\systolic_inst.B_outs[5][4] ),
    .C(\systolic_inst.A_outs[5][7] ),
    .X(_07398_));
 sky130_fd_sc_hd__a21bo_2 _20464_ (.A1(\systolic_inst.A_outs[5][6] ),
    .A2(_07398_),
    .B1_N(_07397_),
    .X(_07399_));
 sky130_fd_sc_hd__xor2_2 _20465_ (.A(_07364_),
    .B(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__nand2_2 _20466_ (.A(\systolic_inst.B_outs[5][5] ),
    .B(\systolic_inst.A_outs[5][5] ),
    .Y(_07401_));
 sky130_fd_sc_hd__and4b_2 _20467_ (.A_N(\systolic_inst.A_outs[5][3] ),
    .B(\systolic_inst.A_outs[5][4] ),
    .C(\systolic_inst.B_outs[5][6] ),
    .D(\systolic_inst.B_outs[5][7] ),
    .X(_07402_));
 sky130_fd_sc_hd__o2bb2a_2 _20468_ (.A1_N(\systolic_inst.A_outs[5][4] ),
    .A2_N(\systolic_inst.B_outs[5][6] ),
    .B1(_11276_),
    .B2(\systolic_inst.A_outs[5][3] ),
    .X(_07403_));
 sky130_fd_sc_hd__nor2_2 _20469_ (.A(_07402_),
    .B(_07403_),
    .Y(_07404_));
 sky130_fd_sc_hd__xnor2_2 _20470_ (.A(_07401_),
    .B(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__o21ba_2 _20471_ (.A1(_07369_),
    .A2(_07371_),
    .B1_N(_07370_),
    .X(_07406_));
 sky130_fd_sc_hd__nand2b_2 _20472_ (.A_N(_07406_),
    .B(_07405_),
    .Y(_07407_));
 sky130_fd_sc_hd__xnor2_2 _20473_ (.A(_07405_),
    .B(_07406_),
    .Y(_07408_));
 sky130_fd_sc_hd__nand2_2 _20474_ (.A(_07400_),
    .B(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__or2_2 _20475_ (.A(_07400_),
    .B(_07408_),
    .X(_07410_));
 sky130_fd_sc_hd__nand2_2 _20476_ (.A(_07409_),
    .B(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__a21bo_2 _20477_ (.A1(_07368_),
    .A2(_07376_),
    .B1_N(_07375_),
    .X(_07412_));
 sky130_fd_sc_hd__nand2b_2 _20478_ (.A_N(_07411_),
    .B(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__xor2_2 _20479_ (.A(_07411_),
    .B(_07412_),
    .X(_07414_));
 sky130_fd_sc_hd__xor2_2 _20480_ (.A(_07396_),
    .B(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__o21a_2 _20481_ (.A1(_07377_),
    .A2(_07378_),
    .B1(_07380_),
    .X(_07416_));
 sky130_fd_sc_hd__nand2b_2 _20482_ (.A_N(_07416_),
    .B(_07415_),
    .Y(_07417_));
 sky130_fd_sc_hd__xnor2_2 _20483_ (.A(_07415_),
    .B(_07416_),
    .Y(_07418_));
 sky130_fd_sc_hd__nand2_2 _20484_ (.A(_07361_),
    .B(_07418_),
    .Y(_07419_));
 sky130_fd_sc_hd__xnor2_2 _20485_ (.A(_07361_),
    .B(_07418_),
    .Y(_07420_));
 sky130_fd_sc_hd__a21boi_2 _20486_ (.A1(_07359_),
    .A2(_07385_),
    .B1_N(_07384_),
    .Y(_07421_));
 sky130_fd_sc_hd__or2_2 _20487_ (.A(_07420_),
    .B(_07421_),
    .X(_07422_));
 sky130_fd_sc_hd__nand2_2 _20488_ (.A(_07420_),
    .B(_07421_),
    .Y(_07423_));
 sky130_fd_sc_hd__nand2_2 _20489_ (.A(_07422_),
    .B(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__nand2_2 _20490_ (.A(_07388_),
    .B(_07389_),
    .Y(_07425_));
 sky130_fd_sc_hd__and3_2 _20491_ (.A(_07387_),
    .B(_07424_),
    .C(_07425_),
    .X(_07426_));
 sky130_fd_sc_hd__a21o_2 _20492_ (.A1(_07387_),
    .A2(_07425_),
    .B1(_07424_),
    .X(_07427_));
 sky130_fd_sc_hd__nand2_2 _20493_ (.A(\systolic_inst.ce_local ),
    .B(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__a2bb2o_2 _20494_ (.A1_N(_07428_),
    .A2_N(_07426_),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[10] ),
    .B2(_11258_),
    .X(_01612_));
 sky130_fd_sc_hd__o2bb2a_2 _20495_ (.A1_N(\systolic_inst.A_outs[5][6] ),
    .A2_N(_07398_),
    .B1(_07399_),
    .B2(_07364_),
    .X(_07429_));
 sky130_fd_sc_hd__nor2_2 _20496_ (.A(_07322_),
    .B(_07429_),
    .Y(_07430_));
 sky130_fd_sc_hd__and2_2 _20497_ (.A(_07322_),
    .B(_07429_),
    .X(_07431_));
 sky130_fd_sc_hd__or2_2 _20498_ (.A(_07430_),
    .B(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__or2_2 _20499_ (.A(\systolic_inst.B_outs[5][3] ),
    .B(\systolic_inst.B_outs[5][4] ),
    .X(_07433_));
 sky130_fd_sc_hd__and3b_2 _20500_ (.A_N(_07398_),
    .B(_07433_),
    .C(\systolic_inst.A_outs[5][7] ),
    .X(_07434_));
 sky130_fd_sc_hd__xnor2_2 _20501_ (.A(_07364_),
    .B(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__nand2_2 _20502_ (.A(\systolic_inst.B_outs[5][5] ),
    .B(\systolic_inst.A_outs[5][6] ),
    .Y(_07436_));
 sky130_fd_sc_hd__and4b_2 _20503_ (.A_N(\systolic_inst.A_outs[5][4] ),
    .B(\systolic_inst.A_outs[5][5] ),
    .C(\systolic_inst.B_outs[5][6] ),
    .D(\systolic_inst.B_outs[5][7] ),
    .X(_07437_));
 sky130_fd_sc_hd__o2bb2a_2 _20504_ (.A1_N(\systolic_inst.A_outs[5][5] ),
    .A2_N(\systolic_inst.B_outs[5][6] ),
    .B1(_11276_),
    .B2(\systolic_inst.A_outs[5][4] ),
    .X(_07438_));
 sky130_fd_sc_hd__or2_2 _20505_ (.A(_07437_),
    .B(_07438_),
    .X(_07439_));
 sky130_fd_sc_hd__xor2_2 _20506_ (.A(_07436_),
    .B(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__o21ba_2 _20507_ (.A1(_07401_),
    .A2(_07403_),
    .B1_N(_07402_),
    .X(_07441_));
 sky130_fd_sc_hd__nand2b_2 _20508_ (.A_N(_07441_),
    .B(_07440_),
    .Y(_07442_));
 sky130_fd_sc_hd__xnor2_2 _20509_ (.A(_07440_),
    .B(_07441_),
    .Y(_07443_));
 sky130_fd_sc_hd__nand2_2 _20510_ (.A(_07435_),
    .B(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__xnor2_2 _20511_ (.A(_07435_),
    .B(_07443_),
    .Y(_07445_));
 sky130_fd_sc_hd__a21o_2 _20512_ (.A1(_07407_),
    .A2(_07409_),
    .B1(_07445_),
    .X(_07446_));
 sky130_fd_sc_hd__nand3_2 _20513_ (.A(_07407_),
    .B(_07409_),
    .C(_07445_),
    .Y(_07447_));
 sky130_fd_sc_hd__nand2_2 _20514_ (.A(_07446_),
    .B(_07447_),
    .Y(_07448_));
 sky130_fd_sc_hd__xor2_2 _20515_ (.A(_07432_),
    .B(_07448_),
    .X(_07449_));
 sky130_fd_sc_hd__o21a_2 _20516_ (.A1(_07396_),
    .A2(_07414_),
    .B1(_07413_),
    .X(_07450_));
 sky130_fd_sc_hd__and2b_2 _20517_ (.A_N(_07450_),
    .B(_07449_),
    .X(_07451_));
 sky130_fd_sc_hd__and2b_2 _20518_ (.A_N(_07449_),
    .B(_07450_),
    .X(_07452_));
 sky130_fd_sc_hd__nor2_2 _20519_ (.A(_07451_),
    .B(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__xnor2_2 _20520_ (.A(_07394_),
    .B(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__nand3_2 _20521_ (.A(_07417_),
    .B(_07419_),
    .C(_07454_),
    .Y(_07455_));
 sky130_fd_sc_hd__inv_2 _20522_ (.A(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__a21o_2 _20523_ (.A1(_07417_),
    .A2(_07419_),
    .B1(_07454_),
    .X(_07457_));
 sky130_fd_sc_hd__nand2_2 _20524_ (.A(_07455_),
    .B(_07457_),
    .Y(_07458_));
 sky130_fd_sc_hd__a21oi_2 _20525_ (.A1(_07422_),
    .A2(_07427_),
    .B1(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__a31o_2 _20526_ (.A1(_07422_),
    .A2(_07427_),
    .A3(_07458_),
    .B1(_11258_),
    .X(_07460_));
 sky130_fd_sc_hd__a2bb2o_2 _20527_ (.A1_N(_07460_),
    .A2_N(_07459_),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[11] ),
    .B2(_11258_),
    .X(_01613_));
 sky130_fd_sc_hd__a31o_2 _20528_ (.A1(\systolic_inst.B_outs[5][2] ),
    .A2(\systolic_inst.A_outs[5][7] ),
    .A3(_07433_),
    .B1(_07398_),
    .X(_07461_));
 sky130_fd_sc_hd__or2_2 _20529_ (.A(_07323_),
    .B(_07461_),
    .X(_07462_));
 sky130_fd_sc_hd__nand2_2 _20530_ (.A(_07323_),
    .B(_07461_),
    .Y(_07463_));
 sky130_fd_sc_hd__nand2_2 _20531_ (.A(_07462_),
    .B(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__inv_2 _20532_ (.A(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__o2bb2a_2 _20533_ (.A1_N(\systolic_inst.B_outs[5][6] ),
    .A2_N(\systolic_inst.A_outs[5][6] ),
    .B1(_11276_),
    .B2(\systolic_inst.A_outs[5][5] ),
    .X(_07466_));
 sky130_fd_sc_hd__and4b_2 _20534_ (.A_N(\systolic_inst.A_outs[5][5] ),
    .B(\systolic_inst.B_outs[5][6] ),
    .C(\systolic_inst.A_outs[5][6] ),
    .D(\systolic_inst.B_outs[5][7] ),
    .X(_07467_));
 sky130_fd_sc_hd__nor2_2 _20535_ (.A(_07466_),
    .B(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__nand2_2 _20536_ (.A(\systolic_inst.B_outs[5][5] ),
    .B(\systolic_inst.A_outs[5][7] ),
    .Y(_07469_));
 sky130_fd_sc_hd__and3_2 _20537_ (.A(\systolic_inst.B_outs[5][5] ),
    .B(\systolic_inst.A_outs[5][7] ),
    .C(_07468_),
    .X(_07470_));
 sky130_fd_sc_hd__xnor2_2 _20538_ (.A(_07468_),
    .B(_07469_),
    .Y(_07471_));
 sky130_fd_sc_hd__o21ba_2 _20539_ (.A1(_07436_),
    .A2(_07438_),
    .B1_N(_07437_),
    .X(_07472_));
 sky130_fd_sc_hd__nand2b_2 _20540_ (.A_N(_07472_),
    .B(_07471_),
    .Y(_07473_));
 sky130_fd_sc_hd__xnor2_2 _20541_ (.A(_07471_),
    .B(_07472_),
    .Y(_07474_));
 sky130_fd_sc_hd__xnor2_2 _20542_ (.A(_07435_),
    .B(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__a21o_2 _20543_ (.A1(_07442_),
    .A2(_07444_),
    .B1(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__nand3_2 _20544_ (.A(_07442_),
    .B(_07444_),
    .C(_07475_),
    .Y(_07477_));
 sky130_fd_sc_hd__nand2_2 _20545_ (.A(_07476_),
    .B(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__xnor2_2 _20546_ (.A(_07465_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__o21a_2 _20547_ (.A1(_07432_),
    .A2(_07448_),
    .B1(_07446_),
    .X(_07480_));
 sky130_fd_sc_hd__and2b_2 _20548_ (.A_N(_07480_),
    .B(_07479_),
    .X(_07481_));
 sky130_fd_sc_hd__xnor2_2 _20549_ (.A(_07479_),
    .B(_07480_),
    .Y(_07482_));
 sky130_fd_sc_hd__and2_2 _20550_ (.A(_07430_),
    .B(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__nor2_2 _20551_ (.A(_07430_),
    .B(_07482_),
    .Y(_07484_));
 sky130_fd_sc_hd__or2_2 _20552_ (.A(_07483_),
    .B(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__a21oi_2 _20553_ (.A1(_07394_),
    .A2(_07453_),
    .B1(_07451_),
    .Y(_07486_));
 sky130_fd_sc_hd__nor2_2 _20554_ (.A(_07485_),
    .B(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__and2_2 _20555_ (.A(_07485_),
    .B(_07486_),
    .X(_07488_));
 sky130_fd_sc_hd__or2_2 _20556_ (.A(_07487_),
    .B(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__a31o_2 _20557_ (.A1(_07422_),
    .A2(_07427_),
    .A3(_07457_),
    .B1(_07456_),
    .X(_07490_));
 sky130_fd_sc_hd__a311oi_2 _20558_ (.A1(_07422_),
    .A2(_07427_),
    .A3(_07457_),
    .B1(_07489_),
    .C1(_07456_),
    .Y(_07491_));
 sky130_fd_sc_hd__and2_2 _20559_ (.A(_07489_),
    .B(_07490_),
    .X(_07492_));
 sky130_fd_sc_hd__nor2_2 _20560_ (.A(_07491_),
    .B(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__mux2_1 _20561_ (.A0(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[12] ),
    .A1(_07493_),
    .S(\systolic_inst.ce_local ),
    .X(_01614_));
 sky130_fd_sc_hd__nand2_2 _20562_ (.A(\systolic_inst.B_outs[5][6] ),
    .B(\systolic_inst.A_outs[5][7] ),
    .Y(_07494_));
 sky130_fd_sc_hd__nor2_2 _20563_ (.A(\systolic_inst.A_outs[5][6] ),
    .B(_11276_),
    .Y(_07495_));
 sky130_fd_sc_hd__xnor2_2 _20564_ (.A(_07494_),
    .B(_07495_),
    .Y(_07496_));
 sky130_fd_sc_hd__nand2b_2 _20565_ (.A_N(_07469_),
    .B(_07496_),
    .Y(_07497_));
 sky130_fd_sc_hd__xnor2_2 _20566_ (.A(_07469_),
    .B(_07496_),
    .Y(_07498_));
 sky130_fd_sc_hd__o21ai_2 _20567_ (.A1(_07467_),
    .A2(_07470_),
    .B1(_07498_),
    .Y(_07499_));
 sky130_fd_sc_hd__or3_2 _20568_ (.A(_07467_),
    .B(_07470_),
    .C(_07498_),
    .X(_07500_));
 sky130_fd_sc_hd__and2_2 _20569_ (.A(_07499_),
    .B(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__nand2_2 _20570_ (.A(_07435_),
    .B(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__or2_2 _20571_ (.A(_07435_),
    .B(_07501_),
    .X(_07503_));
 sky130_fd_sc_hd__nand2_2 _20572_ (.A(_07502_),
    .B(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__a21bo_2 _20573_ (.A1(_07435_),
    .A2(_07474_),
    .B1_N(_07473_),
    .X(_07505_));
 sky130_fd_sc_hd__nand2b_2 _20574_ (.A_N(_07504_),
    .B(_07505_),
    .Y(_07506_));
 sky130_fd_sc_hd__xor2_2 _20575_ (.A(_07504_),
    .B(_07505_),
    .X(_07507_));
 sky130_fd_sc_hd__xnor2_2 _20576_ (.A(_07465_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__o21a_2 _20577_ (.A1(_07464_),
    .A2(_07478_),
    .B1(_07476_),
    .X(_07509_));
 sky130_fd_sc_hd__and2b_2 _20578_ (.A_N(_07509_),
    .B(_07508_),
    .X(_07510_));
 sky130_fd_sc_hd__and2b_2 _20579_ (.A_N(_07508_),
    .B(_07509_),
    .X(_07511_));
 sky130_fd_sc_hd__nor2_2 _20580_ (.A(_07510_),
    .B(_07511_),
    .Y(_07512_));
 sky130_fd_sc_hd__xnor2_2 _20581_ (.A(_07463_),
    .B(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__o21ai_2 _20582_ (.A1(_07481_),
    .A2(_07483_),
    .B1(_07513_),
    .Y(_07514_));
 sky130_fd_sc_hd__or3_2 _20583_ (.A(_07481_),
    .B(_07483_),
    .C(_07513_),
    .X(_07515_));
 sky130_fd_sc_hd__and2_2 _20584_ (.A(_07514_),
    .B(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__or3_2 _20585_ (.A(_07487_),
    .B(_07491_),
    .C(_07516_),
    .X(_07517_));
 sky130_fd_sc_hd__nand2_2 _20586_ (.A(_07491_),
    .B(_07516_),
    .Y(_07518_));
 sky130_fd_sc_hd__nand2_2 _20587_ (.A(_07487_),
    .B(_07516_),
    .Y(_07519_));
 sky130_fd_sc_hd__and3_2 _20588_ (.A(\systolic_inst.ce_local ),
    .B(_07517_),
    .C(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__a22o_2 _20589_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[13] ),
    .B1(_07518_),
    .B2(_07520_),
    .X(_01615_));
 sky130_fd_sc_hd__and2_2 _20590_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[14] ),
    .X(_07521_));
 sky130_fd_sc_hd__o211ai_2 _20591_ (.A1(_11276_),
    .A2(\systolic_inst.A_outs[5][7] ),
    .B1(_07469_),
    .C1(_07494_),
    .Y(_07522_));
 sky130_fd_sc_hd__o311a_2 _20592_ (.A1(\systolic_inst.A_outs[5][6] ),
    .A2(_11276_),
    .A3(_07494_),
    .B1(_07497_),
    .C1(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__a31o_2 _20593_ (.A1(\systolic_inst.B_outs[5][5] ),
    .A2(\systolic_inst.B_outs[5][6] ),
    .A3(\systolic_inst.A_outs[5][7] ),
    .B1(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__nor2_2 _20594_ (.A(_07435_),
    .B(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__and2_2 _20595_ (.A(_07435_),
    .B(_07524_),
    .X(_07526_));
 sky130_fd_sc_hd__or2_2 _20596_ (.A(_07525_),
    .B(_07526_),
    .X(_07527_));
 sky130_fd_sc_hd__a21oi_2 _20597_ (.A1(_07499_),
    .A2(_07502_),
    .B1(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__and3_2 _20598_ (.A(_07499_),
    .B(_07502_),
    .C(_07527_),
    .X(_07529_));
 sky130_fd_sc_hd__nor2_2 _20599_ (.A(_07528_),
    .B(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__xnor2_2 _20600_ (.A(_07464_),
    .B(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__o21a_2 _20601_ (.A1(_07464_),
    .A2(_07507_),
    .B1(_07506_),
    .X(_07532_));
 sky130_fd_sc_hd__and2b_2 _20602_ (.A_N(_07532_),
    .B(_07531_),
    .X(_07533_));
 sky130_fd_sc_hd__and2b_2 _20603_ (.A_N(_07531_),
    .B(_07532_),
    .X(_07534_));
 sky130_fd_sc_hd__nor2_2 _20604_ (.A(_07533_),
    .B(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__xnor2_2 _20605_ (.A(_07463_),
    .B(_07535_),
    .Y(_07536_));
 sky130_fd_sc_hd__a31o_2 _20606_ (.A1(_07323_),
    .A2(_07461_),
    .A3(_07512_),
    .B1(_07510_),
    .X(_07537_));
 sky130_fd_sc_hd__xnor2_2 _20607_ (.A(_07536_),
    .B(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand4_2 _20608_ (.A(_07514_),
    .B(_07518_),
    .C(_07519_),
    .D(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__a31o_2 _20609_ (.A1(_07514_),
    .A2(_07518_),
    .A3(_07519_),
    .B1(_07538_),
    .X(_07540_));
 sky130_fd_sc_hd__a31o_2 _20610_ (.A1(\systolic_inst.ce_local ),
    .A2(_07539_),
    .A3(_07540_),
    .B1(_07521_),
    .X(_01616_));
 sky130_fd_sc_hd__and2_2 _20611_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .X(_07541_));
 sky130_fd_sc_hd__a31o_2 _20612_ (.A1(_07323_),
    .A2(_07461_),
    .A3(_07535_),
    .B1(_07533_),
    .X(_07542_));
 sky130_fd_sc_hd__a21oi_2 _20613_ (.A1(_07465_),
    .A2(_07530_),
    .B1(_07528_),
    .Y(_07543_));
 sky130_fd_sc_hd__xnor2_2 _20614_ (.A(_07462_),
    .B(_07525_),
    .Y(_07544_));
 sky130_fd_sc_hd__xnor2_2 _20615_ (.A(_07543_),
    .B(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__xnor2_2 _20616_ (.A(_07542_),
    .B(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__a21oi_2 _20617_ (.A1(_07536_),
    .A2(_07537_),
    .B1(_07546_),
    .Y(_07547_));
 sky130_fd_sc_hd__a31o_2 _20618_ (.A1(\systolic_inst.ce_local ),
    .A2(_07540_),
    .A3(_07547_),
    .B1(_07541_),
    .X(_01617_));
 sky130_fd_sc_hd__a21o_2 _20619_ (.A1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[5][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_07548_));
 sky130_fd_sc_hd__a21oi_2 _20620_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[5][0] ),
    .Y(_07549_));
 sky130_fd_sc_hd__a21oi_2 _20621_ (.A1(\systolic_inst.ce_local ),
    .A2(_07548_),
    .B1(_07549_),
    .Y(_01618_));
 sky130_fd_sc_hd__and2_2 _20622_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[5][1] ),
    .X(_07550_));
 sky130_fd_sc_hd__nand2_2 _20623_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[5][1] ),
    .Y(_07551_));
 sky130_fd_sc_hd__or2_2 _20624_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[5][1] ),
    .X(_07552_));
 sky130_fd_sc_hd__and4_2 _20625_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[5][0] ),
    .C(_07551_),
    .D(_07552_),
    .X(_07553_));
 sky130_fd_sc_hd__inv_2 _20626_ (.A(_07553_),
    .Y(_07554_));
 sky130_fd_sc_hd__a22o_2 _20627_ (.A1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[5][0] ),
    .B1(_07551_),
    .B2(_07552_),
    .X(_07555_));
 sky130_fd_sc_hd__a32o_2 _20628_ (.A1(_11712_),
    .A2(_07554_),
    .A3(_07555_),
    .B1(\systolic_inst.acc_wires[5][1] ),
    .B2(_11258_),
    .X(_01619_));
 sky130_fd_sc_hd__nand2_2 _20629_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[5][2] ),
    .Y(_07556_));
 sky130_fd_sc_hd__or2_2 _20630_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[5][2] ),
    .X(_07557_));
 sky130_fd_sc_hd__a31o_2 _20631_ (.A1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[5][0] ),
    .A3(_07552_),
    .B1(_07550_),
    .X(_07558_));
 sky130_fd_sc_hd__a21o_2 _20632_ (.A1(_07556_),
    .A2(_07557_),
    .B1(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__and3_2 _20633_ (.A(_07556_),
    .B(_07557_),
    .C(_07558_),
    .X(_07560_));
 sky130_fd_sc_hd__inv_2 _20634_ (.A(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__a32o_2 _20635_ (.A1(_11712_),
    .A2(_07559_),
    .A3(_07561_),
    .B1(\systolic_inst.acc_wires[5][2] ),
    .B2(_11258_),
    .X(_01620_));
 sky130_fd_sc_hd__nand2_2 _20636_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[5][3] ),
    .Y(_07562_));
 sky130_fd_sc_hd__or2_2 _20637_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[5][3] ),
    .X(_07563_));
 sky130_fd_sc_hd__a21bo_2 _20638_ (.A1(_07557_),
    .A2(_07558_),
    .B1_N(_07556_),
    .X(_07564_));
 sky130_fd_sc_hd__and3_2 _20639_ (.A(_07562_),
    .B(_07563_),
    .C(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__inv_2 _20640_ (.A(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__a21o_2 _20641_ (.A1(_07562_),
    .A2(_07563_),
    .B1(_07564_),
    .X(_07567_));
 sky130_fd_sc_hd__a32o_2 _20642_ (.A1(_11712_),
    .A2(_07566_),
    .A3(_07567_),
    .B1(\systolic_inst.acc_wires[5][3] ),
    .B2(_11258_),
    .X(_01621_));
 sky130_fd_sc_hd__nand2_2 _20643_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[5][4] ),
    .Y(_07568_));
 sky130_fd_sc_hd__or2_2 _20644_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[5][4] ),
    .X(_07569_));
 sky130_fd_sc_hd__a21bo_2 _20645_ (.A1(_07563_),
    .A2(_07564_),
    .B1_N(_07562_),
    .X(_07570_));
 sky130_fd_sc_hd__a21o_2 _20646_ (.A1(_07568_),
    .A2(_07569_),
    .B1(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__and3_2 _20647_ (.A(_07568_),
    .B(_07569_),
    .C(_07570_),
    .X(_07572_));
 sky130_fd_sc_hd__inv_2 _20648_ (.A(_07572_),
    .Y(_07573_));
 sky130_fd_sc_hd__a32o_2 _20649_ (.A1(_11712_),
    .A2(_07571_),
    .A3(_07573_),
    .B1(\systolic_inst.acc_wires[5][4] ),
    .B2(_11258_),
    .X(_01622_));
 sky130_fd_sc_hd__nand2_2 _20650_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[5][5] ),
    .Y(_07574_));
 sky130_fd_sc_hd__or2_2 _20651_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[5][5] ),
    .X(_07575_));
 sky130_fd_sc_hd__a21bo_2 _20652_ (.A1(_07569_),
    .A2(_07570_),
    .B1_N(_07568_),
    .X(_07576_));
 sky130_fd_sc_hd__a21o_2 _20653_ (.A1(_07574_),
    .A2(_07575_),
    .B1(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__and3_2 _20654_ (.A(_07574_),
    .B(_07575_),
    .C(_07576_),
    .X(_07578_));
 sky130_fd_sc_hd__inv_2 _20655_ (.A(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__a32o_2 _20656_ (.A1(_11712_),
    .A2(_07577_),
    .A3(_07579_),
    .B1(\systolic_inst.acc_wires[5][5] ),
    .B2(_11258_),
    .X(_01623_));
 sky130_fd_sc_hd__nand2_2 _20657_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[5][6] ),
    .Y(_07580_));
 sky130_fd_sc_hd__or2_2 _20658_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[5][6] ),
    .X(_07581_));
 sky130_fd_sc_hd__a21bo_2 _20659_ (.A1(_07575_),
    .A2(_07576_),
    .B1_N(_07574_),
    .X(_07582_));
 sky130_fd_sc_hd__a21o_2 _20660_ (.A1(_07580_),
    .A2(_07581_),
    .B1(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__and3_2 _20661_ (.A(_07580_),
    .B(_07581_),
    .C(_07582_),
    .X(_07584_));
 sky130_fd_sc_hd__inv_2 _20662_ (.A(_07584_),
    .Y(_07585_));
 sky130_fd_sc_hd__a32o_2 _20663_ (.A1(_11712_),
    .A2(_07583_),
    .A3(_07585_),
    .B1(\systolic_inst.acc_wires[5][6] ),
    .B2(_11258_),
    .X(_01624_));
 sky130_fd_sc_hd__nand2_2 _20664_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[5][7] ),
    .Y(_07586_));
 sky130_fd_sc_hd__or2_2 _20665_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[5][7] ),
    .X(_07587_));
 sky130_fd_sc_hd__a21bo_2 _20666_ (.A1(_07581_),
    .A2(_07582_),
    .B1_N(_07580_),
    .X(_07588_));
 sky130_fd_sc_hd__nand3_2 _20667_ (.A(_07586_),
    .B(_07587_),
    .C(_07588_),
    .Y(_07589_));
 sky130_fd_sc_hd__a21o_2 _20668_ (.A1(_07586_),
    .A2(_07587_),
    .B1(_07588_),
    .X(_07590_));
 sky130_fd_sc_hd__a32o_2 _20669_ (.A1(_11712_),
    .A2(_07589_),
    .A3(_07590_),
    .B1(\systolic_inst.acc_wires[5][7] ),
    .B2(_11258_),
    .X(_01625_));
 sky130_fd_sc_hd__a21bo_2 _20670_ (.A1(_07587_),
    .A2(_07588_),
    .B1_N(_07586_),
    .X(_07591_));
 sky130_fd_sc_hd__xor2_2 _20671_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[5][8] ),
    .X(_07592_));
 sky130_fd_sc_hd__and2_2 _20672_ (.A(_07591_),
    .B(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__o21ai_2 _20673_ (.A1(_07591_),
    .A2(_07592_),
    .B1(_11712_),
    .Y(_07594_));
 sky130_fd_sc_hd__a2bb2o_2 _20674_ (.A1_N(_07594_),
    .A2_N(_07593_),
    .B1(\systolic_inst.acc_wires[5][8] ),
    .B2(_11258_),
    .X(_01626_));
 sky130_fd_sc_hd__xor2_2 _20675_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[5][9] ),
    .X(_07595_));
 sky130_fd_sc_hd__a211o_2 _20676_ (.A1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[5][8] ),
    .B1(_07593_),
    .C1(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__nand2_2 _20677_ (.A(_07592_),
    .B(_07595_),
    .Y(_07597_));
 sky130_fd_sc_hd__nand2_2 _20678_ (.A(_07593_),
    .B(_07595_),
    .Y(_07598_));
 sky130_fd_sc_hd__and3_2 _20679_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[5][8] ),
    .C(_07595_),
    .X(_07599_));
 sky130_fd_sc_hd__nor2_2 _20680_ (.A(_11713_),
    .B(_07599_),
    .Y(_07600_));
 sky130_fd_sc_hd__a32o_2 _20681_ (.A1(_07596_),
    .A2(_07598_),
    .A3(_07600_),
    .B1(\systolic_inst.acc_wires[5][9] ),
    .B2(_11258_),
    .X(_01627_));
 sky130_fd_sc_hd__nand2_2 _20682_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[5][10] ),
    .Y(_07601_));
 sky130_fd_sc_hd__or2_2 _20683_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[5][10] ),
    .X(_07602_));
 sky130_fd_sc_hd__and2_2 _20684_ (.A(_07601_),
    .B(_07602_),
    .X(_07603_));
 sky130_fd_sc_hd__a21oi_2 _20685_ (.A1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[5][9] ),
    .B1(_07599_),
    .Y(_07604_));
 sky130_fd_sc_hd__nand2_2 _20686_ (.A(_07598_),
    .B(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__xor2_2 _20687_ (.A(_07603_),
    .B(_07605_),
    .X(_07606_));
 sky130_fd_sc_hd__a22o_2 _20688_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][10] ),
    .B1(_11712_),
    .B2(_07606_),
    .X(_01628_));
 sky130_fd_sc_hd__nor2_2 _20689_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[5][11] ),
    .Y(_07607_));
 sky130_fd_sc_hd__or2_2 _20690_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[5][11] ),
    .X(_07608_));
 sky130_fd_sc_hd__nand2_2 _20691_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[5][11] ),
    .Y(_07609_));
 sky130_fd_sc_hd__nand2_2 _20692_ (.A(_07608_),
    .B(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__a21bo_2 _20693_ (.A1(_07603_),
    .A2(_07605_),
    .B1_N(_07601_),
    .X(_07611_));
 sky130_fd_sc_hd__xnor2_2 _20694_ (.A(_07610_),
    .B(_07611_),
    .Y(_07612_));
 sky130_fd_sc_hd__a22o_2 _20695_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][11] ),
    .B1(_11712_),
    .B2(_07612_),
    .X(_01629_));
 sky130_fd_sc_hd__nand3_2 _20696_ (.A(_07603_),
    .B(_07608_),
    .C(_07609_),
    .Y(_07613_));
 sky130_fd_sc_hd__nor2_2 _20697_ (.A(_07597_),
    .B(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__o2bb2a_2 _20698_ (.A1_N(_07591_),
    .A2_N(_07614_),
    .B1(_07604_),
    .B2(_07613_),
    .X(_07615_));
 sky130_fd_sc_hd__o21a_2 _20699_ (.A1(_07601_),
    .A2(_07607_),
    .B1(_07609_),
    .X(_07616_));
 sky130_fd_sc_hd__xnor2_2 _20700_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[5][12] ),
    .Y(_07617_));
 sky130_fd_sc_hd__and3_2 _20701_ (.A(_07615_),
    .B(_07616_),
    .C(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__a21oi_2 _20702_ (.A1(_07615_),
    .A2(_07616_),
    .B1(_07617_),
    .Y(_07619_));
 sky130_fd_sc_hd__nor2_2 _20703_ (.A(_07618_),
    .B(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__a22o_2 _20704_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][12] ),
    .B1(_11712_),
    .B2(_07620_),
    .X(_01630_));
 sky130_fd_sc_hd__xor2_2 _20705_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[5][13] ),
    .X(_07621_));
 sky130_fd_sc_hd__a211o_2 _20706_ (.A1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[5][12] ),
    .B1(_07619_),
    .C1(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__nand2b_2 _20707_ (.A_N(_07617_),
    .B(_07621_),
    .Y(_07623_));
 sky130_fd_sc_hd__a21o_2 _20708_ (.A1(_07615_),
    .A2(_07616_),
    .B1(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__and3_2 _20709_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[5][12] ),
    .C(_07621_),
    .X(_07625_));
 sky130_fd_sc_hd__nor2_2 _20710_ (.A(_11713_),
    .B(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__a32o_2 _20711_ (.A1(_07622_),
    .A2(_07624_),
    .A3(_07626_),
    .B1(\systolic_inst.acc_wires[5][13] ),
    .B2(_11258_),
    .X(_01631_));
 sky130_fd_sc_hd__or2_2 _20712_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[5][14] ),
    .X(_07627_));
 sky130_fd_sc_hd__nand2_2 _20713_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[5][14] ),
    .Y(_07628_));
 sky130_fd_sc_hd__and2_2 _20714_ (.A(_07627_),
    .B(_07628_),
    .X(_07629_));
 sky130_fd_sc_hd__a21oi_2 _20715_ (.A1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[5][13] ),
    .B1(_07625_),
    .Y(_07630_));
 sky130_fd_sc_hd__nand2_2 _20716_ (.A(_07624_),
    .B(_07630_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_2 _20717_ (.A(_07629_),
    .B(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__or2_2 _20718_ (.A(_07629_),
    .B(_07631_),
    .X(_07633_));
 sky130_fd_sc_hd__a32o_2 _20719_ (.A1(_11712_),
    .A2(_07632_),
    .A3(_07633_),
    .B1(\systolic_inst.acc_wires[5][14] ),
    .B2(_11258_),
    .X(_01632_));
 sky130_fd_sc_hd__nor2_2 _20720_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][15] ),
    .Y(_07634_));
 sky130_fd_sc_hd__and2_2 _20721_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][15] ),
    .X(_07635_));
 sky130_fd_sc_hd__a211o_2 _20722_ (.A1(_07628_),
    .A2(_07632_),
    .B1(_07634_),
    .C1(_07635_),
    .X(_07636_));
 sky130_fd_sc_hd__o211ai_2 _20723_ (.A1(_07634_),
    .A2(_07635_),
    .B1(_07628_),
    .C1(_07632_),
    .Y(_07637_));
 sky130_fd_sc_hd__a32o_2 _20724_ (.A1(_11712_),
    .A2(_07636_),
    .A3(_07637_),
    .B1(\systolic_inst.acc_wires[5][15] ),
    .B2(_11258_),
    .X(_01633_));
 sky130_fd_sc_hd__or3b_2 _20725_ (.A(_07634_),
    .B(_07635_),
    .C_N(_07629_),
    .X(_07638_));
 sky130_fd_sc_hd__a21o_2 _20726_ (.A1(_07624_),
    .A2(_07630_),
    .B1(_07638_),
    .X(_07639_));
 sky130_fd_sc_hd__o21ba_2 _20727_ (.A1(_07628_),
    .A2(_07634_),
    .B1_N(_07635_),
    .X(_07640_));
 sky130_fd_sc_hd__and2_2 _20728_ (.A(_07639_),
    .B(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__xnor2_2 _20729_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][16] ),
    .Y(_07642_));
 sky130_fd_sc_hd__nand2_2 _20730_ (.A(_07641_),
    .B(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__nor2_2 _20731_ (.A(_07641_),
    .B(_07642_),
    .Y(_07644_));
 sky130_fd_sc_hd__nor2_2 _20732_ (.A(_11713_),
    .B(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__a22o_2 _20733_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][16] ),
    .B1(_07643_),
    .B2(_07645_),
    .X(_01634_));
 sky130_fd_sc_hd__xor2_2 _20734_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][17] ),
    .X(_07646_));
 sky130_fd_sc_hd__inv_2 _20735_ (.A(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__a21oi_2 _20736_ (.A1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[5][16] ),
    .B1(_07644_),
    .Y(_07648_));
 sky130_fd_sc_hd__xnor2_2 _20737_ (.A(_07646_),
    .B(_07648_),
    .Y(_07649_));
 sky130_fd_sc_hd__a22o_2 _20738_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][17] ),
    .B1(_11712_),
    .B2(_07649_),
    .X(_01635_));
 sky130_fd_sc_hd__or2_2 _20739_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][18] ),
    .X(_07650_));
 sky130_fd_sc_hd__nand2_2 _20740_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][18] ),
    .Y(_07651_));
 sky130_fd_sc_hd__nand2_2 _20741_ (.A(_07650_),
    .B(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__o21a_2 _20742_ (.A1(\systolic_inst.acc_wires[5][16] ),
    .A2(\systolic_inst.acc_wires[5][17] ),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .X(_07653_));
 sky130_fd_sc_hd__a21oi_2 _20743_ (.A1(_07644_),
    .A2(_07646_),
    .B1(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__xor2_2 _20744_ (.A(_07652_),
    .B(_07654_),
    .X(_07655_));
 sky130_fd_sc_hd__a22o_2 _20745_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][18] ),
    .B1(_11712_),
    .B2(_07655_),
    .X(_01636_));
 sky130_fd_sc_hd__xnor2_2 _20746_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][19] ),
    .Y(_07656_));
 sky130_fd_sc_hd__o21ai_2 _20747_ (.A1(_07652_),
    .A2(_07654_),
    .B1(_07651_),
    .Y(_07657_));
 sky130_fd_sc_hd__xnor2_2 _20748_ (.A(_07656_),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__a22o_2 _20749_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][19] ),
    .B1(_11712_),
    .B2(_07658_),
    .X(_01637_));
 sky130_fd_sc_hd__or2_2 _20750_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][20] ),
    .X(_07659_));
 sky130_fd_sc_hd__nand2_2 _20751_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][20] ),
    .Y(_07660_));
 sky130_fd_sc_hd__and2_2 _20752_ (.A(_07659_),
    .B(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__or4_2 _20753_ (.A(_07642_),
    .B(_07647_),
    .C(_07652_),
    .D(_07656_),
    .X(_07662_));
 sky130_fd_sc_hd__nor2_2 _20754_ (.A(_07641_),
    .B(_07662_),
    .Y(_07663_));
 sky130_fd_sc_hd__o41a_2 _20755_ (.A1(\systolic_inst.acc_wires[5][16] ),
    .A2(\systolic_inst.acc_wires[5][17] ),
    .A3(\systolic_inst.acc_wires[5][18] ),
    .A4(\systolic_inst.acc_wires[5][19] ),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .X(_07664_));
 sky130_fd_sc_hd__or3_2 _20756_ (.A(_07661_),
    .B(_07663_),
    .C(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__o21ai_2 _20757_ (.A1(_07663_),
    .A2(_07664_),
    .B1(_07661_),
    .Y(_07666_));
 sky130_fd_sc_hd__a32o_2 _20758_ (.A1(_11712_),
    .A2(_07665_),
    .A3(_07666_),
    .B1(\systolic_inst.acc_wires[5][20] ),
    .B2(_11258_),
    .X(_01638_));
 sky130_fd_sc_hd__xnor2_2 _20759_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][21] ),
    .Y(_07667_));
 sky130_fd_sc_hd__inv_2 _20760_ (.A(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__a21oi_2 _20761_ (.A1(_07660_),
    .A2(_07666_),
    .B1(_07667_),
    .Y(_07669_));
 sky130_fd_sc_hd__a31o_2 _20762_ (.A1(_07660_),
    .A2(_07666_),
    .A3(_07667_),
    .B1(_11713_),
    .X(_07670_));
 sky130_fd_sc_hd__a2bb2o_2 _20763_ (.A1_N(_07670_),
    .A2_N(_07669_),
    .B1(\systolic_inst.acc_wires[5][21] ),
    .B2(_11258_),
    .X(_01639_));
 sky130_fd_sc_hd__or2_2 _20764_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][22] ),
    .X(_07671_));
 sky130_fd_sc_hd__nand2_2 _20765_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][22] ),
    .Y(_07672_));
 sky130_fd_sc_hd__and2_2 _20766_ (.A(_07671_),
    .B(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__o21a_2 _20767_ (.A1(\systolic_inst.acc_wires[5][20] ),
    .A2(\systolic_inst.acc_wires[5][21] ),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .X(_07674_));
 sky130_fd_sc_hd__nor2_2 _20768_ (.A(_07666_),
    .B(_07667_),
    .Y(_07675_));
 sky130_fd_sc_hd__o21ai_2 _20769_ (.A1(_07674_),
    .A2(_07675_),
    .B1(_07673_),
    .Y(_07676_));
 sky130_fd_sc_hd__or3_2 _20770_ (.A(_07673_),
    .B(_07674_),
    .C(_07675_),
    .X(_07677_));
 sky130_fd_sc_hd__a32o_2 _20771_ (.A1(_11712_),
    .A2(_07676_),
    .A3(_07677_),
    .B1(\systolic_inst.acc_wires[5][22] ),
    .B2(_11258_),
    .X(_01640_));
 sky130_fd_sc_hd__xor2_2 _20772_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][23] ),
    .X(_07678_));
 sky130_fd_sc_hd__inv_2 _20773_ (.A(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__nand3_2 _20774_ (.A(_07672_),
    .B(_07676_),
    .C(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__a21o_2 _20775_ (.A1(_07672_),
    .A2(_07676_),
    .B1(_07679_),
    .X(_07681_));
 sky130_fd_sc_hd__a32o_2 _20776_ (.A1(_11712_),
    .A2(_07680_),
    .A3(_07681_),
    .B1(\systolic_inst.acc_wires[5][23] ),
    .B2(_11258_),
    .X(_01641_));
 sky130_fd_sc_hd__nand4_2 _20777_ (.A(_07661_),
    .B(_07668_),
    .C(_07673_),
    .D(_07678_),
    .Y(_07682_));
 sky130_fd_sc_hd__a211o_2 _20778_ (.A1(_07639_),
    .A2(_07640_),
    .B1(_07662_),
    .C1(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__o41a_2 _20779_ (.A1(\systolic_inst.acc_wires[5][20] ),
    .A2(\systolic_inst.acc_wires[5][21] ),
    .A3(\systolic_inst.acc_wires[5][22] ),
    .A4(\systolic_inst.acc_wires[5][23] ),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .X(_07684_));
 sky130_fd_sc_hd__nor2_2 _20780_ (.A(_07664_),
    .B(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__nor2_2 _20781_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][24] ),
    .Y(_07686_));
 sky130_fd_sc_hd__and2_2 _20782_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][24] ),
    .X(_07687_));
 sky130_fd_sc_hd__or2_2 _20783_ (.A(_07686_),
    .B(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__a21oi_2 _20784_ (.A1(_07683_),
    .A2(_07685_),
    .B1(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__a31o_2 _20785_ (.A1(_07683_),
    .A2(_07685_),
    .A3(_07688_),
    .B1(_11713_),
    .X(_07690_));
 sky130_fd_sc_hd__a2bb2o_2 _20786_ (.A1_N(_07690_),
    .A2_N(_07689_),
    .B1(\systolic_inst.acc_wires[5][24] ),
    .B2(_11258_),
    .X(_01642_));
 sky130_fd_sc_hd__xor2_2 _20787_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][25] ),
    .X(_07691_));
 sky130_fd_sc_hd__or3_2 _20788_ (.A(_07687_),
    .B(_07689_),
    .C(_07691_),
    .X(_07692_));
 sky130_fd_sc_hd__o21ai_2 _20789_ (.A1(_07687_),
    .A2(_07689_),
    .B1(_07691_),
    .Y(_07693_));
 sky130_fd_sc_hd__a32o_2 _20790_ (.A1(_11712_),
    .A2(_07692_),
    .A3(_07693_),
    .B1(\systolic_inst.acc_wires[5][25] ),
    .B2(_11258_),
    .X(_01643_));
 sky130_fd_sc_hd__or2_2 _20791_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][26] ),
    .X(_07694_));
 sky130_fd_sc_hd__nand2_2 _20792_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][26] ),
    .Y(_07695_));
 sky130_fd_sc_hd__nand2_2 _20793_ (.A(_07694_),
    .B(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__o21a_2 _20794_ (.A1(\systolic_inst.acc_wires[5][24] ),
    .A2(\systolic_inst.acc_wires[5][25] ),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .X(_07697_));
 sky130_fd_sc_hd__a21o_2 _20795_ (.A1(_07689_),
    .A2(_07691_),
    .B1(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__xnor2_2 _20796_ (.A(_07696_),
    .B(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__a22o_2 _20797_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][26] ),
    .B1(_11712_),
    .B2(_07699_),
    .X(_01644_));
 sky130_fd_sc_hd__xnor2_2 _20798_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][27] ),
    .Y(_07700_));
 sky130_fd_sc_hd__a21bo_2 _20799_ (.A1(_07694_),
    .A2(_07698_),
    .B1_N(_07695_),
    .X(_07701_));
 sky130_fd_sc_hd__xnor2_2 _20800_ (.A(_07700_),
    .B(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__a22o_2 _20801_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][27] ),
    .B1(_11712_),
    .B2(_07702_),
    .X(_01645_));
 sky130_fd_sc_hd__nor2_2 _20802_ (.A(_07696_),
    .B(_07700_),
    .Y(_07703_));
 sky130_fd_sc_hd__o21a_2 _20803_ (.A1(\systolic_inst.acc_wires[5][26] ),
    .A2(\systolic_inst.acc_wires[5][27] ),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .X(_07704_));
 sky130_fd_sc_hd__a311oi_2 _20804_ (.A1(_07689_),
    .A2(_07691_),
    .A3(_07703_),
    .B1(_07704_),
    .C1(_07697_),
    .Y(_07705_));
 sky130_fd_sc_hd__or2_2 _20805_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][28] ),
    .X(_07706_));
 sky130_fd_sc_hd__nand2_2 _20806_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][28] ),
    .Y(_07707_));
 sky130_fd_sc_hd__nand2_2 _20807_ (.A(_07706_),
    .B(_07707_),
    .Y(_07708_));
 sky130_fd_sc_hd__xor2_2 _20808_ (.A(_07705_),
    .B(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__a22o_2 _20809_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][28] ),
    .B1(_11712_),
    .B2(_07709_),
    .X(_01646_));
 sky130_fd_sc_hd__xor2_2 _20810_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][29] ),
    .X(_07710_));
 sky130_fd_sc_hd__inv_2 _20811_ (.A(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__o21a_2 _20812_ (.A1(_07705_),
    .A2(_07708_),
    .B1(_07707_),
    .X(_07712_));
 sky130_fd_sc_hd__xnor2_2 _20813_ (.A(_07710_),
    .B(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__a22o_2 _20814_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[5][29] ),
    .B1(_11712_),
    .B2(_07713_),
    .X(_01647_));
 sky130_fd_sc_hd__o21ai_2 _20815_ (.A1(\systolic_inst.acc_wires[5][28] ),
    .A2(\systolic_inst.acc_wires[5][29] ),
    .B1(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .Y(_07714_));
 sky130_fd_sc_hd__o31a_2 _20816_ (.A1(_07705_),
    .A2(_07708_),
    .A3(_07711_),
    .B1(_07714_),
    .X(_07715_));
 sky130_fd_sc_hd__nand2_2 _20817_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][30] ),
    .Y(_07716_));
 sky130_fd_sc_hd__or2_2 _20818_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][30] ),
    .X(_07717_));
 sky130_fd_sc_hd__nand2_2 _20819_ (.A(_07716_),
    .B(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__nand2_2 _20820_ (.A(_07715_),
    .B(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__or2_2 _20821_ (.A(_07715_),
    .B(_07718_),
    .X(_07720_));
 sky130_fd_sc_hd__a32o_2 _20822_ (.A1(_11712_),
    .A2(_07719_),
    .A3(_07720_),
    .B1(\systolic_inst.acc_wires[5][30] ),
    .B2(_11258_),
    .X(_01648_));
 sky130_fd_sc_hd__xnor2_2 _20823_ (.A(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[5][31] ),
    .Y(_07721_));
 sky130_fd_sc_hd__a21oi_2 _20824_ (.A1(_07716_),
    .A2(_07720_),
    .B1(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__a31o_2 _20825_ (.A1(_07716_),
    .A2(_07720_),
    .A3(_07721_),
    .B1(_11713_),
    .X(_07723_));
 sky130_fd_sc_hd__a2bb2o_2 _20826_ (.A1_N(_07723_),
    .A2_N(_07722_),
    .B1(\systolic_inst.acc_wires[5][31] ),
    .B2(_11258_),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _20827_ (.A0(\systolic_inst.A_outs[4][0] ),
    .A1(\systolic_inst.A_shift[8][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _20828_ (.A0(\systolic_inst.A_outs[4][1] ),
    .A1(\systolic_inst.A_shift[8][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _20829_ (.A0(\systolic_inst.A_outs[4][2] ),
    .A1(\systolic_inst.A_shift[8][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _20830_ (.A0(\systolic_inst.A_outs[4][3] ),
    .A1(\systolic_inst.A_shift[8][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _20831_ (.A0(\systolic_inst.A_outs[4][4] ),
    .A1(\systolic_inst.A_shift[8][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _20832_ (.A0(\systolic_inst.A_outs[4][5] ),
    .A1(\systolic_inst.A_shift[8][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _20833_ (.A0(\systolic_inst.A_outs[4][6] ),
    .A1(\systolic_inst.A_shift[8][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _20834_ (.A0(\systolic_inst.A_outs[4][7] ),
    .A1(\systolic_inst.A_shift[8][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _20835_ (.A0(\systolic_inst.B_outs[3][0] ),
    .A1(\systolic_inst.B_shift[3][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _20836_ (.A0(\systolic_inst.B_outs[3][1] ),
    .A1(\systolic_inst.B_shift[3][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _20837_ (.A0(\systolic_inst.B_outs[3][2] ),
    .A1(\systolic_inst.B_shift[3][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _20838_ (.A0(\systolic_inst.B_outs[3][3] ),
    .A1(\systolic_inst.B_shift[3][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _20839_ (.A0(\systolic_inst.B_outs[3][4] ),
    .A1(\systolic_inst.B_shift[3][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _20840_ (.A0(\systolic_inst.B_outs[3][5] ),
    .A1(\systolic_inst.B_shift[3][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _20841_ (.A0(\systolic_inst.B_outs[3][6] ),
    .A1(\systolic_inst.B_shift[3][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _20842_ (.A0(\systolic_inst.B_outs[3][7] ),
    .A1(\systolic_inst.B_shift[3][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01665_));
 sky130_fd_sc_hd__and3_2 _20843_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[4][0] ),
    .C(\systolic_inst.A_outs[4][0] ),
    .X(_07724_));
 sky130_fd_sc_hd__a21o_2 _20844_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[0] ),
    .B1(_07724_),
    .X(_01666_));
 sky130_fd_sc_hd__and4_2 _20845_ (.A(\systolic_inst.B_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][0] ),
    .C(\systolic_inst.A_outs[4][1] ),
    .D(\systolic_inst.B_outs[4][1] ),
    .X(_07725_));
 sky130_fd_sc_hd__a22o_2 _20846_ (.A1(\systolic_inst.B_outs[4][0] ),
    .A2(\systolic_inst.A_outs[4][1] ),
    .B1(\systolic_inst.B_outs[4][1] ),
    .B2(\systolic_inst.A_outs[4][0] ),
    .X(_07726_));
 sky130_fd_sc_hd__nand2_2 _20847_ (.A(\systolic_inst.ce_local ),
    .B(_07726_),
    .Y(_07727_));
 sky130_fd_sc_hd__a2bb2o_2 _20848_ (.A1_N(_07727_),
    .A2_N(_07725_),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01667_));
 sky130_fd_sc_hd__a22o_2 _20849_ (.A1(\systolic_inst.A_outs[4][1] ),
    .A2(\systolic_inst.B_outs[4][1] ),
    .B1(\systolic_inst.B_outs[4][2] ),
    .B2(\systolic_inst.A_outs[4][0] ),
    .X(_07728_));
 sky130_fd_sc_hd__and4_2 _20850_ (.A(\systolic_inst.A_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][1] ),
    .C(\systolic_inst.B_outs[4][1] ),
    .D(\systolic_inst.B_outs[4][2] ),
    .X(_07729_));
 sky130_fd_sc_hd__inv_2 _20851_ (.A(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__and4_2 _20852_ (.A(\systolic_inst.B_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][2] ),
    .C(_07728_),
    .D(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__a22oi_2 _20853_ (.A1(\systolic_inst.B_outs[4][0] ),
    .A2(\systolic_inst.A_outs[4][2] ),
    .B1(_07728_),
    .B2(_07730_),
    .Y(_07732_));
 sky130_fd_sc_hd__nor2_2 _20854_ (.A(_07731_),
    .B(_07732_),
    .Y(_07733_));
 sky130_fd_sc_hd__or2_2 _20855_ (.A(_07725_),
    .B(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__and2_2 _20856_ (.A(_07725_),
    .B(_07733_),
    .X(_07735_));
 sky130_fd_sc_hd__nor2_2 _20857_ (.A(_11258_),
    .B(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__a22o_2 _20858_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[2] ),
    .B1(_07734_),
    .B2(_07736_),
    .X(_01668_));
 sky130_fd_sc_hd__a21o_2 _20859_ (.A1(\systolic_inst.A_outs[4][0] ),
    .A2(\systolic_inst.B_outs[4][3] ),
    .B1(_07729_),
    .X(_07737_));
 sky130_fd_sc_hd__nand2_2 _20860_ (.A(\systolic_inst.B_outs[4][3] ),
    .B(_07729_),
    .Y(_07738_));
 sky130_fd_sc_hd__and2_2 _20861_ (.A(_07737_),
    .B(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__a22o_2 _20862_ (.A1(\systolic_inst.B_outs[4][1] ),
    .A2(\systolic_inst.A_outs[4][2] ),
    .B1(\systolic_inst.B_outs[4][2] ),
    .B2(\systolic_inst.A_outs[4][1] ),
    .X(_07740_));
 sky130_fd_sc_hd__nand4_2 _20863_ (.A(\systolic_inst.A_outs[4][1] ),
    .B(\systolic_inst.B_outs[4][1] ),
    .C(\systolic_inst.A_outs[4][2] ),
    .D(\systolic_inst.B_outs[4][2] ),
    .Y(_07741_));
 sky130_fd_sc_hd__nand4_2 _20864_ (.A(\systolic_inst.B_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][3] ),
    .C(_07740_),
    .D(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__a22o_2 _20865_ (.A1(\systolic_inst.B_outs[4][0] ),
    .A2(\systolic_inst.A_outs[4][3] ),
    .B1(_07740_),
    .B2(_07741_),
    .X(_07743_));
 sky130_fd_sc_hd__and3_2 _20866_ (.A(_07731_),
    .B(_07742_),
    .C(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__a21o_2 _20867_ (.A1(_07742_),
    .A2(_07743_),
    .B1(_07731_),
    .X(_07745_));
 sky130_fd_sc_hd__nand2b_2 _20868_ (.A_N(_07744_),
    .B(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__xnor2_2 _20869_ (.A(_07739_),
    .B(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__and2_2 _20870_ (.A(_07735_),
    .B(_07747_),
    .X(_07748_));
 sky130_fd_sc_hd__o21ai_2 _20871_ (.A1(_07735_),
    .A2(_07747_),
    .B1(\systolic_inst.ce_local ),
    .Y(_07749_));
 sky130_fd_sc_hd__a2bb2o_2 _20872_ (.A1_N(_07749_),
    .A2_N(_07748_),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[3] ),
    .B2(_11258_),
    .X(_01669_));
 sky130_fd_sc_hd__and4_2 _20873_ (.A(\systolic_inst.A_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][1] ),
    .C(\systolic_inst.B_outs[4][3] ),
    .D(\systolic_inst.B_outs[4][4] ),
    .X(_07750_));
 sky130_fd_sc_hd__inv_2 _20874_ (.A(_07750_),
    .Y(_07751_));
 sky130_fd_sc_hd__a22oi_2 _20875_ (.A1(\systolic_inst.A_outs[4][1] ),
    .A2(\systolic_inst.B_outs[4][3] ),
    .B1(\systolic_inst.B_outs[4][4] ),
    .B2(\systolic_inst.A_outs[4][0] ),
    .Y(_07752_));
 sky130_fd_sc_hd__or2_2 _20876_ (.A(_07750_),
    .B(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__nor2_2 _20877_ (.A(_07741_),
    .B(_07753_),
    .Y(_07754_));
 sky130_fd_sc_hd__and2_2 _20878_ (.A(_07741_),
    .B(_07753_),
    .X(_07755_));
 sky130_fd_sc_hd__nor2_2 _20879_ (.A(_07754_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__a22o_2 _20880_ (.A1(\systolic_inst.A_outs[4][2] ),
    .A2(\systolic_inst.B_outs[4][2] ),
    .B1(\systolic_inst.A_outs[4][3] ),
    .B2(\systolic_inst.B_outs[4][1] ),
    .X(_07757_));
 sky130_fd_sc_hd__nand2_2 _20881_ (.A(\systolic_inst.B_outs[4][2] ),
    .B(\systolic_inst.A_outs[4][3] ),
    .Y(_07758_));
 sky130_fd_sc_hd__nand4_2 _20882_ (.A(\systolic_inst.B_outs[4][1] ),
    .B(\systolic_inst.A_outs[4][2] ),
    .C(\systolic_inst.B_outs[4][2] ),
    .D(\systolic_inst.A_outs[4][3] ),
    .Y(_07759_));
 sky130_fd_sc_hd__and4_2 _20883_ (.A(\systolic_inst.B_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][4] ),
    .C(_07757_),
    .D(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__a22oi_2 _20884_ (.A1(\systolic_inst.B_outs[4][0] ),
    .A2(\systolic_inst.A_outs[4][4] ),
    .B1(_07757_),
    .B2(_07759_),
    .Y(_07761_));
 sky130_fd_sc_hd__or3_2 _20885_ (.A(_07742_),
    .B(_07760_),
    .C(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__o21ai_2 _20886_ (.A1(_07760_),
    .A2(_07761_),
    .B1(_07742_),
    .Y(_07763_));
 sky130_fd_sc_hd__nand2_2 _20887_ (.A(_07762_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__xnor2_2 _20888_ (.A(_07756_),
    .B(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__a21oi_2 _20889_ (.A1(_07739_),
    .A2(_07745_),
    .B1(_07744_),
    .Y(_07766_));
 sky130_fd_sc_hd__and2b_2 _20890_ (.A_N(_07766_),
    .B(_07765_),
    .X(_07767_));
 sky130_fd_sc_hd__and2b_2 _20891_ (.A_N(_07765_),
    .B(_07766_),
    .X(_07768_));
 sky130_fd_sc_hd__nor2_2 _20892_ (.A(_07767_),
    .B(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__xnor2_2 _20893_ (.A(_07738_),
    .B(_07769_),
    .Y(_07770_));
 sky130_fd_sc_hd__or2_2 _20894_ (.A(_07748_),
    .B(_07770_),
    .X(_07771_));
 sky130_fd_sc_hd__and2_2 _20895_ (.A(_07748_),
    .B(_07770_),
    .X(_07772_));
 sky130_fd_sc_hd__nor2_2 _20896_ (.A(_11258_),
    .B(_07772_),
    .Y(_07773_));
 sky130_fd_sc_hd__a22o_2 _20897_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[4] ),
    .B1(_07771_),
    .B2(_07773_),
    .X(_01670_));
 sky130_fd_sc_hd__a22oi_2 _20898_ (.A1(\systolic_inst.A_outs[4][2] ),
    .A2(\systolic_inst.B_outs[4][3] ),
    .B1(\systolic_inst.B_outs[4][4] ),
    .B2(\systolic_inst.A_outs[4][1] ),
    .Y(_07774_));
 sky130_fd_sc_hd__and4_2 _20899_ (.A(\systolic_inst.A_outs[4][1] ),
    .B(\systolic_inst.A_outs[4][2] ),
    .C(\systolic_inst.B_outs[4][3] ),
    .D(\systolic_inst.B_outs[4][4] ),
    .X(_07775_));
 sky130_fd_sc_hd__or2_2 _20900_ (.A(_07774_),
    .B(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__xnor2_2 _20901_ (.A(_07759_),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__or2_2 _20902_ (.A(_07751_),
    .B(_07777_),
    .X(_07778_));
 sky130_fd_sc_hd__xnor2_2 _20903_ (.A(_07750_),
    .B(_07777_),
    .Y(_07779_));
 sky130_fd_sc_hd__nand4_2 _20904_ (.A(\systolic_inst.A_outs[4][0] ),
    .B(\systolic_inst.B_outs[4][1] ),
    .C(\systolic_inst.A_outs[4][4] ),
    .D(\systolic_inst.B_outs[4][5] ),
    .Y(_07780_));
 sky130_fd_sc_hd__a22o_2 _20905_ (.A1(\systolic_inst.B_outs[4][1] ),
    .A2(\systolic_inst.A_outs[4][4] ),
    .B1(\systolic_inst.B_outs[4][5] ),
    .B2(\systolic_inst.A_outs[4][0] ),
    .X(_07781_));
 sky130_fd_sc_hd__nand3b_2 _20906_ (.A_N(_07758_),
    .B(_07780_),
    .C(_07781_),
    .Y(_07782_));
 sky130_fd_sc_hd__a21bo_2 _20907_ (.A1(_07780_),
    .A2(_07781_),
    .B1_N(_07758_),
    .X(_07783_));
 sky130_fd_sc_hd__nand4_2 _20908_ (.A(\systolic_inst.B_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][5] ),
    .C(_07782_),
    .D(_07783_),
    .Y(_07784_));
 sky130_fd_sc_hd__a22o_2 _20909_ (.A1(\systolic_inst.B_outs[4][0] ),
    .A2(\systolic_inst.A_outs[4][5] ),
    .B1(_07782_),
    .B2(_07783_),
    .X(_07785_));
 sky130_fd_sc_hd__nand3_2 _20910_ (.A(_07760_),
    .B(_07784_),
    .C(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__a21o_2 _20911_ (.A1(_07784_),
    .A2(_07785_),
    .B1(_07760_),
    .X(_07787_));
 sky130_fd_sc_hd__nand3_2 _20912_ (.A(_07779_),
    .B(_07786_),
    .C(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__a21o_2 _20913_ (.A1(_07786_),
    .A2(_07787_),
    .B1(_07779_),
    .X(_07789_));
 sky130_fd_sc_hd__a21bo_2 _20914_ (.A1(_07756_),
    .A2(_07763_),
    .B1_N(_07762_),
    .X(_07790_));
 sky130_fd_sc_hd__nand3_2 _20915_ (.A(_07788_),
    .B(_07789_),
    .C(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__a21o_2 _20916_ (.A1(_07788_),
    .A2(_07789_),
    .B1(_07790_),
    .X(_07792_));
 sky130_fd_sc_hd__and3_2 _20917_ (.A(_07754_),
    .B(_07791_),
    .C(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__a21oi_2 _20918_ (.A1(_07791_),
    .A2(_07792_),
    .B1(_07754_),
    .Y(_07794_));
 sky130_fd_sc_hd__a31o_2 _20919_ (.A1(\systolic_inst.B_outs[4][3] ),
    .A2(_07729_),
    .A3(_07769_),
    .B1(_07767_),
    .X(_07795_));
 sky130_fd_sc_hd__nor3b_2 _20920_ (.A(_07793_),
    .B(_07794_),
    .C_N(_07795_),
    .Y(_07796_));
 sky130_fd_sc_hd__o21bai_2 _20921_ (.A1(_07793_),
    .A2(_07794_),
    .B1_N(_07795_),
    .Y(_07797_));
 sky130_fd_sc_hd__nand2b_2 _20922_ (.A_N(_07796_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__and3b_2 _20923_ (.A_N(_07796_),
    .B(_07797_),
    .C(_07772_),
    .X(_07799_));
 sky130_fd_sc_hd__xnor2_2 _20924_ (.A(_07772_),
    .B(_07798_),
    .Y(_07800_));
 sky130_fd_sc_hd__mux2_1 _20925_ (.A0(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[5] ),
    .A1(_07800_),
    .S(\systolic_inst.ce_local ),
    .X(_01671_));
 sky130_fd_sc_hd__o21a_2 _20926_ (.A1(_07759_),
    .A2(_07776_),
    .B1(_07778_),
    .X(_07801_));
 sky130_fd_sc_hd__nand2_2 _20927_ (.A(_07780_),
    .B(_07782_),
    .Y(_07802_));
 sky130_fd_sc_hd__a22oi_2 _20928_ (.A1(\systolic_inst.A_outs[4][3] ),
    .A2(\systolic_inst.B_outs[4][3] ),
    .B1(\systolic_inst.B_outs[4][4] ),
    .B2(\systolic_inst.A_outs[4][2] ),
    .Y(_07803_));
 sky130_fd_sc_hd__nand2_2 _20929_ (.A(\systolic_inst.A_outs[4][3] ),
    .B(\systolic_inst.B_outs[4][4] ),
    .Y(_07804_));
 sky130_fd_sc_hd__and4_2 _20930_ (.A(\systolic_inst.A_outs[4][2] ),
    .B(\systolic_inst.A_outs[4][3] ),
    .C(\systolic_inst.B_outs[4][3] ),
    .D(\systolic_inst.B_outs[4][4] ),
    .X(_07805_));
 sky130_fd_sc_hd__or2_2 _20931_ (.A(_07803_),
    .B(_07805_),
    .X(_07806_));
 sky130_fd_sc_hd__a21oi_2 _20932_ (.A1(_07780_),
    .A2(_07782_),
    .B1(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__xnor2_2 _20933_ (.A(_07802_),
    .B(_07806_),
    .Y(_07808_));
 sky130_fd_sc_hd__xnor2_2 _20934_ (.A(_07775_),
    .B(_07808_),
    .Y(_07809_));
 sky130_fd_sc_hd__nand2_2 _20935_ (.A(\systolic_inst.B_outs[4][2] ),
    .B(\systolic_inst.A_outs[4][4] ),
    .Y(_07810_));
 sky130_fd_sc_hd__nand4_2 _20936_ (.A(\systolic_inst.A_outs[4][1] ),
    .B(\systolic_inst.B_outs[4][1] ),
    .C(\systolic_inst.A_outs[4][5] ),
    .D(\systolic_inst.B_outs[4][5] ),
    .Y(_07811_));
 sky130_fd_sc_hd__a22o_2 _20937_ (.A1(\systolic_inst.B_outs[4][1] ),
    .A2(\systolic_inst.A_outs[4][5] ),
    .B1(\systolic_inst.B_outs[4][5] ),
    .B2(\systolic_inst.A_outs[4][1] ),
    .X(_07812_));
 sky130_fd_sc_hd__nand2_2 _20938_ (.A(_07811_),
    .B(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__xor2_2 _20939_ (.A(_07810_),
    .B(_07813_),
    .X(_07814_));
 sky130_fd_sc_hd__a22o_2 _20940_ (.A1(\systolic_inst.B_outs[4][0] ),
    .A2(\systolic_inst.A_outs[4][6] ),
    .B1(\systolic_inst.B_outs[4][6] ),
    .B2(\systolic_inst.A_outs[4][0] ),
    .X(_07815_));
 sky130_fd_sc_hd__inv_2 _20941_ (.A(_07815_),
    .Y(_07816_));
 sky130_fd_sc_hd__and4_2 _20942_ (.A(\systolic_inst.B_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][0] ),
    .C(\systolic_inst.A_outs[4][6] ),
    .D(\systolic_inst.B_outs[4][6] ),
    .X(_07817_));
 sky130_fd_sc_hd__nor2_2 _20943_ (.A(_07816_),
    .B(_07817_),
    .Y(_07818_));
 sky130_fd_sc_hd__xnor2_2 _20944_ (.A(_07814_),
    .B(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__or2_2 _20945_ (.A(_07784_),
    .B(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__xnor2_2 _20946_ (.A(_07784_),
    .B(_07819_),
    .Y(_07821_));
 sky130_fd_sc_hd__xor2_2 _20947_ (.A(_07809_),
    .B(_07821_),
    .X(_07822_));
 sky130_fd_sc_hd__nand2_2 _20948_ (.A(_07786_),
    .B(_07788_),
    .Y(_07823_));
 sky130_fd_sc_hd__xnor2_2 _20949_ (.A(_07822_),
    .B(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__nor2_2 _20950_ (.A(_07801_),
    .B(_07824_),
    .Y(_07825_));
 sky130_fd_sc_hd__xor2_2 _20951_ (.A(_07801_),
    .B(_07824_),
    .X(_07826_));
 sky130_fd_sc_hd__a31o_2 _20952_ (.A1(_07788_),
    .A2(_07789_),
    .A3(_07790_),
    .B1(_07793_),
    .X(_07827_));
 sky130_fd_sc_hd__and2_2 _20953_ (.A(_07826_),
    .B(_07827_),
    .X(_07828_));
 sky130_fd_sc_hd__nor2_2 _20954_ (.A(_07826_),
    .B(_07827_),
    .Y(_07829_));
 sky130_fd_sc_hd__nor2_2 _20955_ (.A(_07828_),
    .B(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__o21a_2 _20956_ (.A1(_07796_),
    .A2(_07799_),
    .B1(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__or3_2 _20957_ (.A(_07796_),
    .B(_07799_),
    .C(_07830_),
    .X(_07832_));
 sky130_fd_sc_hd__or3b_2 _20958_ (.A(_11258_),
    .B(_07831_),
    .C_N(_07832_),
    .X(_07833_));
 sky130_fd_sc_hd__a21bo_2 _20959_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[6] ),
    .B1_N(_07833_),
    .X(_01672_));
 sky130_fd_sc_hd__a21oi_2 _20960_ (.A1(_07822_),
    .A2(_07823_),
    .B1(_07825_),
    .Y(_07834_));
 sky130_fd_sc_hd__a21oi_2 _20961_ (.A1(_07775_),
    .A2(_07808_),
    .B1(_07807_),
    .Y(_07835_));
 sky130_fd_sc_hd__o21ai_2 _20962_ (.A1(_07810_),
    .A2(_07813_),
    .B1(_07811_),
    .Y(_07836_));
 sky130_fd_sc_hd__nand2_2 _20963_ (.A(\systolic_inst.B_outs[4][3] ),
    .B(\systolic_inst.A_outs[4][4] ),
    .Y(_07837_));
 sky130_fd_sc_hd__or2_2 _20964_ (.A(_07804_),
    .B(_07837_),
    .X(_07838_));
 sky130_fd_sc_hd__xor2_2 _20965_ (.A(_07804_),
    .B(_07837_),
    .X(_07839_));
 sky130_fd_sc_hd__xnor2_2 _20966_ (.A(\systolic_inst.B_outs[4][7] ),
    .B(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__nand2b_2 _20967_ (.A_N(_07840_),
    .B(_07836_),
    .Y(_07841_));
 sky130_fd_sc_hd__xnor2_2 _20968_ (.A(_07836_),
    .B(_07840_),
    .Y(_07842_));
 sky130_fd_sc_hd__xnor2_2 _20969_ (.A(_07805_),
    .B(_07842_),
    .Y(_07843_));
 sky130_fd_sc_hd__nand2_2 _20970_ (.A(\systolic_inst.B_outs[4][2] ),
    .B(\systolic_inst.A_outs[4][5] ),
    .Y(_07844_));
 sky130_fd_sc_hd__and3_2 _20971_ (.A(\systolic_inst.B_outs[4][1] ),
    .B(\systolic_inst.A_outs[4][2] ),
    .C(\systolic_inst.A_outs[4][6] ),
    .X(_07845_));
 sky130_fd_sc_hd__a22o_2 _20972_ (.A1(\systolic_inst.A_outs[4][2] ),
    .A2(\systolic_inst.B_outs[4][5] ),
    .B1(\systolic_inst.A_outs[4][6] ),
    .B2(\systolic_inst.B_outs[4][1] ),
    .X(_07846_));
 sky130_fd_sc_hd__a21bo_2 _20973_ (.A1(\systolic_inst.B_outs[4][5] ),
    .A2(_07845_),
    .B1_N(_07846_),
    .X(_07847_));
 sky130_fd_sc_hd__xor2_2 _20974_ (.A(_07844_),
    .B(_07847_),
    .X(_07848_));
 sky130_fd_sc_hd__nand2_2 _20975_ (.A(\systolic_inst.A_outs[4][1] ),
    .B(\systolic_inst.B_outs[4][6] ),
    .Y(_07849_));
 sky130_fd_sc_hd__nand2_2 _20976_ (.A(\systolic_inst.B_outs[4][0] ),
    .B(\systolic_inst.A_outs[4][7] ),
    .Y(_07850_));
 sky130_fd_sc_hd__and2b_2 _20977_ (.A_N(\systolic_inst.A_outs[4][0] ),
    .B(\systolic_inst.B_outs[4][7] ),
    .X(_07851_));
 sky130_fd_sc_hd__nand3_2 _20978_ (.A(\systolic_inst.B_outs[4][0] ),
    .B(\systolic_inst.B_outs[4][7] ),
    .C(\systolic_inst.A_outs[4][7] ),
    .Y(_07852_));
 sky130_fd_sc_hd__nor2_2 _20979_ (.A(\systolic_inst.A_outs[4][0] ),
    .B(_07852_),
    .Y(_07853_));
 sky130_fd_sc_hd__xnor2_2 _20980_ (.A(_07850_),
    .B(_07851_),
    .Y(_07854_));
 sky130_fd_sc_hd__xnor2_2 _20981_ (.A(_07849_),
    .B(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__and2_2 _20982_ (.A(_07817_),
    .B(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__xor2_2 _20983_ (.A(_07817_),
    .B(_07855_),
    .X(_07857_));
 sky130_fd_sc_hd__xnor2_2 _20984_ (.A(_07848_),
    .B(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__or4b_2 _20985_ (.A(_07816_),
    .B(_07817_),
    .C(_07858_),
    .D_N(_07814_),
    .X(_07859_));
 sky130_fd_sc_hd__a21bo_2 _20986_ (.A1(_07814_),
    .A2(_07818_),
    .B1_N(_07858_),
    .X(_07860_));
 sky130_fd_sc_hd__nand2_2 _20987_ (.A(_07859_),
    .B(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__xor2_2 _20988_ (.A(_07843_),
    .B(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__o21a_2 _20989_ (.A1(_07809_),
    .A2(_07821_),
    .B1(_07820_),
    .X(_07863_));
 sky130_fd_sc_hd__nand2b_2 _20990_ (.A_N(_07863_),
    .B(_07862_),
    .Y(_07864_));
 sky130_fd_sc_hd__xnor2_2 _20991_ (.A(_07862_),
    .B(_07863_),
    .Y(_07865_));
 sky130_fd_sc_hd__nand2b_2 _20992_ (.A_N(_07835_),
    .B(_07865_),
    .Y(_07866_));
 sky130_fd_sc_hd__xnor2_2 _20993_ (.A(_07835_),
    .B(_07865_),
    .Y(_07867_));
 sky130_fd_sc_hd__and2b_2 _20994_ (.A_N(_07834_),
    .B(_07867_),
    .X(_07868_));
 sky130_fd_sc_hd__xnor2_2 _20995_ (.A(_07834_),
    .B(_07867_),
    .Y(_07869_));
 sky130_fd_sc_hd__o21a_2 _20996_ (.A1(_07828_),
    .A2(_07831_),
    .B1(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__o31ai_2 _20997_ (.A1(_07828_),
    .A2(_07831_),
    .A3(_07869_),
    .B1(\systolic_inst.ce_local ),
    .Y(_07871_));
 sky130_fd_sc_hd__a2bb2o_2 _20998_ (.A1_N(_07871_),
    .A2_N(_07870_),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[7] ),
    .B2(_11258_),
    .X(_01673_));
 sky130_fd_sc_hd__a21bo_2 _20999_ (.A1(_07805_),
    .A2(_07842_),
    .B1_N(_07841_),
    .X(_07872_));
 sky130_fd_sc_hd__a21bo_2 _21000_ (.A1(\systolic_inst.B_outs[4][7] ),
    .A2(_07839_),
    .B1_N(_07838_),
    .X(_07873_));
 sky130_fd_sc_hd__a32o_2 _21001_ (.A1(\systolic_inst.B_outs[4][2] ),
    .A2(\systolic_inst.A_outs[4][5] ),
    .A3(_07846_),
    .B1(_07845_),
    .B2(\systolic_inst.B_outs[4][5] ),
    .X(_07874_));
 sky130_fd_sc_hd__a22o_2 _21002_ (.A1(\systolic_inst.A_outs[4][4] ),
    .A2(\systolic_inst.B_outs[4][4] ),
    .B1(\systolic_inst.A_outs[4][5] ),
    .B2(\systolic_inst.B_outs[4][3] ),
    .X(_07875_));
 sky130_fd_sc_hd__nand2_2 _21003_ (.A(\systolic_inst.B_outs[4][4] ),
    .B(\systolic_inst.A_outs[4][5] ),
    .Y(_07876_));
 sky130_fd_sc_hd__nor2_2 _21004_ (.A(_07837_),
    .B(_07876_),
    .Y(_07877_));
 sky130_fd_sc_hd__o21a_2 _21005_ (.A1(_07837_),
    .A2(_07876_),
    .B1(_07875_),
    .X(_07878_));
 sky130_fd_sc_hd__nand2_2 _21006_ (.A(_07874_),
    .B(_07878_),
    .Y(_07879_));
 sky130_fd_sc_hd__or2_2 _21007_ (.A(_07874_),
    .B(_07878_),
    .X(_07880_));
 sky130_fd_sc_hd__and2_2 _21008_ (.A(_07879_),
    .B(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__xnor2_2 _21009_ (.A(_07873_),
    .B(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__nand2_2 _21010_ (.A(\systolic_inst.B_outs[4][2] ),
    .B(\systolic_inst.A_outs[4][6] ),
    .Y(_07883_));
 sky130_fd_sc_hd__and3_2 _21011_ (.A(\systolic_inst.B_outs[4][1] ),
    .B(\systolic_inst.B_outs[4][5] ),
    .C(\systolic_inst.A_outs[4][7] ),
    .X(_07884_));
 sky130_fd_sc_hd__a22o_2 _21012_ (.A1(\systolic_inst.A_outs[4][3] ),
    .A2(\systolic_inst.B_outs[4][5] ),
    .B1(\systolic_inst.A_outs[4][7] ),
    .B2(\systolic_inst.B_outs[4][1] ),
    .X(_07885_));
 sky130_fd_sc_hd__a21bo_2 _21013_ (.A1(\systolic_inst.A_outs[4][3] ),
    .A2(_07884_),
    .B1_N(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__xor2_2 _21014_ (.A(_07883_),
    .B(_07886_),
    .X(_07887_));
 sky130_fd_sc_hd__nand2_2 _21015_ (.A(\systolic_inst.A_outs[4][2] ),
    .B(\systolic_inst.B_outs[4][6] ),
    .Y(_07888_));
 sky130_fd_sc_hd__and2b_2 _21016_ (.A_N(\systolic_inst.A_outs[4][1] ),
    .B(\systolic_inst.B_outs[4][7] ),
    .X(_07889_));
 sky130_fd_sc_hd__nor2_2 _21017_ (.A(\systolic_inst.A_outs[4][1] ),
    .B(_07852_),
    .Y(_07890_));
 sky130_fd_sc_hd__xnor2_2 _21018_ (.A(_07850_),
    .B(_07889_),
    .Y(_07891_));
 sky130_fd_sc_hd__xnor2_2 _21019_ (.A(_07888_),
    .B(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__a31o_2 _21020_ (.A1(\systolic_inst.A_outs[4][1] ),
    .A2(\systolic_inst.B_outs[4][6] ),
    .A3(_07854_),
    .B1(_07853_),
    .X(_07893_));
 sky130_fd_sc_hd__and2_2 _21021_ (.A(_07892_),
    .B(_07893_),
    .X(_07894_));
 sky130_fd_sc_hd__xor2_2 _21022_ (.A(_07892_),
    .B(_07893_),
    .X(_07895_));
 sky130_fd_sc_hd__xnor2_2 _21023_ (.A(_07887_),
    .B(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__a21oi_2 _21024_ (.A1(_07848_),
    .A2(_07857_),
    .B1(_07856_),
    .Y(_07897_));
 sky130_fd_sc_hd__xnor2_2 _21025_ (.A(_07896_),
    .B(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__nor2_2 _21026_ (.A(_07882_),
    .B(_07898_),
    .Y(_07899_));
 sky130_fd_sc_hd__and2_2 _21027_ (.A(_07882_),
    .B(_07898_),
    .X(_07900_));
 sky130_fd_sc_hd__nor2_2 _21028_ (.A(_07899_),
    .B(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__o21a_2 _21029_ (.A1(_07843_),
    .A2(_07861_),
    .B1(_07859_),
    .X(_07902_));
 sky130_fd_sc_hd__nand2b_2 _21030_ (.A_N(_07902_),
    .B(_07901_),
    .Y(_07903_));
 sky130_fd_sc_hd__xor2_2 _21031_ (.A(_07901_),
    .B(_07902_),
    .X(_07904_));
 sky130_fd_sc_hd__nand2b_2 _21032_ (.A_N(_07904_),
    .B(_07872_),
    .Y(_07905_));
 sky130_fd_sc_hd__xor2_2 _21033_ (.A(_07872_),
    .B(_07904_),
    .X(_07906_));
 sky130_fd_sc_hd__a21oi_2 _21034_ (.A1(_07864_),
    .A2(_07866_),
    .B1(_07906_),
    .Y(_07907_));
 sky130_fd_sc_hd__and3_2 _21035_ (.A(_07864_),
    .B(_07866_),
    .C(_07906_),
    .X(_07908_));
 sky130_fd_sc_hd__nor2_2 _21036_ (.A(_07907_),
    .B(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__o21a_2 _21037_ (.A1(_07868_),
    .A2(_07870_),
    .B1(_07909_),
    .X(_07910_));
 sky130_fd_sc_hd__nor3_2 _21038_ (.A(_07868_),
    .B(_07870_),
    .C(_07909_),
    .Y(_07911_));
 sky130_fd_sc_hd__nor2_2 _21039_ (.A(_07910_),
    .B(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__mux2_1 _21040_ (.A0(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[8] ),
    .A1(_07912_),
    .S(\systolic_inst.ce_local ),
    .X(_01674_));
 sky130_fd_sc_hd__a21bo_2 _21041_ (.A1(_07873_),
    .A2(_07880_),
    .B1_N(_07879_),
    .X(_07913_));
 sky130_fd_sc_hd__a32o_2 _21042_ (.A1(\systolic_inst.B_outs[4][2] ),
    .A2(\systolic_inst.A_outs[4][6] ),
    .A3(_07885_),
    .B1(_07884_),
    .B2(\systolic_inst.A_outs[4][3] ),
    .X(_07914_));
 sky130_fd_sc_hd__inv_2 _21043_ (.A(_07914_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_2 _21044_ (.A(\systolic_inst.B_outs[4][3] ),
    .B(\systolic_inst.A_outs[4][6] ),
    .Y(_07916_));
 sky130_fd_sc_hd__and4_2 _21045_ (.A(\systolic_inst.B_outs[4][3] ),
    .B(\systolic_inst.B_outs[4][4] ),
    .C(\systolic_inst.A_outs[4][5] ),
    .D(\systolic_inst.A_outs[4][6] ),
    .X(_07917_));
 sky130_fd_sc_hd__a21o_2 _21046_ (.A1(_07876_),
    .A2(_07916_),
    .B1(_07917_),
    .X(_07918_));
 sky130_fd_sc_hd__xnor2_2 _21047_ (.A(_07914_),
    .B(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__nand2_2 _21048_ (.A(_07877_),
    .B(_07919_),
    .Y(_07920_));
 sky130_fd_sc_hd__or2_2 _21049_ (.A(_07877_),
    .B(_07919_),
    .X(_07921_));
 sky130_fd_sc_hd__nand2_2 _21050_ (.A(_07920_),
    .B(_07921_),
    .Y(_07922_));
 sky130_fd_sc_hd__nand2_2 _21051_ (.A(\systolic_inst.B_outs[4][2] ),
    .B(\systolic_inst.A_outs[4][7] ),
    .Y(_07923_));
 sky130_fd_sc_hd__a22o_2 _21052_ (.A1(\systolic_inst.A_outs[4][4] ),
    .A2(\systolic_inst.B_outs[4][5] ),
    .B1(\systolic_inst.A_outs[4][7] ),
    .B2(\systolic_inst.B_outs[4][1] ),
    .X(_07924_));
 sky130_fd_sc_hd__a21bo_2 _21053_ (.A1(\systolic_inst.A_outs[4][4] ),
    .A2(_07884_),
    .B1_N(_07924_),
    .X(_07925_));
 sky130_fd_sc_hd__xor2_2 _21054_ (.A(_07923_),
    .B(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__nand2_2 _21055_ (.A(\systolic_inst.A_outs[4][3] ),
    .B(\systolic_inst.B_outs[4][6] ),
    .Y(_07927_));
 sky130_fd_sc_hd__o21ai_2 _21056_ (.A1(\systolic_inst.A_outs[4][2] ),
    .A2(_11271_),
    .B1(_07850_),
    .Y(_07928_));
 sky130_fd_sc_hd__nor2_2 _21057_ (.A(\systolic_inst.A_outs[4][2] ),
    .B(_07852_),
    .Y(_07929_));
 sky130_fd_sc_hd__o21a_2 _21058_ (.A1(\systolic_inst.A_outs[4][2] ),
    .A2(_07852_),
    .B1(_07928_),
    .X(_07930_));
 sky130_fd_sc_hd__xnor2_2 _21059_ (.A(_07927_),
    .B(_07930_),
    .Y(_07931_));
 sky130_fd_sc_hd__a31o_2 _21060_ (.A1(\systolic_inst.A_outs[4][2] ),
    .A2(\systolic_inst.B_outs[4][6] ),
    .A3(_07891_),
    .B1(_07890_),
    .X(_07932_));
 sky130_fd_sc_hd__and2_2 _21061_ (.A(_07931_),
    .B(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__xor2_2 _21062_ (.A(_07931_),
    .B(_07932_),
    .X(_07934_));
 sky130_fd_sc_hd__xnor2_2 _21063_ (.A(_07926_),
    .B(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__a21o_2 _21064_ (.A1(_07887_),
    .A2(_07895_),
    .B1(_07894_),
    .X(_07936_));
 sky130_fd_sc_hd__and2b_2 _21065_ (.A_N(_07935_),
    .B(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__xor2_2 _21066_ (.A(_07935_),
    .B(_07936_),
    .X(_07938_));
 sky130_fd_sc_hd__nor2_2 _21067_ (.A(_07922_),
    .B(_07938_),
    .Y(_07939_));
 sky130_fd_sc_hd__and2_2 _21068_ (.A(_07922_),
    .B(_07938_),
    .X(_07940_));
 sky130_fd_sc_hd__nor2_2 _21069_ (.A(_07939_),
    .B(_07940_),
    .Y(_07941_));
 sky130_fd_sc_hd__o21ba_2 _21070_ (.A1(_07896_),
    .A2(_07897_),
    .B1_N(_07899_),
    .X(_07942_));
 sky130_fd_sc_hd__nand2b_2 _21071_ (.A_N(_07942_),
    .B(_07941_),
    .Y(_07943_));
 sky130_fd_sc_hd__xnor2_2 _21072_ (.A(_07941_),
    .B(_07942_),
    .Y(_07944_));
 sky130_fd_sc_hd__xnor2_2 _21073_ (.A(_07913_),
    .B(_07944_),
    .Y(_07945_));
 sky130_fd_sc_hd__a21oi_2 _21074_ (.A1(_07903_),
    .A2(_07905_),
    .B1(_07945_),
    .Y(_07946_));
 sky130_fd_sc_hd__and3_2 _21075_ (.A(_07903_),
    .B(_07905_),
    .C(_07945_),
    .X(_07947_));
 sky130_fd_sc_hd__inv_2 _21076_ (.A(_07947_),
    .Y(_07948_));
 sky130_fd_sc_hd__nor2_2 _21077_ (.A(_07946_),
    .B(_07947_),
    .Y(_07949_));
 sky130_fd_sc_hd__nor2_2 _21078_ (.A(_07907_),
    .B(_07910_),
    .Y(_07950_));
 sky130_fd_sc_hd__xnor2_2 _21079_ (.A(_07949_),
    .B(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__mux2_1 _21080_ (.A0(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[9] ),
    .A1(_07951_),
    .S(\systolic_inst.ce_local ),
    .X(_01675_));
 sky130_fd_sc_hd__o21ai_2 _21081_ (.A1(_07915_),
    .A2(_07918_),
    .B1(_07920_),
    .Y(_07952_));
 sky130_fd_sc_hd__a32o_2 _21082_ (.A1(\systolic_inst.B_outs[4][2] ),
    .A2(\systolic_inst.A_outs[4][7] ),
    .A3(_07924_),
    .B1(_07884_),
    .B2(\systolic_inst.A_outs[4][4] ),
    .X(_07953_));
 sky130_fd_sc_hd__a22o_2 _21083_ (.A1(\systolic_inst.B_outs[4][4] ),
    .A2(\systolic_inst.A_outs[4][6] ),
    .B1(\systolic_inst.A_outs[4][7] ),
    .B2(\systolic_inst.B_outs[4][3] ),
    .X(_07954_));
 sky130_fd_sc_hd__and4_2 _21084_ (.A(\systolic_inst.B_outs[4][3] ),
    .B(\systolic_inst.B_outs[4][4] ),
    .C(\systolic_inst.A_outs[4][6] ),
    .D(\systolic_inst.A_outs[4][7] ),
    .X(_07955_));
 sky130_fd_sc_hd__nand4_2 _21085_ (.A(\systolic_inst.B_outs[4][3] ),
    .B(\systolic_inst.B_outs[4][4] ),
    .C(\systolic_inst.A_outs[4][6] ),
    .D(\systolic_inst.A_outs[4][7] ),
    .Y(_07956_));
 sky130_fd_sc_hd__nand2_2 _21086_ (.A(_07954_),
    .B(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__xnor2_2 _21087_ (.A(_07953_),
    .B(_07957_),
    .Y(_07958_));
 sky130_fd_sc_hd__xnor2_2 _21088_ (.A(_07917_),
    .B(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__a22o_2 _21089_ (.A1(\systolic_inst.A_outs[4][5] ),
    .A2(\systolic_inst.B_outs[4][5] ),
    .B1(\systolic_inst.A_outs[4][7] ),
    .B2(\systolic_inst.B_outs[4][1] ),
    .X(_07960_));
 sky130_fd_sc_hd__a21bo_2 _21090_ (.A1(\systolic_inst.A_outs[4][5] ),
    .A2(_07884_),
    .B1_N(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__xor2_2 _21091_ (.A(_07923_),
    .B(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__nand2_2 _21092_ (.A(\systolic_inst.A_outs[4][4] ),
    .B(\systolic_inst.B_outs[4][6] ),
    .Y(_07963_));
 sky130_fd_sc_hd__o21ai_2 _21093_ (.A1(\systolic_inst.A_outs[4][3] ),
    .A2(_11271_),
    .B1(_07850_),
    .Y(_07964_));
 sky130_fd_sc_hd__nor2_2 _21094_ (.A(\systolic_inst.A_outs[4][3] ),
    .B(_07852_),
    .Y(_07965_));
 sky130_fd_sc_hd__o21a_2 _21095_ (.A1(\systolic_inst.A_outs[4][3] ),
    .A2(_07852_),
    .B1(_07964_),
    .X(_07966_));
 sky130_fd_sc_hd__xnor2_2 _21096_ (.A(_07963_),
    .B(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__a31o_2 _21097_ (.A1(\systolic_inst.A_outs[4][3] ),
    .A2(\systolic_inst.B_outs[4][6] ),
    .A3(_07928_),
    .B1(_07929_),
    .X(_07968_));
 sky130_fd_sc_hd__and2_2 _21098_ (.A(_07967_),
    .B(_07968_),
    .X(_07969_));
 sky130_fd_sc_hd__xor2_2 _21099_ (.A(_07967_),
    .B(_07968_),
    .X(_07970_));
 sky130_fd_sc_hd__xnor2_2 _21100_ (.A(_07962_),
    .B(_07970_),
    .Y(_07971_));
 sky130_fd_sc_hd__a21o_2 _21101_ (.A1(_07926_),
    .A2(_07934_),
    .B1(_07933_),
    .X(_07972_));
 sky130_fd_sc_hd__and2b_2 _21102_ (.A_N(_07971_),
    .B(_07972_),
    .X(_07973_));
 sky130_fd_sc_hd__xor2_2 _21103_ (.A(_07971_),
    .B(_07972_),
    .X(_07974_));
 sky130_fd_sc_hd__xor2_2 _21104_ (.A(_07959_),
    .B(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__o21ai_2 _21105_ (.A1(_07937_),
    .A2(_07939_),
    .B1(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__or3_2 _21106_ (.A(_07937_),
    .B(_07939_),
    .C(_07975_),
    .X(_07977_));
 sky130_fd_sc_hd__and2_2 _21107_ (.A(_07976_),
    .B(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__nand2_2 _21108_ (.A(_07952_),
    .B(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__xnor2_2 _21109_ (.A(_07952_),
    .B(_07978_),
    .Y(_07980_));
 sky130_fd_sc_hd__a21boi_2 _21110_ (.A1(_07913_),
    .A2(_07944_),
    .B1_N(_07943_),
    .Y(_07981_));
 sky130_fd_sc_hd__nor2_2 _21111_ (.A(_07980_),
    .B(_07981_),
    .Y(_07982_));
 sky130_fd_sc_hd__xnor2_2 _21112_ (.A(_07980_),
    .B(_07981_),
    .Y(_07983_));
 sky130_fd_sc_hd__inv_2 _21113_ (.A(_07983_),
    .Y(_07984_));
 sky130_fd_sc_hd__o31a_2 _21114_ (.A1(_07907_),
    .A2(_07910_),
    .A3(_07946_),
    .B1(_07948_),
    .X(_07985_));
 sky130_fd_sc_hd__o311a_2 _21115_ (.A1(_07907_),
    .A2(_07910_),
    .A3(_07946_),
    .B1(_07948_),
    .C1(_07984_),
    .X(_07986_));
 sky130_fd_sc_hd__xnor2_2 _21116_ (.A(_07983_),
    .B(_07985_),
    .Y(_07987_));
 sky130_fd_sc_hd__mux2_1 _21117_ (.A0(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[10] ),
    .A1(_07987_),
    .S(\systolic_inst.ce_local ),
    .X(_01676_));
 sky130_fd_sc_hd__a32o_2 _21118_ (.A1(_07953_),
    .A2(_07954_),
    .A3(_07956_),
    .B1(_07958_),
    .B2(_07917_),
    .X(_07988_));
 sky130_fd_sc_hd__a32o_2 _21119_ (.A1(\systolic_inst.B_outs[4][2] ),
    .A2(\systolic_inst.A_outs[4][7] ),
    .A3(_07960_),
    .B1(_07884_),
    .B2(\systolic_inst.A_outs[4][5] ),
    .X(_07989_));
 sky130_fd_sc_hd__inv_2 _21120_ (.A(_07989_),
    .Y(_07990_));
 sky130_fd_sc_hd__o21a_2 _21121_ (.A1(\systolic_inst.B_outs[4][3] ),
    .A2(\systolic_inst.B_outs[4][4] ),
    .B1(\systolic_inst.A_outs[4][7] ),
    .X(_07991_));
 sky130_fd_sc_hd__o21ai_2 _21122_ (.A1(\systolic_inst.B_outs[4][3] ),
    .A2(\systolic_inst.B_outs[4][4] ),
    .B1(\systolic_inst.A_outs[4][7] ),
    .Y(_07992_));
 sky130_fd_sc_hd__a21o_2 _21123_ (.A1(\systolic_inst.B_outs[4][3] ),
    .A2(\systolic_inst.B_outs[4][4] ),
    .B1(_07992_),
    .X(_07993_));
 sky130_fd_sc_hd__xnor2_2 _21124_ (.A(_07989_),
    .B(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__or2_2 _21125_ (.A(_07955_),
    .B(_07994_),
    .X(_07995_));
 sky130_fd_sc_hd__nand2_2 _21126_ (.A(_07955_),
    .B(_07994_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand2_2 _21127_ (.A(_07995_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__a22o_2 _21128_ (.A1(\systolic_inst.B_outs[4][5] ),
    .A2(\systolic_inst.A_outs[4][6] ),
    .B1(\systolic_inst.A_outs[4][7] ),
    .B2(\systolic_inst.B_outs[4][1] ),
    .X(_07998_));
 sky130_fd_sc_hd__a21bo_2 _21129_ (.A1(\systolic_inst.A_outs[4][6] ),
    .A2(_07884_),
    .B1_N(_07998_),
    .X(_07999_));
 sky130_fd_sc_hd__xor2_2 _21130_ (.A(_07923_),
    .B(_07999_),
    .X(_08000_));
 sky130_fd_sc_hd__o21a_2 _21131_ (.A1(\systolic_inst.A_outs[4][4] ),
    .A2(_11271_),
    .B1(_07850_),
    .X(_08001_));
 sky130_fd_sc_hd__nor2_2 _21132_ (.A(\systolic_inst.A_outs[4][4] ),
    .B(_07852_),
    .Y(_08002_));
 sky130_fd_sc_hd__nor2_2 _21133_ (.A(_08001_),
    .B(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__and3_2 _21134_ (.A(\systolic_inst.A_outs[4][5] ),
    .B(\systolic_inst.B_outs[4][6] ),
    .C(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__a21oi_2 _21135_ (.A1(\systolic_inst.A_outs[4][5] ),
    .A2(\systolic_inst.B_outs[4][6] ),
    .B1(_08003_),
    .Y(_08005_));
 sky130_fd_sc_hd__nor2_2 _21136_ (.A(_08004_),
    .B(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__a31o_2 _21137_ (.A1(\systolic_inst.A_outs[4][4] ),
    .A2(\systolic_inst.B_outs[4][6] ),
    .A3(_07964_),
    .B1(_07965_),
    .X(_08007_));
 sky130_fd_sc_hd__and2_2 _21138_ (.A(_08006_),
    .B(_08007_),
    .X(_08008_));
 sky130_fd_sc_hd__nor2_2 _21139_ (.A(_08006_),
    .B(_08007_),
    .Y(_08009_));
 sky130_fd_sc_hd__nor2_2 _21140_ (.A(_08008_),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__xnor2_2 _21141_ (.A(_08000_),
    .B(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__a21o_2 _21142_ (.A1(_07962_),
    .A2(_07970_),
    .B1(_07969_),
    .X(_08012_));
 sky130_fd_sc_hd__and2b_2 _21143_ (.A_N(_08011_),
    .B(_08012_),
    .X(_08013_));
 sky130_fd_sc_hd__xor2_2 _21144_ (.A(_08011_),
    .B(_08012_),
    .X(_08014_));
 sky130_fd_sc_hd__xor2_2 _21145_ (.A(_07997_),
    .B(_08014_),
    .X(_08015_));
 sky130_fd_sc_hd__o21ba_2 _21146_ (.A1(_07959_),
    .A2(_07974_),
    .B1_N(_07973_),
    .X(_08016_));
 sky130_fd_sc_hd__nand2b_2 _21147_ (.A_N(_08016_),
    .B(_08015_),
    .Y(_08017_));
 sky130_fd_sc_hd__xnor2_2 _21148_ (.A(_08015_),
    .B(_08016_),
    .Y(_08018_));
 sky130_fd_sc_hd__xnor2_2 _21149_ (.A(_07988_),
    .B(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand3_2 _21150_ (.A(_07976_),
    .B(_07979_),
    .C(_08019_),
    .Y(_08020_));
 sky130_fd_sc_hd__inv_2 _21151_ (.A(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__a21oi_2 _21152_ (.A1(_07976_),
    .A2(_07979_),
    .B1(_08019_),
    .Y(_08022_));
 sky130_fd_sc_hd__nor2_2 _21153_ (.A(_08021_),
    .B(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__nor2_2 _21154_ (.A(_07982_),
    .B(_07986_),
    .Y(_08024_));
 sky130_fd_sc_hd__xnor2_2 _21155_ (.A(_08023_),
    .B(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__mux2_1 _21156_ (.A0(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[11] ),
    .A1(_08025_),
    .S(\systolic_inst.ce_local ),
    .X(_01677_));
 sky130_fd_sc_hd__o21ai_2 _21157_ (.A1(_07990_),
    .A2(_07993_),
    .B1(_07996_),
    .Y(_08026_));
 sky130_fd_sc_hd__o2bb2a_2 _21158_ (.A1_N(\systolic_inst.A_outs[4][6] ),
    .A2_N(_07884_),
    .B1(_07923_),
    .B2(_07999_),
    .X(_08027_));
 sky130_fd_sc_hd__nor2_2 _21159_ (.A(_07992_),
    .B(_08027_),
    .Y(_08028_));
 sky130_fd_sc_hd__and2_2 _21160_ (.A(_07992_),
    .B(_08027_),
    .X(_08029_));
 sky130_fd_sc_hd__nor2_2 _21161_ (.A(_08028_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__o21a_2 _21162_ (.A1(\systolic_inst.A_outs[4][5] ),
    .A2(_11271_),
    .B1(_07850_),
    .X(_08031_));
 sky130_fd_sc_hd__nor2_2 _21163_ (.A(\systolic_inst.A_outs[4][5] ),
    .B(_07852_),
    .Y(_08032_));
 sky130_fd_sc_hd__nor2_2 _21164_ (.A(_08031_),
    .B(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__nand2_2 _21165_ (.A(\systolic_inst.A_outs[4][6] ),
    .B(\systolic_inst.B_outs[4][6] ),
    .Y(_08034_));
 sky130_fd_sc_hd__xnor2_2 _21166_ (.A(_08033_),
    .B(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__o21ai_2 _21167_ (.A1(_08002_),
    .A2(_08004_),
    .B1(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__or3_2 _21168_ (.A(_08002_),
    .B(_08004_),
    .C(_08035_),
    .X(_08037_));
 sky130_fd_sc_hd__nand2_2 _21169_ (.A(_08036_),
    .B(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__or2_2 _21170_ (.A(\systolic_inst.B_outs[4][1] ),
    .B(\systolic_inst.B_outs[4][5] ),
    .X(_08039_));
 sky130_fd_sc_hd__and3b_2 _21171_ (.A_N(_07884_),
    .B(_08039_),
    .C(\systolic_inst.A_outs[4][7] ),
    .X(_08040_));
 sky130_fd_sc_hd__xor2_2 _21172_ (.A(_07923_),
    .B(_08040_),
    .X(_08041_));
 sky130_fd_sc_hd__nand2_2 _21173_ (.A(_08038_),
    .B(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__or2_2 _21174_ (.A(_08038_),
    .B(_08041_),
    .X(_08043_));
 sky130_fd_sc_hd__nand2_2 _21175_ (.A(_08042_),
    .B(_08043_),
    .Y(_08044_));
 sky130_fd_sc_hd__a21o_2 _21176_ (.A1(_08000_),
    .A2(_08010_),
    .B1(_08008_),
    .X(_08045_));
 sky130_fd_sc_hd__xnor2_2 _21177_ (.A(_08044_),
    .B(_08045_),
    .Y(_08046_));
 sky130_fd_sc_hd__xor2_2 _21178_ (.A(_08030_),
    .B(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__o21ba_2 _21179_ (.A1(_07997_),
    .A2(_08014_),
    .B1_N(_08013_),
    .X(_08048_));
 sky130_fd_sc_hd__nand2b_2 _21180_ (.A_N(_08048_),
    .B(_08047_),
    .Y(_08049_));
 sky130_fd_sc_hd__xor2_2 _21181_ (.A(_08047_),
    .B(_08048_),
    .X(_08050_));
 sky130_fd_sc_hd__nand2b_2 _21182_ (.A_N(_08050_),
    .B(_08026_),
    .Y(_08051_));
 sky130_fd_sc_hd__xor2_2 _21183_ (.A(_08026_),
    .B(_08050_),
    .X(_08052_));
 sky130_fd_sc_hd__a21boi_2 _21184_ (.A1(_07988_),
    .A2(_08018_),
    .B1_N(_08017_),
    .Y(_08053_));
 sky130_fd_sc_hd__xnor2_2 _21185_ (.A(_08052_),
    .B(_08053_),
    .Y(_08054_));
 sky130_fd_sc_hd__inv_2 _21186_ (.A(_08054_),
    .Y(_08055_));
 sky130_fd_sc_hd__o31a_2 _21187_ (.A1(_07982_),
    .A2(_07986_),
    .A3(_08022_),
    .B1(_08020_),
    .X(_08056_));
 sky130_fd_sc_hd__o311a_2 _21188_ (.A1(_07982_),
    .A2(_07986_),
    .A3(_08022_),
    .B1(_08055_),
    .C1(_08020_),
    .X(_08057_));
 sky130_fd_sc_hd__nor2_2 _21189_ (.A(_08055_),
    .B(_08056_),
    .Y(_08058_));
 sky130_fd_sc_hd__nor2_2 _21190_ (.A(_08057_),
    .B(_08058_),
    .Y(_08059_));
 sky130_fd_sc_hd__mux2_1 _21191_ (.A0(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[12] ),
    .A1(_08059_),
    .S(\systolic_inst.ce_local ),
    .X(_01678_));
 sky130_fd_sc_hd__o21a_2 _21192_ (.A1(\systolic_inst.A_outs[4][6] ),
    .A2(_11271_),
    .B1(_07850_),
    .X(_08060_));
 sky130_fd_sc_hd__o21ba_2 _21193_ (.A1(\systolic_inst.A_outs[4][6] ),
    .A2(_07852_),
    .B1_N(_08060_),
    .X(_08061_));
 sky130_fd_sc_hd__nand2_2 _21194_ (.A(\systolic_inst.B_outs[4][6] ),
    .B(\systolic_inst.A_outs[4][7] ),
    .Y(_08062_));
 sky130_fd_sc_hd__xor2_2 _21195_ (.A(_08061_),
    .B(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__o21ba_2 _21196_ (.A1(_08031_),
    .A2(_08034_),
    .B1_N(_08032_),
    .X(_08064_));
 sky130_fd_sc_hd__xnor2_2 _21197_ (.A(_08063_),
    .B(_08064_),
    .Y(_08065_));
 sky130_fd_sc_hd__nor2_2 _21198_ (.A(_08041_),
    .B(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__and2_2 _21199_ (.A(_08041_),
    .B(_08065_),
    .X(_08067_));
 sky130_fd_sc_hd__or2_2 _21200_ (.A(_08066_),
    .B(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__a21oi_2 _21201_ (.A1(_08036_),
    .A2(_08043_),
    .B1(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__and3_2 _21202_ (.A(_08036_),
    .B(_08043_),
    .C(_08068_),
    .X(_08070_));
 sky130_fd_sc_hd__or2_2 _21203_ (.A(_08069_),
    .B(_08070_),
    .X(_08071_));
 sky130_fd_sc_hd__a31o_2 _21204_ (.A1(\systolic_inst.B_outs[4][2] ),
    .A2(\systolic_inst.A_outs[4][7] ),
    .A3(_08039_),
    .B1(_07884_),
    .X(_08072_));
 sky130_fd_sc_hd__nand2_2 _21205_ (.A(_07991_),
    .B(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__xnor2_2 _21206_ (.A(_07991_),
    .B(_08072_),
    .Y(_08074_));
 sky130_fd_sc_hd__and2_2 _21207_ (.A(_08071_),
    .B(_08074_),
    .X(_08075_));
 sky130_fd_sc_hd__nor2_2 _21208_ (.A(_08071_),
    .B(_08074_),
    .Y(_08076_));
 sky130_fd_sc_hd__or2_2 _21209_ (.A(_08075_),
    .B(_08076_),
    .X(_08077_));
 sky130_fd_sc_hd__a32o_2 _21210_ (.A1(_08042_),
    .A2(_08043_),
    .A3(_08045_),
    .B1(_08046_),
    .B2(_08030_),
    .X(_08078_));
 sky130_fd_sc_hd__nand2b_2 _21211_ (.A_N(_08077_),
    .B(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__xnor2_2 _21212_ (.A(_08077_),
    .B(_08078_),
    .Y(_08080_));
 sky130_fd_sc_hd__nand2_2 _21213_ (.A(_08028_),
    .B(_08080_),
    .Y(_08081_));
 sky130_fd_sc_hd__xnor2_2 _21214_ (.A(_08028_),
    .B(_08080_),
    .Y(_08082_));
 sky130_fd_sc_hd__and3_2 _21215_ (.A(_08049_),
    .B(_08051_),
    .C(_08082_),
    .X(_08083_));
 sky130_fd_sc_hd__a21o_2 _21216_ (.A1(_08049_),
    .A2(_08051_),
    .B1(_08082_),
    .X(_08084_));
 sky130_fd_sc_hd__and2b_2 _21217_ (.A_N(_08083_),
    .B(_08084_),
    .X(_08085_));
 sky130_fd_sc_hd__o21ba_2 _21218_ (.A1(_08052_),
    .A2(_08053_),
    .B1_N(_08057_),
    .X(_08086_));
 sky130_fd_sc_hd__xnor2_2 _21219_ (.A(_08085_),
    .B(_08086_),
    .Y(_08087_));
 sky130_fd_sc_hd__mux2_1 _21220_ (.A0(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[13] ),
    .A1(_08087_),
    .S(\systolic_inst.ce_local ),
    .X(_01679_));
 sky130_fd_sc_hd__and2_2 _21221_ (.A(_11258_),
    .B(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[14] ),
    .X(_08088_));
 sky130_fd_sc_hd__o211a_2 _21222_ (.A1(_11271_),
    .A2(\systolic_inst.A_outs[4][7] ),
    .B1(_07850_),
    .C1(_08062_),
    .X(_08089_));
 sky130_fd_sc_hd__o22a_2 _21223_ (.A1(\systolic_inst.A_outs[4][6] ),
    .A2(_07852_),
    .B1(_08060_),
    .B2(_08062_),
    .X(_08090_));
 sky130_fd_sc_hd__a31oi_2 _21224_ (.A1(\systolic_inst.B_outs[4][0] ),
    .A2(\systolic_inst.B_outs[4][6] ),
    .A3(\systolic_inst.A_outs[4][7] ),
    .B1(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__or3_2 _21225_ (.A(_08041_),
    .B(_08089_),
    .C(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__o21ai_2 _21226_ (.A1(_08089_),
    .A2(_08091_),
    .B1(_08041_),
    .Y(_08093_));
 sky130_fd_sc_hd__nand2_2 _21227_ (.A(_08092_),
    .B(_08093_),
    .Y(_08094_));
 sky130_fd_sc_hd__o21ba_2 _21228_ (.A1(_08063_),
    .A2(_08064_),
    .B1_N(_08066_),
    .X(_08095_));
 sky130_fd_sc_hd__xnor2_2 _21229_ (.A(_08094_),
    .B(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__or2_2 _21230_ (.A(_08074_),
    .B(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__nand2_2 _21231_ (.A(_08074_),
    .B(_08096_),
    .Y(_08098_));
 sky130_fd_sc_hd__and2_2 _21232_ (.A(_08097_),
    .B(_08098_),
    .X(_08099_));
 sky130_fd_sc_hd__or3_2 _21233_ (.A(_08069_),
    .B(_08076_),
    .C(_08099_),
    .X(_08100_));
 sky130_fd_sc_hd__o21ai_2 _21234_ (.A1(_08069_),
    .A2(_08076_),
    .B1(_08099_),
    .Y(_08101_));
 sky130_fd_sc_hd__nand2_2 _21235_ (.A(_08100_),
    .B(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__xnor2_2 _21236_ (.A(_08073_),
    .B(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__a21oi_2 _21237_ (.A1(_08079_),
    .A2(_08081_),
    .B1(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__and3_2 _21238_ (.A(_08079_),
    .B(_08081_),
    .C(_08103_),
    .X(_08105_));
 sky130_fd_sc_hd__or2_2 _21239_ (.A(_08104_),
    .B(_08105_),
    .X(_08106_));
 sky130_fd_sc_hd__nand2_2 _21240_ (.A(_08057_),
    .B(_08085_),
    .Y(_08107_));
 sky130_fd_sc_hd__or3_2 _21241_ (.A(_08052_),
    .B(_08053_),
    .C(_08083_),
    .X(_08108_));
 sky130_fd_sc_hd__nand4_2 _21242_ (.A(_08084_),
    .B(_08106_),
    .C(_08107_),
    .D(_08108_),
    .Y(_08109_));
 sky130_fd_sc_hd__a31o_2 _21243_ (.A1(_08084_),
    .A2(_08107_),
    .A3(_08108_),
    .B1(_08106_),
    .X(_08110_));
 sky130_fd_sc_hd__a31o_2 _21244_ (.A1(\systolic_inst.ce_local ),
    .A2(_08109_),
    .A3(_08110_),
    .B1(_08088_),
    .X(_01680_));
 sky130_fd_sc_hd__xor2_2 _21245_ (.A(_08074_),
    .B(_08093_),
    .X(_08111_));
 sky130_fd_sc_hd__o21a_2 _21246_ (.A1(_08094_),
    .A2(_08095_),
    .B1(_08097_),
    .X(_08112_));
 sky130_fd_sc_hd__xnor2_2 _21247_ (.A(_08111_),
    .B(_08112_),
    .Y(_08113_));
 sky130_fd_sc_hd__mux2_1 _21248_ (.A0(_08100_),
    .A1(_08101_),
    .S(_08073_),
    .X(_08114_));
 sky130_fd_sc_hd__o21ai_2 _21249_ (.A1(_08113_),
    .A2(_08114_),
    .B1(\systolic_inst.ce_local ),
    .Y(_08115_));
 sky130_fd_sc_hd__a211oi_2 _21250_ (.A1(_08113_),
    .A2(_08114_),
    .B1(_08115_),
    .C1(_08104_),
    .Y(_08116_));
 sky130_fd_sc_hd__a22o_2 _21251_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B1(_08110_),
    .B2(_08116_),
    .X(_01681_));
 sky130_fd_sc_hd__a21o_2 _21252_ (.A1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[4][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_08117_));
 sky130_fd_sc_hd__a21oi_2 _21253_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[4][0] ),
    .Y(_08118_));
 sky130_fd_sc_hd__a21oi_2 _21254_ (.A1(\systolic_inst.ce_local ),
    .A2(_08117_),
    .B1(_08118_),
    .Y(_01682_));
 sky130_fd_sc_hd__and2_2 _21255_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[4][1] ),
    .X(_08119_));
 sky130_fd_sc_hd__nand2_2 _21256_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[4][1] ),
    .Y(_08120_));
 sky130_fd_sc_hd__or2_2 _21257_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[4][1] ),
    .X(_08121_));
 sky130_fd_sc_hd__and4_2 _21258_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[4][0] ),
    .C(_08120_),
    .D(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__inv_2 _21259_ (.A(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__a22o_2 _21260_ (.A1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[4][0] ),
    .B1(_08120_),
    .B2(_08121_),
    .X(_08124_));
 sky130_fd_sc_hd__a32o_2 _21261_ (.A1(_11712_),
    .A2(_08123_),
    .A3(_08124_),
    .B1(\systolic_inst.acc_wires[4][1] ),
    .B2(_11258_),
    .X(_01683_));
 sky130_fd_sc_hd__and2_2 _21262_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[4][2] ),
    .X(_08125_));
 sky130_fd_sc_hd__nand2_2 _21263_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[4][2] ),
    .Y(_08126_));
 sky130_fd_sc_hd__or2_2 _21264_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[4][2] ),
    .X(_08127_));
 sky130_fd_sc_hd__a211o_2 _21265_ (.A1(_08126_),
    .A2(_08127_),
    .B1(_08119_),
    .C1(_08122_),
    .X(_08128_));
 sky130_fd_sc_hd__o211a_2 _21266_ (.A1(_08119_),
    .A2(_08122_),
    .B1(_08126_),
    .C1(_08127_),
    .X(_08129_));
 sky130_fd_sc_hd__inv_2 _21267_ (.A(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__a32o_2 _21268_ (.A1(_11712_),
    .A2(_08128_),
    .A3(_08130_),
    .B1(\systolic_inst.acc_wires[4][2] ),
    .B2(_11258_),
    .X(_01684_));
 sky130_fd_sc_hd__and2_2 _21269_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[4][3] ),
    .X(_08131_));
 sky130_fd_sc_hd__nand2_2 _21270_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[4][3] ),
    .Y(_08132_));
 sky130_fd_sc_hd__or2_2 _21271_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[4][3] ),
    .X(_08133_));
 sky130_fd_sc_hd__a211o_2 _21272_ (.A1(_08132_),
    .A2(_08133_),
    .B1(_08125_),
    .C1(_08129_),
    .X(_08134_));
 sky130_fd_sc_hd__o211a_2 _21273_ (.A1(_08125_),
    .A2(_08129_),
    .B1(_08132_),
    .C1(_08133_),
    .X(_08135_));
 sky130_fd_sc_hd__inv_2 _21274_ (.A(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__a32o_2 _21275_ (.A1(_11712_),
    .A2(_08134_),
    .A3(_08136_),
    .B1(\systolic_inst.acc_wires[4][3] ),
    .B2(_11258_),
    .X(_01685_));
 sky130_fd_sc_hd__and2_2 _21276_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[4][4] ),
    .X(_08137_));
 sky130_fd_sc_hd__nand2_2 _21277_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[4][4] ),
    .Y(_08138_));
 sky130_fd_sc_hd__or2_2 _21278_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[4][4] ),
    .X(_08139_));
 sky130_fd_sc_hd__a211o_2 _21279_ (.A1(_08138_),
    .A2(_08139_),
    .B1(_08131_),
    .C1(_08135_),
    .X(_08140_));
 sky130_fd_sc_hd__o211a_2 _21280_ (.A1(_08131_),
    .A2(_08135_),
    .B1(_08138_),
    .C1(_08139_),
    .X(_08141_));
 sky130_fd_sc_hd__inv_2 _21281_ (.A(_08141_),
    .Y(_08142_));
 sky130_fd_sc_hd__a32o_2 _21282_ (.A1(_11712_),
    .A2(_08140_),
    .A3(_08142_),
    .B1(\systolic_inst.acc_wires[4][4] ),
    .B2(_11258_),
    .X(_01686_));
 sky130_fd_sc_hd__and2_2 _21283_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[4][5] ),
    .X(_08143_));
 sky130_fd_sc_hd__nand2_2 _21284_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[4][5] ),
    .Y(_08144_));
 sky130_fd_sc_hd__or2_2 _21285_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[4][5] ),
    .X(_08145_));
 sky130_fd_sc_hd__a211o_2 _21286_ (.A1(_08144_),
    .A2(_08145_),
    .B1(_08137_),
    .C1(_08141_),
    .X(_08146_));
 sky130_fd_sc_hd__o211a_2 _21287_ (.A1(_08137_),
    .A2(_08141_),
    .B1(_08144_),
    .C1(_08145_),
    .X(_08147_));
 sky130_fd_sc_hd__inv_2 _21288_ (.A(_08147_),
    .Y(_08148_));
 sky130_fd_sc_hd__a32o_2 _21289_ (.A1(_11712_),
    .A2(_08146_),
    .A3(_08148_),
    .B1(\systolic_inst.acc_wires[4][5] ),
    .B2(_11258_),
    .X(_01687_));
 sky130_fd_sc_hd__and2_2 _21290_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[4][6] ),
    .X(_08149_));
 sky130_fd_sc_hd__nand2_2 _21291_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[4][6] ),
    .Y(_08150_));
 sky130_fd_sc_hd__or2_2 _21292_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[4][6] ),
    .X(_08151_));
 sky130_fd_sc_hd__a211o_2 _21293_ (.A1(_08150_),
    .A2(_08151_),
    .B1(_08143_),
    .C1(_08147_),
    .X(_08152_));
 sky130_fd_sc_hd__o211a_2 _21294_ (.A1(_08143_),
    .A2(_08147_),
    .B1(_08150_),
    .C1(_08151_),
    .X(_08153_));
 sky130_fd_sc_hd__inv_2 _21295_ (.A(_08153_),
    .Y(_08154_));
 sky130_fd_sc_hd__a32o_2 _21296_ (.A1(_11712_),
    .A2(_08152_),
    .A3(_08154_),
    .B1(\systolic_inst.acc_wires[4][6] ),
    .B2(_11258_),
    .X(_01688_));
 sky130_fd_sc_hd__nand2_2 _21297_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[4][7] ),
    .Y(_08155_));
 sky130_fd_sc_hd__or2_2 _21298_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[4][7] ),
    .X(_08156_));
 sky130_fd_sc_hd__o211ai_2 _21299_ (.A1(_08149_),
    .A2(_08153_),
    .B1(_08155_),
    .C1(_08156_),
    .Y(_08157_));
 sky130_fd_sc_hd__a211o_2 _21300_ (.A1(_08155_),
    .A2(_08156_),
    .B1(_08149_),
    .C1(_08153_),
    .X(_08158_));
 sky130_fd_sc_hd__a32o_2 _21301_ (.A1(_11712_),
    .A2(_08157_),
    .A3(_08158_),
    .B1(\systolic_inst.acc_wires[4][7] ),
    .B2(_11258_),
    .X(_01689_));
 sky130_fd_sc_hd__or2_2 _21302_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[4][8] ),
    .X(_08159_));
 sky130_fd_sc_hd__nand2_2 _21303_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[4][8] ),
    .Y(_08160_));
 sky130_fd_sc_hd__nand2_2 _21304_ (.A(_08159_),
    .B(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__nand3_2 _21305_ (.A(_08155_),
    .B(_08157_),
    .C(_08161_),
    .Y(_08162_));
 sky130_fd_sc_hd__a21o_2 _21306_ (.A1(_08155_),
    .A2(_08157_),
    .B1(_08161_),
    .X(_08163_));
 sky130_fd_sc_hd__a32o_2 _21307_ (.A1(_11712_),
    .A2(_08162_),
    .A3(_08163_),
    .B1(\systolic_inst.acc_wires[4][8] ),
    .B2(_11258_),
    .X(_01690_));
 sky130_fd_sc_hd__nor2_2 _21308_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[4][9] ),
    .Y(_08164_));
 sky130_fd_sc_hd__nand2_2 _21309_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[4][9] ),
    .Y(_08165_));
 sky130_fd_sc_hd__and2b_2 _21310_ (.A_N(_08164_),
    .B(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__nand2_2 _21311_ (.A(_08160_),
    .B(_08163_),
    .Y(_08167_));
 sky130_fd_sc_hd__or2_2 _21312_ (.A(_08166_),
    .B(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__a21bo_2 _21313_ (.A1(_08160_),
    .A2(_08163_),
    .B1_N(_08166_),
    .X(_08169_));
 sky130_fd_sc_hd__a32o_2 _21314_ (.A1(_11712_),
    .A2(_08168_),
    .A3(_08169_),
    .B1(\systolic_inst.acc_wires[4][9] ),
    .B2(_11258_),
    .X(_01691_));
 sky130_fd_sc_hd__or2_2 _21315_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[4][10] ),
    .X(_08170_));
 sky130_fd_sc_hd__nand2_2 _21316_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[4][10] ),
    .Y(_08171_));
 sky130_fd_sc_hd__nand2_2 _21317_ (.A(_08170_),
    .B(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand3_2 _21318_ (.A(_08165_),
    .B(_08169_),
    .C(_08172_),
    .Y(_08173_));
 sky130_fd_sc_hd__a21o_2 _21319_ (.A1(_08165_),
    .A2(_08169_),
    .B1(_08172_),
    .X(_08174_));
 sky130_fd_sc_hd__a32o_2 _21320_ (.A1(_11712_),
    .A2(_08173_),
    .A3(_08174_),
    .B1(\systolic_inst.acc_wires[4][10] ),
    .B2(_11258_),
    .X(_01692_));
 sky130_fd_sc_hd__or2_2 _21321_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[4][11] ),
    .X(_08175_));
 sky130_fd_sc_hd__nand2_2 _21322_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[4][11] ),
    .Y(_08176_));
 sky130_fd_sc_hd__nand2_2 _21323_ (.A(_08175_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__nand3_2 _21324_ (.A(_08171_),
    .B(_08174_),
    .C(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__a21o_2 _21325_ (.A1(_08171_),
    .A2(_08174_),
    .B1(_08177_),
    .X(_08179_));
 sky130_fd_sc_hd__a32o_2 _21326_ (.A1(_11712_),
    .A2(_08178_),
    .A3(_08179_),
    .B1(\systolic_inst.acc_wires[4][11] ),
    .B2(_11258_),
    .X(_01693_));
 sky130_fd_sc_hd__nor2_2 _21327_ (.A(_08172_),
    .B(_08177_),
    .Y(_08180_));
 sky130_fd_sc_hd__nand2_2 _21328_ (.A(_08166_),
    .B(_08180_),
    .Y(_08181_));
 sky130_fd_sc_hd__a211o_2 _21329_ (.A1(_08155_),
    .A2(_08157_),
    .B1(_08161_),
    .C1(_08181_),
    .X(_08182_));
 sky130_fd_sc_hd__o21ai_2 _21330_ (.A1(_08160_),
    .A2(_08164_),
    .B1(_08165_),
    .Y(_08183_));
 sky130_fd_sc_hd__and3_2 _21331_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[4][10] ),
    .C(_08175_),
    .X(_08184_));
 sky130_fd_sc_hd__a221oi_2 _21332_ (.A1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[11] ),
    .A2(\systolic_inst.acc_wires[4][11] ),
    .B1(_08180_),
    .B2(_08183_),
    .C1(_08184_),
    .Y(_08185_));
 sky130_fd_sc_hd__and2_2 _21333_ (.A(_08182_),
    .B(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__or2_2 _21334_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[4][12] ),
    .X(_08187_));
 sky130_fd_sc_hd__nand2_2 _21335_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[4][12] ),
    .Y(_08188_));
 sky130_fd_sc_hd__nand2_2 _21336_ (.A(_08187_),
    .B(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__xor2_2 _21337_ (.A(_08186_),
    .B(_08189_),
    .X(_08190_));
 sky130_fd_sc_hd__a22o_2 _21338_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[4][12] ),
    .B1(_11712_),
    .B2(_08190_),
    .X(_01694_));
 sky130_fd_sc_hd__or2_2 _21339_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[4][13] ),
    .X(_08191_));
 sky130_fd_sc_hd__nand2_2 _21340_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[4][13] ),
    .Y(_08192_));
 sky130_fd_sc_hd__nand2_2 _21341_ (.A(_08191_),
    .B(_08192_),
    .Y(_08193_));
 sky130_fd_sc_hd__o211a_2 _21342_ (.A1(_08186_),
    .A2(_08189_),
    .B1(_08193_),
    .C1(_08188_),
    .X(_08194_));
 sky130_fd_sc_hd__a211o_2 _21343_ (.A1(_08182_),
    .A2(_08185_),
    .B1(_08189_),
    .C1(_08193_),
    .X(_08195_));
 sky130_fd_sc_hd__o211ai_2 _21344_ (.A1(_08188_),
    .A2(_08193_),
    .B1(_08195_),
    .C1(_11712_),
    .Y(_08196_));
 sky130_fd_sc_hd__a2bb2o_2 _21345_ (.A1_N(_08196_),
    .A2_N(_08194_),
    .B1(\systolic_inst.acc_wires[4][13] ),
    .B2(_11258_),
    .X(_01695_));
 sky130_fd_sc_hd__or2_2 _21346_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[4][14] ),
    .X(_08197_));
 sky130_fd_sc_hd__nand2_2 _21347_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[4][14] ),
    .Y(_08198_));
 sky130_fd_sc_hd__and2_2 _21348_ (.A(_08197_),
    .B(_08198_),
    .X(_08199_));
 sky130_fd_sc_hd__o21a_2 _21349_ (.A1(_08188_),
    .A2(_08193_),
    .B1(_08192_),
    .X(_08200_));
 sky130_fd_sc_hd__nand2_2 _21350_ (.A(_08195_),
    .B(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__nand2_2 _21351_ (.A(_08199_),
    .B(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__or2_2 _21352_ (.A(_08199_),
    .B(_08201_),
    .X(_08203_));
 sky130_fd_sc_hd__a32o_2 _21353_ (.A1(_11712_),
    .A2(_08202_),
    .A3(_08203_),
    .B1(\systolic_inst.acc_wires[4][14] ),
    .B2(_11258_),
    .X(_01696_));
 sky130_fd_sc_hd__nor2_2 _21354_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][15] ),
    .Y(_08204_));
 sky130_fd_sc_hd__and2_2 _21355_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][15] ),
    .X(_08205_));
 sky130_fd_sc_hd__a211o_2 _21356_ (.A1(_08198_),
    .A2(_08202_),
    .B1(_08204_),
    .C1(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__o211ai_2 _21357_ (.A1(_08204_),
    .A2(_08205_),
    .B1(_08198_),
    .C1(_08202_),
    .Y(_08207_));
 sky130_fd_sc_hd__a32o_2 _21358_ (.A1(_11712_),
    .A2(_08206_),
    .A3(_08207_),
    .B1(\systolic_inst.acc_wires[4][15] ),
    .B2(_11258_),
    .X(_01697_));
 sky130_fd_sc_hd__or3b_2 _21359_ (.A(_08204_),
    .B(_08205_),
    .C_N(_08199_),
    .X(_08208_));
 sky130_fd_sc_hd__a21o_2 _21360_ (.A1(_08195_),
    .A2(_08200_),
    .B1(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__o21ba_2 _21361_ (.A1(_08198_),
    .A2(_08204_),
    .B1_N(_08205_),
    .X(_08210_));
 sky130_fd_sc_hd__and2_2 _21362_ (.A(_08209_),
    .B(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__or2_2 _21363_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][16] ),
    .X(_08212_));
 sky130_fd_sc_hd__nand2_2 _21364_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][16] ),
    .Y(_08213_));
 sky130_fd_sc_hd__nand2_2 _21365_ (.A(_08212_),
    .B(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__nand2_2 _21366_ (.A(_08211_),
    .B(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__nor2_2 _21367_ (.A(_08211_),
    .B(_08214_),
    .Y(_08216_));
 sky130_fd_sc_hd__nor2_2 _21368_ (.A(_11713_),
    .B(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__a22o_2 _21369_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[4][16] ),
    .B1(_08215_),
    .B2(_08217_),
    .X(_01698_));
 sky130_fd_sc_hd__xor2_2 _21370_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][17] ),
    .X(_08218_));
 sky130_fd_sc_hd__o21a_2 _21371_ (.A1(_08211_),
    .A2(_08214_),
    .B1(_08213_),
    .X(_08219_));
 sky130_fd_sc_hd__xnor2_2 _21372_ (.A(_08218_),
    .B(_08219_),
    .Y(_08220_));
 sky130_fd_sc_hd__a22o_2 _21373_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[4][17] ),
    .B1(_11712_),
    .B2(_08220_),
    .X(_01699_));
 sky130_fd_sc_hd__or2_2 _21374_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][18] ),
    .X(_08221_));
 sky130_fd_sc_hd__nand2_2 _21375_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][18] ),
    .Y(_08222_));
 sky130_fd_sc_hd__nand2_2 _21376_ (.A(_08221_),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__o21ai_2 _21377_ (.A1(\systolic_inst.acc_wires[4][16] ),
    .A2(\systolic_inst.acc_wires[4][17] ),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .Y(_08224_));
 sky130_fd_sc_hd__nand2_2 _21378_ (.A(_08216_),
    .B(_08218_),
    .Y(_08225_));
 sky130_fd_sc_hd__a21o_2 _21379_ (.A1(_08224_),
    .A2(_08225_),
    .B1(_08223_),
    .X(_08226_));
 sky130_fd_sc_hd__nand3_2 _21380_ (.A(_08223_),
    .B(_08224_),
    .C(_08225_),
    .Y(_08227_));
 sky130_fd_sc_hd__a32o_2 _21381_ (.A1(_11712_),
    .A2(_08226_),
    .A3(_08227_),
    .B1(\systolic_inst.acc_wires[4][18] ),
    .B2(_11258_),
    .X(_01700_));
 sky130_fd_sc_hd__xnor2_2 _21382_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][19] ),
    .Y(_08228_));
 sky130_fd_sc_hd__a21oi_2 _21383_ (.A1(_08222_),
    .A2(_08226_),
    .B1(_08228_),
    .Y(_08229_));
 sky130_fd_sc_hd__a31o_2 _21384_ (.A1(_08222_),
    .A2(_08226_),
    .A3(_08228_),
    .B1(_11713_),
    .X(_08230_));
 sky130_fd_sc_hd__a2bb2o_2 _21385_ (.A1_N(_08230_),
    .A2_N(_08229_),
    .B1(\systolic_inst.acc_wires[4][19] ),
    .B2(_11258_),
    .X(_01701_));
 sky130_fd_sc_hd__or2_2 _21386_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][20] ),
    .X(_08231_));
 sky130_fd_sc_hd__nand2_2 _21387_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][20] ),
    .Y(_08232_));
 sky130_fd_sc_hd__and2_2 _21388_ (.A(_08231_),
    .B(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__and3_2 _21389_ (.A(_08212_),
    .B(_08213_),
    .C(_08218_),
    .X(_08234_));
 sky130_fd_sc_hd__or3b_2 _21390_ (.A(_08223_),
    .B(_08228_),
    .C_N(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__nor2_2 _21391_ (.A(_08211_),
    .B(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__o41a_2 _21392_ (.A1(\systolic_inst.acc_wires[4][16] ),
    .A2(\systolic_inst.acc_wires[4][17] ),
    .A3(\systolic_inst.acc_wires[4][18] ),
    .A4(\systolic_inst.acc_wires[4][19] ),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .X(_08237_));
 sky130_fd_sc_hd__or3_2 _21393_ (.A(_08233_),
    .B(_08236_),
    .C(_08237_),
    .X(_08238_));
 sky130_fd_sc_hd__o21ai_2 _21394_ (.A1(_08236_),
    .A2(_08237_),
    .B1(_08233_),
    .Y(_08239_));
 sky130_fd_sc_hd__a32o_2 _21395_ (.A1(_11712_),
    .A2(_08238_),
    .A3(_08239_),
    .B1(\systolic_inst.acc_wires[4][20] ),
    .B2(_11258_),
    .X(_01702_));
 sky130_fd_sc_hd__xnor2_2 _21396_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][21] ),
    .Y(_08240_));
 sky130_fd_sc_hd__inv_2 _21397_ (.A(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__a21oi_2 _21398_ (.A1(_08232_),
    .A2(_08239_),
    .B1(_08240_),
    .Y(_08242_));
 sky130_fd_sc_hd__a31o_2 _21399_ (.A1(_08232_),
    .A2(_08239_),
    .A3(_08240_),
    .B1(_11713_),
    .X(_08243_));
 sky130_fd_sc_hd__a2bb2o_2 _21400_ (.A1_N(_08243_),
    .A2_N(_08242_),
    .B1(\systolic_inst.acc_wires[4][21] ),
    .B2(_11258_),
    .X(_01703_));
 sky130_fd_sc_hd__or2_2 _21401_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][22] ),
    .X(_08244_));
 sky130_fd_sc_hd__nand2_2 _21402_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][22] ),
    .Y(_08245_));
 sky130_fd_sc_hd__and2_2 _21403_ (.A(_08244_),
    .B(_08245_),
    .X(_08246_));
 sky130_fd_sc_hd__o21a_2 _21404_ (.A1(\systolic_inst.acc_wires[4][20] ),
    .A2(\systolic_inst.acc_wires[4][21] ),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .X(_08247_));
 sky130_fd_sc_hd__nor2_2 _21405_ (.A(_08239_),
    .B(_08240_),
    .Y(_08248_));
 sky130_fd_sc_hd__o21ai_2 _21406_ (.A1(_08247_),
    .A2(_08248_),
    .B1(_08246_),
    .Y(_08249_));
 sky130_fd_sc_hd__or3_2 _21407_ (.A(_08246_),
    .B(_08247_),
    .C(_08248_),
    .X(_08250_));
 sky130_fd_sc_hd__a32o_2 _21408_ (.A1(_11712_),
    .A2(_08249_),
    .A3(_08250_),
    .B1(\systolic_inst.acc_wires[4][22] ),
    .B2(_11258_),
    .X(_01704_));
 sky130_fd_sc_hd__xor2_2 _21409_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][23] ),
    .X(_08251_));
 sky130_fd_sc_hd__inv_2 _21410_ (.A(_08251_),
    .Y(_08252_));
 sky130_fd_sc_hd__nand3_2 _21411_ (.A(_08245_),
    .B(_08249_),
    .C(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__a21o_2 _21412_ (.A1(_08245_),
    .A2(_08249_),
    .B1(_08252_),
    .X(_08254_));
 sky130_fd_sc_hd__a32o_2 _21413_ (.A1(_11712_),
    .A2(_08253_),
    .A3(_08254_),
    .B1(\systolic_inst.acc_wires[4][23] ),
    .B2(_11258_),
    .X(_01705_));
 sky130_fd_sc_hd__nand4_2 _21414_ (.A(_08233_),
    .B(_08241_),
    .C(_08246_),
    .D(_08251_),
    .Y(_08255_));
 sky130_fd_sc_hd__a211o_2 _21415_ (.A1(_08209_),
    .A2(_08210_),
    .B1(_08235_),
    .C1(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__o41a_2 _21416_ (.A1(\systolic_inst.acc_wires[4][20] ),
    .A2(\systolic_inst.acc_wires[4][21] ),
    .A3(\systolic_inst.acc_wires[4][22] ),
    .A4(\systolic_inst.acc_wires[4][23] ),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .X(_08257_));
 sky130_fd_sc_hd__nor2_2 _21417_ (.A(_08237_),
    .B(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__nor2_2 _21418_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][24] ),
    .Y(_08259_));
 sky130_fd_sc_hd__and2_2 _21419_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][24] ),
    .X(_08260_));
 sky130_fd_sc_hd__or2_2 _21420_ (.A(_08259_),
    .B(_08260_),
    .X(_08261_));
 sky130_fd_sc_hd__a21oi_2 _21421_ (.A1(_08256_),
    .A2(_08258_),
    .B1(_08261_),
    .Y(_08262_));
 sky130_fd_sc_hd__a31o_2 _21422_ (.A1(_08256_),
    .A2(_08258_),
    .A3(_08261_),
    .B1(_11713_),
    .X(_08263_));
 sky130_fd_sc_hd__a2bb2o_2 _21423_ (.A1_N(_08263_),
    .A2_N(_08262_),
    .B1(\systolic_inst.acc_wires[4][24] ),
    .B2(_11258_),
    .X(_01706_));
 sky130_fd_sc_hd__xor2_2 _21424_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][25] ),
    .X(_08264_));
 sky130_fd_sc_hd__or3_2 _21425_ (.A(_08260_),
    .B(_08262_),
    .C(_08264_),
    .X(_08265_));
 sky130_fd_sc_hd__o21ai_2 _21426_ (.A1(_08260_),
    .A2(_08262_),
    .B1(_08264_),
    .Y(_08266_));
 sky130_fd_sc_hd__a32o_2 _21427_ (.A1(_11712_),
    .A2(_08265_),
    .A3(_08266_),
    .B1(\systolic_inst.acc_wires[4][25] ),
    .B2(_11258_),
    .X(_01707_));
 sky130_fd_sc_hd__or2_2 _21428_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][26] ),
    .X(_08267_));
 sky130_fd_sc_hd__nand2_2 _21429_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][26] ),
    .Y(_08268_));
 sky130_fd_sc_hd__nand2_2 _21430_ (.A(_08267_),
    .B(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__o21a_2 _21431_ (.A1(\systolic_inst.acc_wires[4][24] ),
    .A2(\systolic_inst.acc_wires[4][25] ),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .X(_08270_));
 sky130_fd_sc_hd__a21o_2 _21432_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08270_),
    .X(_08271_));
 sky130_fd_sc_hd__xnor2_2 _21433_ (.A(_08269_),
    .B(_08271_),
    .Y(_08272_));
 sky130_fd_sc_hd__a22o_2 _21434_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[4][26] ),
    .B1(_11712_),
    .B2(_08272_),
    .X(_01708_));
 sky130_fd_sc_hd__xnor2_2 _21435_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][27] ),
    .Y(_08273_));
 sky130_fd_sc_hd__a21bo_2 _21436_ (.A1(_08267_),
    .A2(_08271_),
    .B1_N(_08268_),
    .X(_08274_));
 sky130_fd_sc_hd__xnor2_2 _21437_ (.A(_08273_),
    .B(_08274_),
    .Y(_08275_));
 sky130_fd_sc_hd__a22o_2 _21438_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[4][27] ),
    .B1(_11712_),
    .B2(_08275_),
    .X(_01709_));
 sky130_fd_sc_hd__nor2_2 _21439_ (.A(_08269_),
    .B(_08273_),
    .Y(_08276_));
 sky130_fd_sc_hd__o21a_2 _21440_ (.A1(\systolic_inst.acc_wires[4][26] ),
    .A2(\systolic_inst.acc_wires[4][27] ),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .X(_08277_));
 sky130_fd_sc_hd__a311oi_2 _21441_ (.A1(_08262_),
    .A2(_08264_),
    .A3(_08276_),
    .B1(_08277_),
    .C1(_08270_),
    .Y(_08278_));
 sky130_fd_sc_hd__or2_2 _21442_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][28] ),
    .X(_08279_));
 sky130_fd_sc_hd__nand2_2 _21443_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][28] ),
    .Y(_08280_));
 sky130_fd_sc_hd__nand2_2 _21444_ (.A(_08279_),
    .B(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__xor2_2 _21445_ (.A(_08278_),
    .B(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__a22o_2 _21446_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[4][28] ),
    .B1(_11712_),
    .B2(_08282_),
    .X(_01710_));
 sky130_fd_sc_hd__xor2_2 _21447_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][29] ),
    .X(_08283_));
 sky130_fd_sc_hd__inv_2 _21448_ (.A(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__o21a_2 _21449_ (.A1(_08278_),
    .A2(_08281_),
    .B1(_08280_),
    .X(_08285_));
 sky130_fd_sc_hd__xnor2_2 _21450_ (.A(_08283_),
    .B(_08285_),
    .Y(_08286_));
 sky130_fd_sc_hd__a22o_2 _21451_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[4][29] ),
    .B1(_11712_),
    .B2(_08286_),
    .X(_01711_));
 sky130_fd_sc_hd__o21ai_2 _21452_ (.A1(\systolic_inst.acc_wires[4][28] ),
    .A2(\systolic_inst.acc_wires[4][29] ),
    .B1(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .Y(_08287_));
 sky130_fd_sc_hd__o31a_2 _21453_ (.A1(_08278_),
    .A2(_08281_),
    .A3(_08284_),
    .B1(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__nand2_2 _21454_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][30] ),
    .Y(_08289_));
 sky130_fd_sc_hd__or2_2 _21455_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][30] ),
    .X(_08290_));
 sky130_fd_sc_hd__nand2_2 _21456_ (.A(_08289_),
    .B(_08290_),
    .Y(_08291_));
 sky130_fd_sc_hd__nand2_2 _21457_ (.A(_08288_),
    .B(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__or2_2 _21458_ (.A(_08288_),
    .B(_08291_),
    .X(_08293_));
 sky130_fd_sc_hd__a32o_2 _21459_ (.A1(_11712_),
    .A2(_08292_),
    .A3(_08293_),
    .B1(\systolic_inst.acc_wires[4][30] ),
    .B2(_11258_),
    .X(_01712_));
 sky130_fd_sc_hd__xnor2_2 _21460_ (.A(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[4][31] ),
    .Y(_08294_));
 sky130_fd_sc_hd__a21oi_2 _21461_ (.A1(_08289_),
    .A2(_08293_),
    .B1(_08294_),
    .Y(_08295_));
 sky130_fd_sc_hd__a31o_2 _21462_ (.A1(_08289_),
    .A2(_08293_),
    .A3(_08294_),
    .B1(_11713_),
    .X(_08296_));
 sky130_fd_sc_hd__a2bb2o_2 _21463_ (.A1_N(_08296_),
    .A2_N(_08295_),
    .B1(\systolic_inst.acc_wires[4][31] ),
    .B2(_11258_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _21464_ (.A0(\systolic_inst.A_outs[3][0] ),
    .A1(\systolic_inst.A_outs[2][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _21465_ (.A0(\systolic_inst.A_outs[3][1] ),
    .A1(\systolic_inst.A_outs[2][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _21466_ (.A0(\systolic_inst.A_outs[3][2] ),
    .A1(\systolic_inst.A_outs[2][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _21467_ (.A0(\systolic_inst.A_outs[3][3] ),
    .A1(\systolic_inst.A_outs[2][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _21468_ (.A0(\systolic_inst.A_outs[3][4] ),
    .A1(\systolic_inst.A_outs[2][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _21469_ (.A0(\systolic_inst.A_outs[3][5] ),
    .A1(\systolic_inst.A_outs[2][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _21470_ (.A0(\systolic_inst.A_outs[3][6] ),
    .A1(\systolic_inst.A_outs[2][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _21471_ (.A0(\systolic_inst.A_outs[3][7] ),
    .A1(\systolic_inst.A_outs[2][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _21472_ (.A0(\systolic_inst.B_outs[2][0] ),
    .A1(\systolic_inst.B_shift[2][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _21473_ (.A0(\systolic_inst.B_outs[2][1] ),
    .A1(\systolic_inst.B_shift[2][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _21474_ (.A0(\systolic_inst.B_outs[2][2] ),
    .A1(\systolic_inst.B_shift[2][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _21475_ (.A0(\systolic_inst.B_outs[2][3] ),
    .A1(\systolic_inst.B_shift[2][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _21476_ (.A0(\systolic_inst.B_outs[2][4] ),
    .A1(\systolic_inst.B_shift[2][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _21477_ (.A0(\systolic_inst.B_outs[2][5] ),
    .A1(\systolic_inst.B_shift[2][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _21478_ (.A0(\systolic_inst.B_outs[2][6] ),
    .A1(\systolic_inst.B_shift[2][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _21479_ (.A0(\systolic_inst.B_outs[2][7] ),
    .A1(\systolic_inst.B_shift[2][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01729_));
 sky130_fd_sc_hd__and3_2 _21480_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[3][0] ),
    .C(\systolic_inst.A_outs[3][0] ),
    .X(_08297_));
 sky130_fd_sc_hd__a21o_2 _21481_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[0] ),
    .B1(_08297_),
    .X(_01730_));
 sky130_fd_sc_hd__and4_2 _21482_ (.A(\systolic_inst.B_outs[3][0] ),
    .B(\systolic_inst.A_outs[3][0] ),
    .C(\systolic_inst.B_outs[3][1] ),
    .D(\systolic_inst.A_outs[3][1] ),
    .X(_08298_));
 sky130_fd_sc_hd__inv_2 _21483_ (.A(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__a22o_2 _21484_ (.A1(\systolic_inst.A_outs[3][0] ),
    .A2(\systolic_inst.B_outs[3][1] ),
    .B1(\systolic_inst.A_outs[3][1] ),
    .B2(\systolic_inst.B_outs[3][0] ),
    .X(_08300_));
 sky130_fd_sc_hd__and2_2 _21485_ (.A(\systolic_inst.ce_local ),
    .B(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__a22o_2 _21486_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[1] ),
    .B1(_08299_),
    .B2(_08301_),
    .X(_01731_));
 sky130_fd_sc_hd__nand2_2 _21487_ (.A(\systolic_inst.B_outs[3][1] ),
    .B(\systolic_inst.A_outs[3][1] ),
    .Y(_08302_));
 sky130_fd_sc_hd__nand2_2 _21488_ (.A(\systolic_inst.B_outs[3][0] ),
    .B(\systolic_inst.A_outs[3][2] ),
    .Y(_08303_));
 sky130_fd_sc_hd__and4_2 _21489_ (.A(\systolic_inst.B_outs[3][0] ),
    .B(\systolic_inst.B_outs[3][1] ),
    .C(\systolic_inst.A_outs[3][1] ),
    .D(\systolic_inst.A_outs[3][2] ),
    .X(_08304_));
 sky130_fd_sc_hd__a21o_2 _21490_ (.A1(_08302_),
    .A2(_08303_),
    .B1(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__xnor2_2 _21491_ (.A(_08298_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__and2_2 _21492_ (.A(\systolic_inst.A_outs[3][0] ),
    .B(\systolic_inst.B_outs[3][2] ),
    .X(_08307_));
 sky130_fd_sc_hd__nand2_2 _21493_ (.A(_08306_),
    .B(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__o21a_2 _21494_ (.A1(_08306_),
    .A2(_08307_),
    .B1(\systolic_inst.ce_local ),
    .X(_08309_));
 sky130_fd_sc_hd__a22o_2 _21495_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[2] ),
    .B1(_08308_),
    .B2(_08309_),
    .X(_01732_));
 sky130_fd_sc_hd__a22oi_2 _21496_ (.A1(\systolic_inst.A_outs[3][1] ),
    .A2(\systolic_inst.B_outs[3][2] ),
    .B1(\systolic_inst.B_outs[3][3] ),
    .B2(\systolic_inst.A_outs[3][0] ),
    .Y(_08310_));
 sky130_fd_sc_hd__and4_2 _21497_ (.A(\systolic_inst.A_outs[3][0] ),
    .B(\systolic_inst.A_outs[3][1] ),
    .C(\systolic_inst.B_outs[3][2] ),
    .D(\systolic_inst.B_outs[3][3] ),
    .X(_08311_));
 sky130_fd_sc_hd__or2_2 _21498_ (.A(_08310_),
    .B(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__nand2_2 _21499_ (.A(\systolic_inst.B_outs[3][1] ),
    .B(\systolic_inst.A_outs[3][3] ),
    .Y(_08313_));
 sky130_fd_sc_hd__or2_2 _21500_ (.A(_08303_),
    .B(_08313_),
    .X(_08314_));
 sky130_fd_sc_hd__a22o_2 _21501_ (.A1(\systolic_inst.B_outs[3][1] ),
    .A2(\systolic_inst.A_outs[3][2] ),
    .B1(\systolic_inst.A_outs[3][3] ),
    .B2(\systolic_inst.B_outs[3][0] ),
    .X(_08315_));
 sky130_fd_sc_hd__nand3_2 _21502_ (.A(_08304_),
    .B(_08314_),
    .C(_08315_),
    .Y(_08316_));
 sky130_fd_sc_hd__a21o_2 _21503_ (.A1(_08314_),
    .A2(_08315_),
    .B1(_08304_),
    .X(_08317_));
 sky130_fd_sc_hd__nand2_2 _21504_ (.A(_08316_),
    .B(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__or2_2 _21505_ (.A(_08312_),
    .B(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__xnor2_2 _21506_ (.A(_08312_),
    .B(_08318_),
    .Y(_08320_));
 sky130_fd_sc_hd__o21ai_2 _21507_ (.A1(_08299_),
    .A2(_08305_),
    .B1(_08308_),
    .Y(_08321_));
 sky130_fd_sc_hd__and2b_2 _21508_ (.A_N(_08320_),
    .B(_08321_),
    .X(_08322_));
 sky130_fd_sc_hd__xnor2_2 _21509_ (.A(_08320_),
    .B(_08321_),
    .Y(_08323_));
 sky130_fd_sc_hd__mux2_1 _21510_ (.A0(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[3] ),
    .A1(_08323_),
    .S(\systolic_inst.ce_local ),
    .X(_01733_));
 sky130_fd_sc_hd__and2_2 _21511_ (.A(\systolic_inst.B_outs[3][2] ),
    .B(\systolic_inst.A_outs[3][2] ),
    .X(_08324_));
 sky130_fd_sc_hd__nand4_2 _21512_ (.A(\systolic_inst.A_outs[3][0] ),
    .B(\systolic_inst.A_outs[3][1] ),
    .C(\systolic_inst.B_outs[3][3] ),
    .D(\systolic_inst.B_outs[3][4] ),
    .Y(_08325_));
 sky130_fd_sc_hd__a22o_2 _21513_ (.A1(\systolic_inst.A_outs[3][1] ),
    .A2(\systolic_inst.B_outs[3][3] ),
    .B1(\systolic_inst.B_outs[3][4] ),
    .B2(\systolic_inst.A_outs[3][0] ),
    .X(_08326_));
 sky130_fd_sc_hd__nand2_2 _21514_ (.A(_08325_),
    .B(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__xnor2_2 _21515_ (.A(_08324_),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__inv_2 _21516_ (.A(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__nand2_2 _21517_ (.A(\systolic_inst.B_outs[3][0] ),
    .B(\systolic_inst.A_outs[3][4] ),
    .Y(_08330_));
 sky130_fd_sc_hd__and4_2 _21518_ (.A(\systolic_inst.B_outs[3][0] ),
    .B(\systolic_inst.B_outs[3][1] ),
    .C(\systolic_inst.A_outs[3][3] ),
    .D(\systolic_inst.A_outs[3][4] ),
    .X(_08331_));
 sky130_fd_sc_hd__a21oi_2 _21519_ (.A1(_08313_),
    .A2(_08330_),
    .B1(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__xnor2_2 _21520_ (.A(_08311_),
    .B(_08332_),
    .Y(_08333_));
 sky130_fd_sc_hd__nor2_2 _21521_ (.A(_08314_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__xnor2_2 _21522_ (.A(_08314_),
    .B(_08333_),
    .Y(_08335_));
 sky130_fd_sc_hd__nor2_2 _21523_ (.A(_08329_),
    .B(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__xnor2_2 _21524_ (.A(_08329_),
    .B(_08335_),
    .Y(_08337_));
 sky130_fd_sc_hd__a21o_2 _21525_ (.A1(_08316_),
    .A2(_08319_),
    .B1(_08337_),
    .X(_08338_));
 sky130_fd_sc_hd__inv_2 _21526_ (.A(_08338_),
    .Y(_08339_));
 sky130_fd_sc_hd__nand3_2 _21527_ (.A(_08316_),
    .B(_08319_),
    .C(_08337_),
    .Y(_08340_));
 sky130_fd_sc_hd__a21oi_2 _21528_ (.A1(_08338_),
    .A2(_08340_),
    .B1(_08322_),
    .Y(_08341_));
 sky130_fd_sc_hd__and3_2 _21529_ (.A(_08322_),
    .B(_08338_),
    .C(_08340_),
    .X(_08342_));
 sky130_fd_sc_hd__or3_2 _21530_ (.A(_11258_),
    .B(_08341_),
    .C(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__a21bo_2 _21531_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[4] ),
    .B1_N(_08343_),
    .X(_01734_));
 sky130_fd_sc_hd__and2_2 _21532_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[5] ),
    .X(_08344_));
 sky130_fd_sc_hd__a21oi_2 _21533_ (.A1(_08311_),
    .A2(_08332_),
    .B1(_08334_),
    .Y(_08345_));
 sky130_fd_sc_hd__a21bo_2 _21534_ (.A1(_08324_),
    .A2(_08326_),
    .B1_N(_08325_),
    .X(_08346_));
 sky130_fd_sc_hd__a22oi_2 _21535_ (.A1(\systolic_inst.B_outs[3][1] ),
    .A2(\systolic_inst.A_outs[3][4] ),
    .B1(\systolic_inst.A_outs[3][5] ),
    .B2(\systolic_inst.B_outs[3][0] ),
    .Y(_08347_));
 sky130_fd_sc_hd__and4_2 _21536_ (.A(\systolic_inst.B_outs[3][0] ),
    .B(\systolic_inst.B_outs[3][1] ),
    .C(\systolic_inst.A_outs[3][4] ),
    .D(\systolic_inst.A_outs[3][5] ),
    .X(_08348_));
 sky130_fd_sc_hd__or2_2 _21537_ (.A(_08347_),
    .B(_08348_),
    .X(_08349_));
 sky130_fd_sc_hd__nand2b_2 _21538_ (.A_N(_08349_),
    .B(_08346_),
    .Y(_08350_));
 sky130_fd_sc_hd__xnor2_2 _21539_ (.A(_08346_),
    .B(_08349_),
    .Y(_08351_));
 sky130_fd_sc_hd__nand2_2 _21540_ (.A(_08331_),
    .B(_08351_),
    .Y(_08352_));
 sky130_fd_sc_hd__xnor2_2 _21541_ (.A(_08331_),
    .B(_08351_),
    .Y(_08353_));
 sky130_fd_sc_hd__nand2_2 _21542_ (.A(\systolic_inst.A_outs[3][0] ),
    .B(\systolic_inst.B_outs[3][5] ),
    .Y(_08354_));
 sky130_fd_sc_hd__nand2_2 _21543_ (.A(\systolic_inst.B_outs[3][2] ),
    .B(\systolic_inst.A_outs[3][3] ),
    .Y(_08355_));
 sky130_fd_sc_hd__and4_2 _21544_ (.A(\systolic_inst.A_outs[3][1] ),
    .B(\systolic_inst.A_outs[3][2] ),
    .C(\systolic_inst.B_outs[3][3] ),
    .D(\systolic_inst.B_outs[3][4] ),
    .X(_08356_));
 sky130_fd_sc_hd__a22o_2 _21545_ (.A1(\systolic_inst.A_outs[3][2] ),
    .A2(\systolic_inst.B_outs[3][3] ),
    .B1(\systolic_inst.B_outs[3][4] ),
    .B2(\systolic_inst.A_outs[3][1] ),
    .X(_08357_));
 sky130_fd_sc_hd__and2b_2 _21546_ (.A_N(_08356_),
    .B(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__xnor2_2 _21547_ (.A(_08355_),
    .B(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__nand2b_2 _21548_ (.A_N(_08354_),
    .B(_08359_),
    .Y(_08360_));
 sky130_fd_sc_hd__xor2_2 _21549_ (.A(_08354_),
    .B(_08359_),
    .X(_08361_));
 sky130_fd_sc_hd__nor2_2 _21550_ (.A(_08353_),
    .B(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__inv_2 _21551_ (.A(_08362_),
    .Y(_08363_));
 sky130_fd_sc_hd__xor2_2 _21552_ (.A(_08353_),
    .B(_08361_),
    .X(_08364_));
 sky130_fd_sc_hd__nand2_2 _21553_ (.A(_08336_),
    .B(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__or2_2 _21554_ (.A(_08336_),
    .B(_08364_),
    .X(_08366_));
 sky130_fd_sc_hd__and2_2 _21555_ (.A(_08365_),
    .B(_08366_),
    .X(_08367_));
 sky130_fd_sc_hd__nand2b_2 _21556_ (.A_N(_08345_),
    .B(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__xnor2_2 _21557_ (.A(_08345_),
    .B(_08367_),
    .Y(_08369_));
 sky130_fd_sc_hd__nor2_2 _21558_ (.A(_08339_),
    .B(_08342_),
    .Y(_08370_));
 sky130_fd_sc_hd__or3_2 _21559_ (.A(_08339_),
    .B(_08342_),
    .C(_08369_),
    .X(_08371_));
 sky130_fd_sc_hd__nand2b_2 _21560_ (.A_N(_08370_),
    .B(_08369_),
    .Y(_08372_));
 sky130_fd_sc_hd__a31o_2 _21561_ (.A1(\systolic_inst.ce_local ),
    .A2(_08371_),
    .A3(_08372_),
    .B1(_08344_),
    .X(_01735_));
 sky130_fd_sc_hd__a31o_2 _21562_ (.A1(\systolic_inst.B_outs[3][2] ),
    .A2(\systolic_inst.A_outs[3][3] ),
    .A3(_08357_),
    .B1(_08356_),
    .X(_08373_));
 sky130_fd_sc_hd__a22oi_2 _21563_ (.A1(\systolic_inst.B_outs[3][1] ),
    .A2(\systolic_inst.A_outs[3][5] ),
    .B1(\systolic_inst.A_outs[3][6] ),
    .B2(\systolic_inst.B_outs[3][0] ),
    .Y(_08374_));
 sky130_fd_sc_hd__and4_2 _21564_ (.A(\systolic_inst.B_outs[3][0] ),
    .B(\systolic_inst.B_outs[3][1] ),
    .C(\systolic_inst.A_outs[3][5] ),
    .D(\systolic_inst.A_outs[3][6] ),
    .X(_08375_));
 sky130_fd_sc_hd__nor2_2 _21565_ (.A(_08374_),
    .B(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__xor2_2 _21566_ (.A(_08373_),
    .B(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__and2_2 _21567_ (.A(_08348_),
    .B(_08377_),
    .X(_08378_));
 sky130_fd_sc_hd__nor2_2 _21568_ (.A(_08348_),
    .B(_08377_),
    .Y(_08379_));
 sky130_fd_sc_hd__or2_2 _21569_ (.A(_08378_),
    .B(_08379_),
    .X(_08380_));
 sky130_fd_sc_hd__nand2_2 _21570_ (.A(\systolic_inst.B_outs[3][2] ),
    .B(\systolic_inst.A_outs[3][4] ),
    .Y(_08381_));
 sky130_fd_sc_hd__and4_2 _21571_ (.A(\systolic_inst.A_outs[3][2] ),
    .B(\systolic_inst.B_outs[3][3] ),
    .C(\systolic_inst.A_outs[3][3] ),
    .D(\systolic_inst.B_outs[3][4] ),
    .X(_08382_));
 sky130_fd_sc_hd__a22oi_2 _21572_ (.A1(\systolic_inst.B_outs[3][3] ),
    .A2(\systolic_inst.A_outs[3][3] ),
    .B1(\systolic_inst.B_outs[3][4] ),
    .B2(\systolic_inst.A_outs[3][2] ),
    .Y(_08383_));
 sky130_fd_sc_hd__or2_2 _21573_ (.A(_08382_),
    .B(_08383_),
    .X(_08384_));
 sky130_fd_sc_hd__xnor2_2 _21574_ (.A(_08381_),
    .B(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__a22oi_2 _21575_ (.A1(\systolic_inst.A_outs[3][1] ),
    .A2(\systolic_inst.B_outs[3][5] ),
    .B1(\systolic_inst.B_outs[3][6] ),
    .B2(\systolic_inst.A_outs[3][0] ),
    .Y(_08386_));
 sky130_fd_sc_hd__nand2_2 _21576_ (.A(\systolic_inst.A_outs[3][1] ),
    .B(\systolic_inst.B_outs[3][6] ),
    .Y(_08387_));
 sky130_fd_sc_hd__nor2_2 _21577_ (.A(_08354_),
    .B(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__nor2_2 _21578_ (.A(_08386_),
    .B(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__or3_2 _21579_ (.A(_08385_),
    .B(_08386_),
    .C(_08388_),
    .X(_08390_));
 sky130_fd_sc_hd__xor2_2 _21580_ (.A(_08385_),
    .B(_08389_),
    .X(_08391_));
 sky130_fd_sc_hd__xnor2_2 _21581_ (.A(_08360_),
    .B(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__xnor2_2 _21582_ (.A(_08380_),
    .B(_08392_),
    .Y(_08393_));
 sky130_fd_sc_hd__xnor2_2 _21583_ (.A(_08363_),
    .B(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__a21oi_2 _21584_ (.A1(_08350_),
    .A2(_08352_),
    .B1(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__and3_2 _21585_ (.A(_08350_),
    .B(_08352_),
    .C(_08394_),
    .X(_08396_));
 sky130_fd_sc_hd__a211oi_2 _21586_ (.A1(_08365_),
    .A2(_08368_),
    .B1(_08395_),
    .C1(_08396_),
    .Y(_08397_));
 sky130_fd_sc_hd__o211a_2 _21587_ (.A1(_08395_),
    .A2(_08396_),
    .B1(_08365_),
    .C1(_08368_),
    .X(_08398_));
 sky130_fd_sc_hd__o21ai_2 _21588_ (.A1(_08397_),
    .A2(_08398_),
    .B1(_08372_),
    .Y(_08399_));
 sky130_fd_sc_hd__nor3_2 _21589_ (.A(_08372_),
    .B(_08397_),
    .C(_08398_),
    .Y(_08400_));
 sky130_fd_sc_hd__nor2_2 _21590_ (.A(_11258_),
    .B(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__a22o_2 _21591_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[6] ),
    .B1(_08399_),
    .B2(_08401_),
    .X(_01736_));
 sky130_fd_sc_hd__o21ba_2 _21592_ (.A1(_08363_),
    .A2(_08393_),
    .B1_N(_08395_),
    .X(_08402_));
 sky130_fd_sc_hd__a21oi_2 _21593_ (.A1(_08373_),
    .A2(_08376_),
    .B1(_08378_),
    .Y(_08403_));
 sky130_fd_sc_hd__o21ba_2 _21594_ (.A1(_08381_),
    .A2(_08383_),
    .B1_N(_08382_),
    .X(_08404_));
 sky130_fd_sc_hd__a22o_2 _21595_ (.A1(\systolic_inst.B_outs[3][1] ),
    .A2(\systolic_inst.A_outs[3][6] ),
    .B1(\systolic_inst.A_outs[3][7] ),
    .B2(\systolic_inst.B_outs[3][0] ),
    .X(_08405_));
 sky130_fd_sc_hd__nand4_2 _21596_ (.A(\systolic_inst.B_outs[3][0] ),
    .B(\systolic_inst.B_outs[3][1] ),
    .C(\systolic_inst.A_outs[3][6] ),
    .D(\systolic_inst.A_outs[3][7] ),
    .Y(_08406_));
 sky130_fd_sc_hd__nand2_2 _21597_ (.A(_08405_),
    .B(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__xnor2_2 _21598_ (.A(_11274_),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__nor2_2 _21599_ (.A(_08404_),
    .B(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__and2_2 _21600_ (.A(_08404_),
    .B(_08408_),
    .X(_08410_));
 sky130_fd_sc_hd__nor2_2 _21601_ (.A(_08409_),
    .B(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__xnor2_2 _21602_ (.A(_08375_),
    .B(_08411_),
    .Y(_08412_));
 sky130_fd_sc_hd__nand2_2 _21603_ (.A(\systolic_inst.B_outs[3][2] ),
    .B(\systolic_inst.A_outs[3][5] ),
    .Y(_08413_));
 sky130_fd_sc_hd__and4_2 _21604_ (.A(\systolic_inst.B_outs[3][3] ),
    .B(\systolic_inst.A_outs[3][3] ),
    .C(\systolic_inst.B_outs[3][4] ),
    .D(\systolic_inst.A_outs[3][4] ),
    .X(_08414_));
 sky130_fd_sc_hd__a22oi_2 _21605_ (.A1(\systolic_inst.A_outs[3][3] ),
    .A2(\systolic_inst.B_outs[3][4] ),
    .B1(\systolic_inst.A_outs[3][4] ),
    .B2(\systolic_inst.B_outs[3][3] ),
    .Y(_08415_));
 sky130_fd_sc_hd__or2_2 _21606_ (.A(_08414_),
    .B(_08415_),
    .X(_08416_));
 sky130_fd_sc_hd__xnor2_2 _21607_ (.A(_08413_),
    .B(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__nand2_2 _21608_ (.A(\systolic_inst.A_outs[3][2] ),
    .B(\systolic_inst.B_outs[3][5] ),
    .Y(_08418_));
 sky130_fd_sc_hd__and2b_2 _21609_ (.A_N(\systolic_inst.A_outs[3][0] ),
    .B(\systolic_inst.B_outs[3][7] ),
    .X(_08419_));
 sky130_fd_sc_hd__and3_2 _21610_ (.A(\systolic_inst.A_outs[3][1] ),
    .B(\systolic_inst.B_outs[3][6] ),
    .C(_08419_),
    .X(_08420_));
 sky130_fd_sc_hd__xnor2_2 _21611_ (.A(_08387_),
    .B(_08419_),
    .Y(_08421_));
 sky130_fd_sc_hd__xnor2_2 _21612_ (.A(_08418_),
    .B(_08421_),
    .Y(_08422_));
 sky130_fd_sc_hd__xnor2_2 _21613_ (.A(_08388_),
    .B(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__nor2_2 _21614_ (.A(_08417_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__xnor2_2 _21615_ (.A(_08417_),
    .B(_08423_),
    .Y(_08425_));
 sky130_fd_sc_hd__or2_2 _21616_ (.A(_08390_),
    .B(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__and2_2 _21617_ (.A(_08390_),
    .B(_08425_),
    .X(_08427_));
 sky130_fd_sc_hd__xor2_2 _21618_ (.A(_08390_),
    .B(_08425_),
    .X(_08428_));
 sky130_fd_sc_hd__xnor2_2 _21619_ (.A(_08412_),
    .B(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__o32a_2 _21620_ (.A1(_08378_),
    .A2(_08379_),
    .A3(_08392_),
    .B1(_08391_),
    .B2(_08360_),
    .X(_08430_));
 sky130_fd_sc_hd__nand2b_2 _21621_ (.A_N(_08430_),
    .B(_08429_),
    .Y(_08431_));
 sky130_fd_sc_hd__xnor2_2 _21622_ (.A(_08429_),
    .B(_08430_),
    .Y(_08432_));
 sky130_fd_sc_hd__nand2b_2 _21623_ (.A_N(_08403_),
    .B(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__xnor2_2 _21624_ (.A(_08403_),
    .B(_08432_),
    .Y(_08434_));
 sky130_fd_sc_hd__nand2b_2 _21625_ (.A_N(_08402_),
    .B(_08434_),
    .Y(_08435_));
 sky130_fd_sc_hd__xnor2_2 _21626_ (.A(_08402_),
    .B(_08434_),
    .Y(_08436_));
 sky130_fd_sc_hd__o21ai_2 _21627_ (.A1(_08397_),
    .A2(_08400_),
    .B1(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__o31a_2 _21628_ (.A1(_08397_),
    .A2(_08400_),
    .A3(_08436_),
    .B1(\systolic_inst.ce_local ),
    .X(_08438_));
 sky130_fd_sc_hd__a22o_2 _21629_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[7] ),
    .B1(_08437_),
    .B2(_08438_),
    .X(_01737_));
 sky130_fd_sc_hd__a21o_2 _21630_ (.A1(_08375_),
    .A2(_08411_),
    .B1(_08409_),
    .X(_08439_));
 sky130_fd_sc_hd__a21bo_2 _21631_ (.A1(\systolic_inst.B_outs[3][7] ),
    .A2(_08405_),
    .B1_N(_08406_),
    .X(_08440_));
 sky130_fd_sc_hd__o21bai_2 _21632_ (.A1(_08413_),
    .A2(_08415_),
    .B1_N(_08414_),
    .Y(_08441_));
 sky130_fd_sc_hd__o21a_2 _21633_ (.A1(\systolic_inst.B_outs[3][0] ),
    .A2(\systolic_inst.B_outs[3][1] ),
    .B1(\systolic_inst.A_outs[3][7] ),
    .X(_08442_));
 sky130_fd_sc_hd__o21ai_2 _21634_ (.A1(\systolic_inst.B_outs[3][0] ),
    .A2(\systolic_inst.B_outs[3][1] ),
    .B1(\systolic_inst.A_outs[3][7] ),
    .Y(_08443_));
 sky130_fd_sc_hd__a21o_2 _21635_ (.A1(\systolic_inst.B_outs[3][0] ),
    .A2(\systolic_inst.B_outs[3][1] ),
    .B1(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__and2b_2 _21636_ (.A_N(_08444_),
    .B(_08441_),
    .X(_08445_));
 sky130_fd_sc_hd__xnor2_2 _21637_ (.A(_08441_),
    .B(_08444_),
    .Y(_08446_));
 sky130_fd_sc_hd__xnor2_2 _21638_ (.A(_08440_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__and4_2 _21639_ (.A(\systolic_inst.B_outs[3][3] ),
    .B(\systolic_inst.B_outs[3][4] ),
    .C(\systolic_inst.A_outs[3][4] ),
    .D(\systolic_inst.A_outs[3][5] ),
    .X(_08448_));
 sky130_fd_sc_hd__a22oi_2 _21640_ (.A1(\systolic_inst.B_outs[3][4] ),
    .A2(\systolic_inst.A_outs[3][4] ),
    .B1(\systolic_inst.A_outs[3][5] ),
    .B2(\systolic_inst.B_outs[3][3] ),
    .Y(_08449_));
 sky130_fd_sc_hd__nor2_2 _21641_ (.A(_08448_),
    .B(_08449_),
    .Y(_08450_));
 sky130_fd_sc_hd__nand2_2 _21642_ (.A(\systolic_inst.B_outs[3][2] ),
    .B(\systolic_inst.A_outs[3][6] ),
    .Y(_08451_));
 sky130_fd_sc_hd__xnor2_2 _21643_ (.A(_08450_),
    .B(_08451_),
    .Y(_08452_));
 sky130_fd_sc_hd__nand2_2 _21644_ (.A(\systolic_inst.A_outs[3][3] ),
    .B(\systolic_inst.B_outs[3][5] ),
    .Y(_08453_));
 sky130_fd_sc_hd__and4b_2 _21645_ (.A_N(\systolic_inst.A_outs[3][1] ),
    .B(\systolic_inst.A_outs[3][2] ),
    .C(\systolic_inst.B_outs[3][6] ),
    .D(\systolic_inst.B_outs[3][7] ),
    .X(_08454_));
 sky130_fd_sc_hd__o2bb2a_2 _21646_ (.A1_N(\systolic_inst.A_outs[3][2] ),
    .A2_N(\systolic_inst.B_outs[3][6] ),
    .B1(_11274_),
    .B2(\systolic_inst.A_outs[3][1] ),
    .X(_08455_));
 sky130_fd_sc_hd__nor2_2 _21647_ (.A(_08454_),
    .B(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__xnor2_2 _21648_ (.A(_08453_),
    .B(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__a31oi_2 _21649_ (.A1(\systolic_inst.A_outs[3][2] ),
    .A2(\systolic_inst.B_outs[3][5] ),
    .A3(_08421_),
    .B1(_08420_),
    .Y(_08458_));
 sky130_fd_sc_hd__nand2b_2 _21650_ (.A_N(_08458_),
    .B(_08457_),
    .Y(_08459_));
 sky130_fd_sc_hd__xnor2_2 _21651_ (.A(_08457_),
    .B(_08458_),
    .Y(_08460_));
 sky130_fd_sc_hd__nand2_2 _21652_ (.A(_08452_),
    .B(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__xnor2_2 _21653_ (.A(_08452_),
    .B(_08460_),
    .Y(_08462_));
 sky130_fd_sc_hd__a21oi_2 _21654_ (.A1(_08388_),
    .A2(_08422_),
    .B1(_08424_),
    .Y(_08463_));
 sky130_fd_sc_hd__xnor2_2 _21655_ (.A(_08462_),
    .B(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__or2_2 _21656_ (.A(_08447_),
    .B(_08464_),
    .X(_08465_));
 sky130_fd_sc_hd__xor2_2 _21657_ (.A(_08447_),
    .B(_08464_),
    .X(_08466_));
 sky130_fd_sc_hd__o21a_2 _21658_ (.A1(_08412_),
    .A2(_08427_),
    .B1(_08426_),
    .X(_08467_));
 sky130_fd_sc_hd__nand2b_2 _21659_ (.A_N(_08467_),
    .B(_08466_),
    .Y(_08468_));
 sky130_fd_sc_hd__xor2_2 _21660_ (.A(_08466_),
    .B(_08467_),
    .X(_08469_));
 sky130_fd_sc_hd__nand2b_2 _21661_ (.A_N(_08469_),
    .B(_08439_),
    .Y(_08470_));
 sky130_fd_sc_hd__xor2_2 _21662_ (.A(_08439_),
    .B(_08469_),
    .X(_08471_));
 sky130_fd_sc_hd__and2_2 _21663_ (.A(_08431_),
    .B(_08433_),
    .X(_08472_));
 sky130_fd_sc_hd__nor2_2 _21664_ (.A(_08471_),
    .B(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__and2_2 _21665_ (.A(_08471_),
    .B(_08472_),
    .X(_08474_));
 sky130_fd_sc_hd__nor2_2 _21666_ (.A(_08473_),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__and2_2 _21667_ (.A(_08435_),
    .B(_08437_),
    .X(_08476_));
 sky130_fd_sc_hd__and2b_2 _21668_ (.A_N(_08476_),
    .B(_08475_),
    .X(_08477_));
 sky130_fd_sc_hd__and2b_2 _21669_ (.A_N(_08475_),
    .B(_08476_),
    .X(_08478_));
 sky130_fd_sc_hd__nor2_2 _21670_ (.A(_08477_),
    .B(_08478_),
    .Y(_08479_));
 sky130_fd_sc_hd__mux2_1 _21671_ (.A0(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[8] ),
    .A1(_08479_),
    .S(\systolic_inst.ce_local ),
    .X(_01738_));
 sky130_fd_sc_hd__a21o_2 _21672_ (.A1(_08440_),
    .A2(_08446_),
    .B1(_08445_),
    .X(_08480_));
 sky130_fd_sc_hd__o21ba_2 _21673_ (.A1(_08449_),
    .A2(_08451_),
    .B1_N(_08448_),
    .X(_08481_));
 sky130_fd_sc_hd__nor2_2 _21674_ (.A(_08443_),
    .B(_08481_),
    .Y(_08482_));
 sky130_fd_sc_hd__and2_2 _21675_ (.A(_08443_),
    .B(_08481_),
    .X(_08483_));
 sky130_fd_sc_hd__or2_2 _21676_ (.A(_08482_),
    .B(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__nand2_2 _21677_ (.A(\systolic_inst.B_outs[3][2] ),
    .B(\systolic_inst.A_outs[3][7] ),
    .Y(_08485_));
 sky130_fd_sc_hd__a22oi_2 _21678_ (.A1(\systolic_inst.B_outs[3][4] ),
    .A2(\systolic_inst.A_outs[3][5] ),
    .B1(\systolic_inst.A_outs[3][6] ),
    .B2(\systolic_inst.B_outs[3][3] ),
    .Y(_08486_));
 sky130_fd_sc_hd__and4_2 _21679_ (.A(\systolic_inst.B_outs[3][3] ),
    .B(\systolic_inst.B_outs[3][4] ),
    .C(\systolic_inst.A_outs[3][5] ),
    .D(\systolic_inst.A_outs[3][6] ),
    .X(_08487_));
 sky130_fd_sc_hd__nor2_2 _21680_ (.A(_08486_),
    .B(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__xnor2_2 _21681_ (.A(_08485_),
    .B(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__nand2_2 _21682_ (.A(\systolic_inst.A_outs[3][4] ),
    .B(\systolic_inst.B_outs[3][5] ),
    .Y(_08490_));
 sky130_fd_sc_hd__and4b_2 _21683_ (.A_N(\systolic_inst.A_outs[3][2] ),
    .B(\systolic_inst.A_outs[3][3] ),
    .C(\systolic_inst.B_outs[3][6] ),
    .D(\systolic_inst.B_outs[3][7] ),
    .X(_08491_));
 sky130_fd_sc_hd__o2bb2a_2 _21684_ (.A1_N(\systolic_inst.A_outs[3][3] ),
    .A2_N(\systolic_inst.B_outs[3][6] ),
    .B1(_11274_),
    .B2(\systolic_inst.A_outs[3][2] ),
    .X(_08492_));
 sky130_fd_sc_hd__nor2_2 _21685_ (.A(_08491_),
    .B(_08492_),
    .Y(_08493_));
 sky130_fd_sc_hd__xnor2_2 _21686_ (.A(_08490_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__o21ba_2 _21687_ (.A1(_08453_),
    .A2(_08455_),
    .B1_N(_08454_),
    .X(_08495_));
 sky130_fd_sc_hd__nand2b_2 _21688_ (.A_N(_08495_),
    .B(_08494_),
    .Y(_08496_));
 sky130_fd_sc_hd__xnor2_2 _21689_ (.A(_08494_),
    .B(_08495_),
    .Y(_08497_));
 sky130_fd_sc_hd__xnor2_2 _21690_ (.A(_08489_),
    .B(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__a21o_2 _21691_ (.A1(_08459_),
    .A2(_08461_),
    .B1(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__nand3_2 _21692_ (.A(_08459_),
    .B(_08461_),
    .C(_08498_),
    .Y(_08500_));
 sky130_fd_sc_hd__nand2_2 _21693_ (.A(_08499_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__xor2_2 _21694_ (.A(_08484_),
    .B(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__o21a_2 _21695_ (.A1(_08462_),
    .A2(_08463_),
    .B1(_08465_),
    .X(_08503_));
 sky130_fd_sc_hd__nand2b_2 _21696_ (.A_N(_08503_),
    .B(_08502_),
    .Y(_08504_));
 sky130_fd_sc_hd__xnor2_2 _21697_ (.A(_08502_),
    .B(_08503_),
    .Y(_08505_));
 sky130_fd_sc_hd__xnor2_2 _21698_ (.A(_08480_),
    .B(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__a21oi_2 _21699_ (.A1(_08468_),
    .A2(_08470_),
    .B1(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__and3_2 _21700_ (.A(_08468_),
    .B(_08470_),
    .C(_08506_),
    .X(_08508_));
 sky130_fd_sc_hd__inv_2 _21701_ (.A(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__nor2_2 _21702_ (.A(_08507_),
    .B(_08508_),
    .Y(_08510_));
 sky130_fd_sc_hd__or3_2 _21703_ (.A(_08473_),
    .B(_08477_),
    .C(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__o21ai_2 _21704_ (.A1(_08473_),
    .A2(_08477_),
    .B1(_08510_),
    .Y(_08512_));
 sky130_fd_sc_hd__and2_2 _21705_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[9] ),
    .X(_08513_));
 sky130_fd_sc_hd__a31o_2 _21706_ (.A1(\systolic_inst.ce_local ),
    .A2(_08511_),
    .A3(_08512_),
    .B1(_08513_),
    .X(_01739_));
 sky130_fd_sc_hd__o21ba_2 _21707_ (.A1(_08485_),
    .A2(_08486_),
    .B1_N(_08487_),
    .X(_08514_));
 sky130_fd_sc_hd__nor2_2 _21708_ (.A(_08443_),
    .B(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__and2_2 _21709_ (.A(_08443_),
    .B(_08514_),
    .X(_08516_));
 sky130_fd_sc_hd__or2_2 _21710_ (.A(_08515_),
    .B(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__a22o_2 _21711_ (.A1(\systolic_inst.B_outs[3][4] ),
    .A2(\systolic_inst.A_outs[3][6] ),
    .B1(\systolic_inst.A_outs[3][7] ),
    .B2(\systolic_inst.B_outs[3][3] ),
    .X(_08518_));
 sky130_fd_sc_hd__and3_2 _21712_ (.A(\systolic_inst.B_outs[3][3] ),
    .B(\systolic_inst.B_outs[3][4] ),
    .C(\systolic_inst.A_outs[3][7] ),
    .X(_08519_));
 sky130_fd_sc_hd__a21bo_2 _21713_ (.A1(\systolic_inst.A_outs[3][6] ),
    .A2(_08519_),
    .B1_N(_08518_),
    .X(_08520_));
 sky130_fd_sc_hd__xor2_2 _21714_ (.A(_08485_),
    .B(_08520_),
    .X(_08521_));
 sky130_fd_sc_hd__nand2_2 _21715_ (.A(\systolic_inst.B_outs[3][5] ),
    .B(\systolic_inst.A_outs[3][5] ),
    .Y(_08522_));
 sky130_fd_sc_hd__and4b_2 _21716_ (.A_N(\systolic_inst.A_outs[3][3] ),
    .B(\systolic_inst.A_outs[3][4] ),
    .C(\systolic_inst.B_outs[3][6] ),
    .D(\systolic_inst.B_outs[3][7] ),
    .X(_08523_));
 sky130_fd_sc_hd__o2bb2a_2 _21717_ (.A1_N(\systolic_inst.A_outs[3][4] ),
    .A2_N(\systolic_inst.B_outs[3][6] ),
    .B1(_11274_),
    .B2(\systolic_inst.A_outs[3][3] ),
    .X(_08524_));
 sky130_fd_sc_hd__nor2_2 _21718_ (.A(_08523_),
    .B(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__xnor2_2 _21719_ (.A(_08522_),
    .B(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__o21ba_2 _21720_ (.A1(_08490_),
    .A2(_08492_),
    .B1_N(_08491_),
    .X(_08527_));
 sky130_fd_sc_hd__nand2b_2 _21721_ (.A_N(_08527_),
    .B(_08526_),
    .Y(_08528_));
 sky130_fd_sc_hd__xnor2_2 _21722_ (.A(_08526_),
    .B(_08527_),
    .Y(_08529_));
 sky130_fd_sc_hd__nand2_2 _21723_ (.A(_08521_),
    .B(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__or2_2 _21724_ (.A(_08521_),
    .B(_08529_),
    .X(_08531_));
 sky130_fd_sc_hd__nand2_2 _21725_ (.A(_08530_),
    .B(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__a21bo_2 _21726_ (.A1(_08489_),
    .A2(_08497_),
    .B1_N(_08496_),
    .X(_08533_));
 sky130_fd_sc_hd__nand2b_2 _21727_ (.A_N(_08532_),
    .B(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__xor2_2 _21728_ (.A(_08532_),
    .B(_08533_),
    .X(_08535_));
 sky130_fd_sc_hd__xor2_2 _21729_ (.A(_08517_),
    .B(_08535_),
    .X(_08536_));
 sky130_fd_sc_hd__o21a_2 _21730_ (.A1(_08484_),
    .A2(_08501_),
    .B1(_08499_),
    .X(_08537_));
 sky130_fd_sc_hd__nand2b_2 _21731_ (.A_N(_08537_),
    .B(_08536_),
    .Y(_08538_));
 sky130_fd_sc_hd__xnor2_2 _21732_ (.A(_08536_),
    .B(_08537_),
    .Y(_08539_));
 sky130_fd_sc_hd__nand2_2 _21733_ (.A(_08482_),
    .B(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__or2_2 _21734_ (.A(_08482_),
    .B(_08539_),
    .X(_08541_));
 sky130_fd_sc_hd__nand2_2 _21735_ (.A(_08540_),
    .B(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__a21boi_2 _21736_ (.A1(_08480_),
    .A2(_08505_),
    .B1_N(_08504_),
    .Y(_08543_));
 sky130_fd_sc_hd__nor2_2 _21737_ (.A(_08542_),
    .B(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__xor2_2 _21738_ (.A(_08542_),
    .B(_08543_),
    .X(_08545_));
 sky130_fd_sc_hd__o31a_2 _21739_ (.A1(_08473_),
    .A2(_08477_),
    .A3(_08507_),
    .B1(_08509_),
    .X(_08546_));
 sky130_fd_sc_hd__or2_2 _21740_ (.A(_08545_),
    .B(_08546_),
    .X(_08547_));
 sky130_fd_sc_hd__o311a_2 _21741_ (.A1(_08473_),
    .A2(_08477_),
    .A3(_08507_),
    .B1(_08509_),
    .C1(_08545_),
    .X(_08548_));
 sky130_fd_sc_hd__nor2_2 _21742_ (.A(_11258_),
    .B(_08548_),
    .Y(_08549_));
 sky130_fd_sc_hd__a22o_2 _21743_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[10] ),
    .B1(_08547_),
    .B2(_08549_),
    .X(_01740_));
 sky130_fd_sc_hd__o2bb2a_2 _21744_ (.A1_N(\systolic_inst.A_outs[3][6] ),
    .A2_N(_08519_),
    .B1(_08520_),
    .B2(_08485_),
    .X(_08550_));
 sky130_fd_sc_hd__or2_2 _21745_ (.A(_08443_),
    .B(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__nand2_2 _21746_ (.A(_08443_),
    .B(_08550_),
    .Y(_08552_));
 sky130_fd_sc_hd__nand2_2 _21747_ (.A(_08551_),
    .B(_08552_),
    .Y(_08553_));
 sky130_fd_sc_hd__or2_2 _21748_ (.A(\systolic_inst.B_outs[3][3] ),
    .B(\systolic_inst.B_outs[3][4] ),
    .X(_08554_));
 sky130_fd_sc_hd__and3b_2 _21749_ (.A_N(_08519_),
    .B(_08554_),
    .C(\systolic_inst.A_outs[3][7] ),
    .X(_08555_));
 sky130_fd_sc_hd__xnor2_2 _21750_ (.A(_08485_),
    .B(_08555_),
    .Y(_08556_));
 sky130_fd_sc_hd__nand2_2 _21751_ (.A(\systolic_inst.B_outs[3][5] ),
    .B(\systolic_inst.A_outs[3][6] ),
    .Y(_08557_));
 sky130_fd_sc_hd__and4b_2 _21752_ (.A_N(\systolic_inst.A_outs[3][4] ),
    .B(\systolic_inst.A_outs[3][5] ),
    .C(\systolic_inst.B_outs[3][6] ),
    .D(\systolic_inst.B_outs[3][7] ),
    .X(_08558_));
 sky130_fd_sc_hd__o2bb2a_2 _21753_ (.A1_N(\systolic_inst.A_outs[3][5] ),
    .A2_N(\systolic_inst.B_outs[3][6] ),
    .B1(_11274_),
    .B2(\systolic_inst.A_outs[3][4] ),
    .X(_08559_));
 sky130_fd_sc_hd__nor2_2 _21754_ (.A(_08558_),
    .B(_08559_),
    .Y(_08560_));
 sky130_fd_sc_hd__xnor2_2 _21755_ (.A(_08557_),
    .B(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__o21ba_2 _21756_ (.A1(_08522_),
    .A2(_08524_),
    .B1_N(_08523_),
    .X(_08562_));
 sky130_fd_sc_hd__nand2b_2 _21757_ (.A_N(_08562_),
    .B(_08561_),
    .Y(_08563_));
 sky130_fd_sc_hd__xnor2_2 _21758_ (.A(_08561_),
    .B(_08562_),
    .Y(_08564_));
 sky130_fd_sc_hd__nand2_2 _21759_ (.A(_08556_),
    .B(_08564_),
    .Y(_08565_));
 sky130_fd_sc_hd__xnor2_2 _21760_ (.A(_08556_),
    .B(_08564_),
    .Y(_08566_));
 sky130_fd_sc_hd__a21o_2 _21761_ (.A1(_08528_),
    .A2(_08530_),
    .B1(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__nand3_2 _21762_ (.A(_08528_),
    .B(_08530_),
    .C(_08566_),
    .Y(_08568_));
 sky130_fd_sc_hd__nand2_2 _21763_ (.A(_08567_),
    .B(_08568_),
    .Y(_08569_));
 sky130_fd_sc_hd__xor2_2 _21764_ (.A(_08553_),
    .B(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__o21a_2 _21765_ (.A1(_08517_),
    .A2(_08535_),
    .B1(_08534_),
    .X(_08571_));
 sky130_fd_sc_hd__and2b_2 _21766_ (.A_N(_08571_),
    .B(_08570_),
    .X(_08572_));
 sky130_fd_sc_hd__xnor2_2 _21767_ (.A(_08570_),
    .B(_08571_),
    .Y(_08573_));
 sky130_fd_sc_hd__xnor2_2 _21768_ (.A(_08515_),
    .B(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__and3_2 _21769_ (.A(_08538_),
    .B(_08540_),
    .C(_08574_),
    .X(_08575_));
 sky130_fd_sc_hd__inv_2 _21770_ (.A(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__a21oi_2 _21771_ (.A1(_08538_),
    .A2(_08540_),
    .B1(_08574_),
    .Y(_08577_));
 sky130_fd_sc_hd__nor2_2 _21772_ (.A(_08575_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__or3_2 _21773_ (.A(_08544_),
    .B(_08548_),
    .C(_08578_),
    .X(_08579_));
 sky130_fd_sc_hd__o21ai_2 _21774_ (.A1(_08544_),
    .A2(_08548_),
    .B1(_08578_),
    .Y(_08580_));
 sky130_fd_sc_hd__and2_2 _21775_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[11] ),
    .X(_08581_));
 sky130_fd_sc_hd__a31o_2 _21776_ (.A1(\systolic_inst.ce_local ),
    .A2(_08579_),
    .A3(_08580_),
    .B1(_08581_),
    .X(_01741_));
 sky130_fd_sc_hd__a31o_2 _21777_ (.A1(\systolic_inst.B_outs[3][2] ),
    .A2(\systolic_inst.A_outs[3][7] ),
    .A3(_08554_),
    .B1(_08519_),
    .X(_08582_));
 sky130_fd_sc_hd__or2_2 _21778_ (.A(_08442_),
    .B(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__nand2_2 _21779_ (.A(_08442_),
    .B(_08582_),
    .Y(_08584_));
 sky130_fd_sc_hd__nand2_2 _21780_ (.A(_08583_),
    .B(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__inv_2 _21781_ (.A(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__o2bb2a_2 _21782_ (.A1_N(\systolic_inst.B_outs[3][6] ),
    .A2_N(\systolic_inst.A_outs[3][6] ),
    .B1(_11274_),
    .B2(\systolic_inst.A_outs[3][5] ),
    .X(_08587_));
 sky130_fd_sc_hd__and4b_2 _21783_ (.A_N(\systolic_inst.A_outs[3][5] ),
    .B(\systolic_inst.B_outs[3][6] ),
    .C(\systolic_inst.A_outs[3][6] ),
    .D(\systolic_inst.B_outs[3][7] ),
    .X(_08588_));
 sky130_fd_sc_hd__nor2_2 _21784_ (.A(_08587_),
    .B(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__nand2_2 _21785_ (.A(\systolic_inst.B_outs[3][5] ),
    .B(\systolic_inst.A_outs[3][7] ),
    .Y(_08590_));
 sky130_fd_sc_hd__and3_2 _21786_ (.A(\systolic_inst.B_outs[3][5] ),
    .B(\systolic_inst.A_outs[3][7] ),
    .C(_08589_),
    .X(_08591_));
 sky130_fd_sc_hd__xnor2_2 _21787_ (.A(_08589_),
    .B(_08590_),
    .Y(_08592_));
 sky130_fd_sc_hd__o21ba_2 _21788_ (.A1(_08557_),
    .A2(_08559_),
    .B1_N(_08558_),
    .X(_08593_));
 sky130_fd_sc_hd__nand2b_2 _21789_ (.A_N(_08593_),
    .B(_08592_),
    .Y(_08594_));
 sky130_fd_sc_hd__xnor2_2 _21790_ (.A(_08592_),
    .B(_08593_),
    .Y(_08595_));
 sky130_fd_sc_hd__xnor2_2 _21791_ (.A(_08556_),
    .B(_08595_),
    .Y(_08596_));
 sky130_fd_sc_hd__a21o_2 _21792_ (.A1(_08563_),
    .A2(_08565_),
    .B1(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__nand3_2 _21793_ (.A(_08563_),
    .B(_08565_),
    .C(_08596_),
    .Y(_08598_));
 sky130_fd_sc_hd__nand2_2 _21794_ (.A(_08597_),
    .B(_08598_),
    .Y(_08599_));
 sky130_fd_sc_hd__xnor2_2 _21795_ (.A(_08586_),
    .B(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__o21a_2 _21796_ (.A1(_08553_),
    .A2(_08569_),
    .B1(_08567_),
    .X(_08601_));
 sky130_fd_sc_hd__and2b_2 _21797_ (.A_N(_08601_),
    .B(_08600_),
    .X(_08602_));
 sky130_fd_sc_hd__xnor2_2 _21798_ (.A(_08600_),
    .B(_08601_),
    .Y(_08603_));
 sky130_fd_sc_hd__and2b_2 _21799_ (.A_N(_08551_),
    .B(_08603_),
    .X(_08604_));
 sky130_fd_sc_hd__xor2_2 _21800_ (.A(_08551_),
    .B(_08603_),
    .X(_08605_));
 sky130_fd_sc_hd__a21oi_2 _21801_ (.A1(_08515_),
    .A2(_08573_),
    .B1(_08572_),
    .Y(_08606_));
 sky130_fd_sc_hd__nor2_2 _21802_ (.A(_08605_),
    .B(_08606_),
    .Y(_08607_));
 sky130_fd_sc_hd__and2_2 _21803_ (.A(_08605_),
    .B(_08606_),
    .X(_08608_));
 sky130_fd_sc_hd__or2_2 _21804_ (.A(_08607_),
    .B(_08608_),
    .X(_08609_));
 sky130_fd_sc_hd__inv_2 _21805_ (.A(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__o31a_2 _21806_ (.A1(_08544_),
    .A2(_08548_),
    .A3(_08577_),
    .B1(_08576_),
    .X(_08611_));
 sky130_fd_sc_hd__o311a_2 _21807_ (.A1(_08544_),
    .A2(_08548_),
    .A3(_08577_),
    .B1(_08610_),
    .C1(_08576_),
    .X(_08612_));
 sky130_fd_sc_hd__nor2_2 _21808_ (.A(_08610_),
    .B(_08611_),
    .Y(_08613_));
 sky130_fd_sc_hd__nor2_2 _21809_ (.A(_08612_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__mux2_1 _21810_ (.A0(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[12] ),
    .A1(_08614_),
    .S(\systolic_inst.ce_local ),
    .X(_01742_));
 sky130_fd_sc_hd__nand2_2 _21811_ (.A(\systolic_inst.B_outs[3][6] ),
    .B(\systolic_inst.A_outs[3][7] ),
    .Y(_08615_));
 sky130_fd_sc_hd__nor2_2 _21812_ (.A(\systolic_inst.A_outs[3][6] ),
    .B(_11274_),
    .Y(_08616_));
 sky130_fd_sc_hd__xnor2_2 _21813_ (.A(_08615_),
    .B(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__nand2b_2 _21814_ (.A_N(_08590_),
    .B(_08617_),
    .Y(_08618_));
 sky130_fd_sc_hd__xnor2_2 _21815_ (.A(_08590_),
    .B(_08617_),
    .Y(_08619_));
 sky130_fd_sc_hd__o21ai_2 _21816_ (.A1(_08588_),
    .A2(_08591_),
    .B1(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__or3_2 _21817_ (.A(_08588_),
    .B(_08591_),
    .C(_08619_),
    .X(_08621_));
 sky130_fd_sc_hd__and2_2 _21818_ (.A(_08620_),
    .B(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__nand2_2 _21819_ (.A(_08556_),
    .B(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__or2_2 _21820_ (.A(_08556_),
    .B(_08622_),
    .X(_08624_));
 sky130_fd_sc_hd__nand2_2 _21821_ (.A(_08623_),
    .B(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__a21bo_2 _21822_ (.A1(_08556_),
    .A2(_08595_),
    .B1_N(_08594_),
    .X(_08626_));
 sky130_fd_sc_hd__nand2b_2 _21823_ (.A_N(_08625_),
    .B(_08626_),
    .Y(_08627_));
 sky130_fd_sc_hd__xor2_2 _21824_ (.A(_08625_),
    .B(_08626_),
    .X(_08628_));
 sky130_fd_sc_hd__xnor2_2 _21825_ (.A(_08586_),
    .B(_08628_),
    .Y(_08629_));
 sky130_fd_sc_hd__o21a_2 _21826_ (.A1(_08585_),
    .A2(_08599_),
    .B1(_08597_),
    .X(_08630_));
 sky130_fd_sc_hd__and2b_2 _21827_ (.A_N(_08630_),
    .B(_08629_),
    .X(_08631_));
 sky130_fd_sc_hd__and2b_2 _21828_ (.A_N(_08629_),
    .B(_08630_),
    .X(_08632_));
 sky130_fd_sc_hd__nor2_2 _21829_ (.A(_08631_),
    .B(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__xnor2_2 _21830_ (.A(_08584_),
    .B(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__nor3_2 _21831_ (.A(_08602_),
    .B(_08604_),
    .C(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__o21a_2 _21832_ (.A1(_08602_),
    .A2(_08604_),
    .B1(_08634_),
    .X(_08636_));
 sky130_fd_sc_hd__nor2_2 _21833_ (.A(_08635_),
    .B(_08636_),
    .Y(_08637_));
 sky130_fd_sc_hd__o21ai_2 _21834_ (.A1(_08607_),
    .A2(_08612_),
    .B1(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__o31a_2 _21835_ (.A1(_08607_),
    .A2(_08612_),
    .A3(_08637_),
    .B1(\systolic_inst.ce_local ),
    .X(_08639_));
 sky130_fd_sc_hd__a22o_2 _21836_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[13] ),
    .B1(_08638_),
    .B2(_08639_),
    .X(_01743_));
 sky130_fd_sc_hd__o211ai_2 _21837_ (.A1(_11274_),
    .A2(\systolic_inst.A_outs[3][7] ),
    .B1(_08590_),
    .C1(_08615_),
    .Y(_08640_));
 sky130_fd_sc_hd__o311a_2 _21838_ (.A1(\systolic_inst.A_outs[3][6] ),
    .A2(_11274_),
    .A3(_08615_),
    .B1(_08618_),
    .C1(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__a31o_2 _21839_ (.A1(\systolic_inst.B_outs[3][5] ),
    .A2(\systolic_inst.B_outs[3][6] ),
    .A3(\systolic_inst.A_outs[3][7] ),
    .B1(_08641_),
    .X(_08642_));
 sky130_fd_sc_hd__nor2_2 _21840_ (.A(_08556_),
    .B(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__and2_2 _21841_ (.A(_08556_),
    .B(_08642_),
    .X(_08644_));
 sky130_fd_sc_hd__or2_2 _21842_ (.A(_08643_),
    .B(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__a21oi_2 _21843_ (.A1(_08620_),
    .A2(_08623_),
    .B1(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__and3_2 _21844_ (.A(_08620_),
    .B(_08623_),
    .C(_08645_),
    .X(_08647_));
 sky130_fd_sc_hd__nor2_2 _21845_ (.A(_08646_),
    .B(_08647_),
    .Y(_08648_));
 sky130_fd_sc_hd__xnor2_2 _21846_ (.A(_08585_),
    .B(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__o21a_2 _21847_ (.A1(_08585_),
    .A2(_08628_),
    .B1(_08627_),
    .X(_08650_));
 sky130_fd_sc_hd__and2b_2 _21848_ (.A_N(_08650_),
    .B(_08649_),
    .X(_08651_));
 sky130_fd_sc_hd__and2b_2 _21849_ (.A_N(_08649_),
    .B(_08650_),
    .X(_08652_));
 sky130_fd_sc_hd__nor2_2 _21850_ (.A(_08651_),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__xnor2_2 _21851_ (.A(_08584_),
    .B(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__o21ba_2 _21852_ (.A1(_08584_),
    .A2(_08632_),
    .B1_N(_08631_),
    .X(_08655_));
 sky130_fd_sc_hd__nand2b_2 _21853_ (.A_N(_08655_),
    .B(_08654_),
    .Y(_08656_));
 sky130_fd_sc_hd__xnor2_2 _21854_ (.A(_08654_),
    .B(_08655_),
    .Y(_08657_));
 sky130_fd_sc_hd__nor2_2 _21855_ (.A(_08607_),
    .B(_08636_),
    .Y(_08658_));
 sky130_fd_sc_hd__a2bb2o_2 _21856_ (.A1_N(_08635_),
    .A2_N(_08658_),
    .B1(_08637_),
    .B2(_08612_),
    .X(_08659_));
 sky130_fd_sc_hd__nand2_2 _21857_ (.A(_08657_),
    .B(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__xor2_2 _21858_ (.A(_08657_),
    .B(_08659_),
    .X(_08661_));
 sky130_fd_sc_hd__mux2_1 _21859_ (.A0(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[14] ),
    .A1(_08661_),
    .S(\systolic_inst.ce_local ),
    .X(_01744_));
 sky130_fd_sc_hd__a31oi_2 _21860_ (.A1(_08442_),
    .A2(_08582_),
    .A3(_08653_),
    .B1(_08651_),
    .Y(_08662_));
 sky130_fd_sc_hd__a21oi_2 _21861_ (.A1(_08586_),
    .A2(_08648_),
    .B1(_08646_),
    .Y(_08663_));
 sky130_fd_sc_hd__xnor2_2 _21862_ (.A(_08583_),
    .B(_08643_),
    .Y(_08664_));
 sky130_fd_sc_hd__xnor2_2 _21863_ (.A(_08663_),
    .B(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__xnor2_2 _21864_ (.A(_08662_),
    .B(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__and3_2 _21865_ (.A(\systolic_inst.ce_local ),
    .B(_08656_),
    .C(_08666_),
    .X(_08667_));
 sky130_fd_sc_hd__a22o_2 _21866_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B1(_08660_),
    .B2(_08667_),
    .X(_01745_));
 sky130_fd_sc_hd__a21o_2 _21867_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[3][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_08668_));
 sky130_fd_sc_hd__a21oi_2 _21868_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[3][0] ),
    .Y(_08669_));
 sky130_fd_sc_hd__a21oi_2 _21869_ (.A1(\systolic_inst.ce_local ),
    .A2(_08668_),
    .B1(_08669_),
    .Y(_01746_));
 sky130_fd_sc_hd__and2_2 _21870_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[3][1] ),
    .X(_08670_));
 sky130_fd_sc_hd__nand2_2 _21871_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[3][1] ),
    .Y(_08671_));
 sky130_fd_sc_hd__or2_2 _21872_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[3][1] ),
    .X(_08672_));
 sky130_fd_sc_hd__and4_2 _21873_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[3][0] ),
    .C(_08671_),
    .D(_08672_),
    .X(_08673_));
 sky130_fd_sc_hd__inv_2 _21874_ (.A(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__a22o_2 _21875_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[3][0] ),
    .B1(_08671_),
    .B2(_08672_),
    .X(_08675_));
 sky130_fd_sc_hd__a32o_2 _21876_ (.A1(_11712_),
    .A2(_08674_),
    .A3(_08675_),
    .B1(\systolic_inst.acc_wires[3][1] ),
    .B2(_11258_),
    .X(_01747_));
 sky130_fd_sc_hd__and2_2 _21877_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[3][2] ),
    .X(_08676_));
 sky130_fd_sc_hd__nand2_2 _21878_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[3][2] ),
    .Y(_08677_));
 sky130_fd_sc_hd__or2_2 _21879_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[3][2] ),
    .X(_08678_));
 sky130_fd_sc_hd__a211o_2 _21880_ (.A1(_08677_),
    .A2(_08678_),
    .B1(_08670_),
    .C1(_08673_),
    .X(_08679_));
 sky130_fd_sc_hd__o211a_2 _21881_ (.A1(_08670_),
    .A2(_08673_),
    .B1(_08677_),
    .C1(_08678_),
    .X(_08680_));
 sky130_fd_sc_hd__inv_2 _21882_ (.A(_08680_),
    .Y(_08681_));
 sky130_fd_sc_hd__a32o_2 _21883_ (.A1(_11712_),
    .A2(_08679_),
    .A3(_08681_),
    .B1(\systolic_inst.acc_wires[3][2] ),
    .B2(_11258_),
    .X(_01748_));
 sky130_fd_sc_hd__and2_2 _21884_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[3][3] ),
    .X(_08682_));
 sky130_fd_sc_hd__nand2_2 _21885_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[3][3] ),
    .Y(_08683_));
 sky130_fd_sc_hd__or2_2 _21886_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[3][3] ),
    .X(_08684_));
 sky130_fd_sc_hd__a211o_2 _21887_ (.A1(_08683_),
    .A2(_08684_),
    .B1(_08676_),
    .C1(_08680_),
    .X(_08685_));
 sky130_fd_sc_hd__o211a_2 _21888_ (.A1(_08676_),
    .A2(_08680_),
    .B1(_08683_),
    .C1(_08684_),
    .X(_08686_));
 sky130_fd_sc_hd__inv_2 _21889_ (.A(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__a32o_2 _21890_ (.A1(_11712_),
    .A2(_08685_),
    .A3(_08687_),
    .B1(\systolic_inst.acc_wires[3][3] ),
    .B2(_11258_),
    .X(_01749_));
 sky130_fd_sc_hd__and2_2 _21891_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[3][4] ),
    .X(_08688_));
 sky130_fd_sc_hd__nand2_2 _21892_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[3][4] ),
    .Y(_08689_));
 sky130_fd_sc_hd__or2_2 _21893_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[3][4] ),
    .X(_08690_));
 sky130_fd_sc_hd__a211o_2 _21894_ (.A1(_08689_),
    .A2(_08690_),
    .B1(_08682_),
    .C1(_08686_),
    .X(_08691_));
 sky130_fd_sc_hd__o211a_2 _21895_ (.A1(_08682_),
    .A2(_08686_),
    .B1(_08689_),
    .C1(_08690_),
    .X(_08692_));
 sky130_fd_sc_hd__inv_2 _21896_ (.A(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__a32o_2 _21897_ (.A1(_11712_),
    .A2(_08691_),
    .A3(_08693_),
    .B1(\systolic_inst.acc_wires[3][4] ),
    .B2(_11258_),
    .X(_01750_));
 sky130_fd_sc_hd__and2_2 _21898_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[3][5] ),
    .X(_08694_));
 sky130_fd_sc_hd__nand2_2 _21899_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[3][5] ),
    .Y(_08695_));
 sky130_fd_sc_hd__or2_2 _21900_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[3][5] ),
    .X(_08696_));
 sky130_fd_sc_hd__a211o_2 _21901_ (.A1(_08695_),
    .A2(_08696_),
    .B1(_08688_),
    .C1(_08692_),
    .X(_08697_));
 sky130_fd_sc_hd__o211a_2 _21902_ (.A1(_08688_),
    .A2(_08692_),
    .B1(_08695_),
    .C1(_08696_),
    .X(_08698_));
 sky130_fd_sc_hd__inv_2 _21903_ (.A(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__a32o_2 _21904_ (.A1(_11712_),
    .A2(_08697_),
    .A3(_08699_),
    .B1(\systolic_inst.acc_wires[3][5] ),
    .B2(_11258_),
    .X(_01751_));
 sky130_fd_sc_hd__nand2_2 _21905_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[3][6] ),
    .Y(_08700_));
 sky130_fd_sc_hd__inv_2 _21906_ (.A(_08700_),
    .Y(_08701_));
 sky130_fd_sc_hd__or2_2 _21907_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[3][6] ),
    .X(_08702_));
 sky130_fd_sc_hd__a211o_2 _21908_ (.A1(_08700_),
    .A2(_08702_),
    .B1(_08694_),
    .C1(_08698_),
    .X(_08703_));
 sky130_fd_sc_hd__o211a_2 _21909_ (.A1(_08694_),
    .A2(_08698_),
    .B1(_08700_),
    .C1(_08702_),
    .X(_08704_));
 sky130_fd_sc_hd__inv_2 _21910_ (.A(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__a32o_2 _21911_ (.A1(_11712_),
    .A2(_08703_),
    .A3(_08705_),
    .B1(\systolic_inst.acc_wires[3][6] ),
    .B2(_11258_),
    .X(_01752_));
 sky130_fd_sc_hd__nand2_2 _21912_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[3][7] ),
    .Y(_08706_));
 sky130_fd_sc_hd__or2_2 _21913_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[3][7] ),
    .X(_08707_));
 sky130_fd_sc_hd__a211o_2 _21914_ (.A1(_08706_),
    .A2(_08707_),
    .B1(_08701_),
    .C1(_08704_),
    .X(_08708_));
 sky130_fd_sc_hd__o211ai_2 _21915_ (.A1(_08701_),
    .A2(_08704_),
    .B1(_08706_),
    .C1(_08707_),
    .Y(_08709_));
 sky130_fd_sc_hd__a32o_2 _21916_ (.A1(_11712_),
    .A2(_08708_),
    .A3(_08709_),
    .B1(\systolic_inst.acc_wires[3][7] ),
    .B2(_11258_),
    .X(_01753_));
 sky130_fd_sc_hd__xnor2_2 _21917_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[3][8] ),
    .Y(_08710_));
 sky130_fd_sc_hd__a21oi_2 _21918_ (.A1(_08706_),
    .A2(_08709_),
    .B1(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__a31o_2 _21919_ (.A1(_08706_),
    .A2(_08709_),
    .A3(_08710_),
    .B1(_11713_),
    .X(_08712_));
 sky130_fd_sc_hd__a2bb2o_2 _21920_ (.A1_N(_08712_),
    .A2_N(_08711_),
    .B1(\systolic_inst.acc_wires[3][8] ),
    .B2(_11258_),
    .X(_01754_));
 sky130_fd_sc_hd__nor2_2 _21921_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[3][9] ),
    .Y(_08713_));
 sky130_fd_sc_hd__and2_2 _21922_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[3][9] ),
    .X(_08714_));
 sky130_fd_sc_hd__nor2_2 _21923_ (.A(_08713_),
    .B(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__a21oi_2 _21924_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[3][8] ),
    .B1(_08711_),
    .Y(_08716_));
 sky130_fd_sc_hd__xnor2_2 _21925_ (.A(_08715_),
    .B(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__a22o_2 _21926_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[3][9] ),
    .B1(_11712_),
    .B2(_08717_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_2 _21927_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[3][10] ),
    .Y(_08718_));
 sky130_fd_sc_hd__or2_2 _21928_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[3][10] ),
    .X(_08719_));
 sky130_fd_sc_hd__and2_2 _21929_ (.A(_08718_),
    .B(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__a31o_2 _21930_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[3][8] ),
    .A3(_08715_),
    .B1(_08714_),
    .X(_08721_));
 sky130_fd_sc_hd__a21o_2 _21931_ (.A1(_08711_),
    .A2(_08715_),
    .B1(_08721_),
    .X(_08722_));
 sky130_fd_sc_hd__or2_2 _21932_ (.A(_08720_),
    .B(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__nand2_2 _21933_ (.A(_08720_),
    .B(_08722_),
    .Y(_08724_));
 sky130_fd_sc_hd__a32o_2 _21934_ (.A1(_11712_),
    .A2(_08723_),
    .A3(_08724_),
    .B1(\systolic_inst.acc_wires[3][10] ),
    .B2(_11258_),
    .X(_01756_));
 sky130_fd_sc_hd__or2_2 _21935_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[3][11] ),
    .X(_08725_));
 sky130_fd_sc_hd__nand2_2 _21936_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[3][11] ),
    .Y(_08726_));
 sky130_fd_sc_hd__inv_2 _21937_ (.A(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__nand2_2 _21938_ (.A(_08725_),
    .B(_08726_),
    .Y(_08728_));
 sky130_fd_sc_hd__a21o_2 _21939_ (.A1(_08718_),
    .A2(_08724_),
    .B1(_08728_),
    .X(_08729_));
 sky130_fd_sc_hd__a31oi_2 _21940_ (.A1(_08718_),
    .A2(_08724_),
    .A3(_08728_),
    .B1(_11713_),
    .Y(_08730_));
 sky130_fd_sc_hd__a22o_2 _21941_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[3][11] ),
    .B1(_08729_),
    .B2(_08730_),
    .X(_01757_));
 sky130_fd_sc_hd__a31o_2 _21942_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[10] ),
    .A2(\systolic_inst.acc_wires[3][10] ),
    .A3(_08725_),
    .B1(_08727_),
    .X(_08731_));
 sky130_fd_sc_hd__and3_2 _21943_ (.A(_08720_),
    .B(_08725_),
    .C(_08726_),
    .X(_08732_));
 sky130_fd_sc_hd__and2_2 _21944_ (.A(_08721_),
    .B(_08732_),
    .X(_08733_));
 sky130_fd_sc_hd__or4b_2 _21945_ (.A(_08710_),
    .B(_08713_),
    .C(_08714_),
    .D_N(_08732_),
    .X(_08734_));
 sky130_fd_sc_hd__a21oi_2 _21946_ (.A1(_08706_),
    .A2(_08709_),
    .B1(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__or2_2 _21947_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[3][12] ),
    .X(_08736_));
 sky130_fd_sc_hd__nand2_2 _21948_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[3][12] ),
    .Y(_08737_));
 sky130_fd_sc_hd__and2_2 _21949_ (.A(_08736_),
    .B(_08737_),
    .X(_08738_));
 sky130_fd_sc_hd__or4_2 _21950_ (.A(_08731_),
    .B(_08733_),
    .C(_08735_),
    .D(_08738_),
    .X(_08739_));
 sky130_fd_sc_hd__o31ai_2 _21951_ (.A1(_08731_),
    .A2(_08733_),
    .A3(_08735_),
    .B1(_08738_),
    .Y(_08740_));
 sky130_fd_sc_hd__a32o_2 _21952_ (.A1(_11712_),
    .A2(_08739_),
    .A3(_08740_),
    .B1(\systolic_inst.acc_wires[3][12] ),
    .B2(_11258_),
    .X(_01758_));
 sky130_fd_sc_hd__or2_2 _21953_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[3][13] ),
    .X(_08741_));
 sky130_fd_sc_hd__nand2_2 _21954_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[3][13] ),
    .Y(_08742_));
 sky130_fd_sc_hd__inv_2 _21955_ (.A(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__nand2_2 _21956_ (.A(_08741_),
    .B(_08742_),
    .Y(_08744_));
 sky130_fd_sc_hd__nand3_2 _21957_ (.A(_08737_),
    .B(_08740_),
    .C(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__a21o_2 _21958_ (.A1(_08737_),
    .A2(_08740_),
    .B1(_08744_),
    .X(_08746_));
 sky130_fd_sc_hd__a32o_2 _21959_ (.A1(_11712_),
    .A2(_08745_),
    .A3(_08746_),
    .B1(\systolic_inst.acc_wires[3][13] ),
    .B2(_11258_),
    .X(_01759_));
 sky130_fd_sc_hd__or2_2 _21960_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[3][14] ),
    .X(_08747_));
 sky130_fd_sc_hd__nand2_2 _21961_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[3][14] ),
    .Y(_08748_));
 sky130_fd_sc_hd__nand2_2 _21962_ (.A(_08747_),
    .B(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand3_2 _21963_ (.A(_08742_),
    .B(_08746_),
    .C(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__a21o_2 _21964_ (.A1(_08742_),
    .A2(_08746_),
    .B1(_08749_),
    .X(_08751_));
 sky130_fd_sc_hd__a32o_2 _21965_ (.A1(_11712_),
    .A2(_08750_),
    .A3(_08751_),
    .B1(\systolic_inst.acc_wires[3][14] ),
    .B2(_11258_),
    .X(_01760_));
 sky130_fd_sc_hd__or2_2 _21966_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][15] ),
    .X(_08752_));
 sky130_fd_sc_hd__nand2_2 _21967_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][15] ),
    .Y(_08753_));
 sky130_fd_sc_hd__nand2_2 _21968_ (.A(_08752_),
    .B(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__a21oi_2 _21969_ (.A1(_08748_),
    .A2(_08751_),
    .B1(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__a31o_2 _21970_ (.A1(_08748_),
    .A2(_08751_),
    .A3(_08754_),
    .B1(_11713_),
    .X(_08756_));
 sky130_fd_sc_hd__a2bb2o_2 _21971_ (.A1_N(_08756_),
    .A2_N(_08755_),
    .B1(\systolic_inst.acc_wires[3][15] ),
    .B2(_11258_),
    .X(_01761_));
 sky130_fd_sc_hd__nor2_2 _21972_ (.A(_08749_),
    .B(_08754_),
    .Y(_08757_));
 sky130_fd_sc_hd__and3_2 _21973_ (.A(_08741_),
    .B(_08742_),
    .C(_08757_),
    .X(_08758_));
 sky130_fd_sc_hd__o311a_2 _21974_ (.A1(_08731_),
    .A2(_08733_),
    .A3(_08735_),
    .B1(_08738_),
    .C1(_08758_),
    .X(_08759_));
 sky130_fd_sc_hd__a31o_2 _21975_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[3][12] ),
    .A3(_08741_),
    .B1(_08743_),
    .X(_08760_));
 sky130_fd_sc_hd__and3_2 _21976_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[3][14] ),
    .C(_08752_),
    .X(_08761_));
 sky130_fd_sc_hd__a221oi_2 _21977_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[3][15] ),
    .B1(_08757_),
    .B2(_08760_),
    .C1(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__inv_2 _21978_ (.A(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__or2_2 _21979_ (.A(_08759_),
    .B(_08763_),
    .X(_08764_));
 sky130_fd_sc_hd__xnor2_2 _21980_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][16] ),
    .Y(_08765_));
 sky130_fd_sc_hd__and2b_2 _21981_ (.A_N(_08765_),
    .B(_08764_),
    .X(_08766_));
 sky130_fd_sc_hd__xnor2_2 _21982_ (.A(_08764_),
    .B(_08765_),
    .Y(_08767_));
 sky130_fd_sc_hd__a22o_2 _21983_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[3][16] ),
    .B1(_11712_),
    .B2(_08767_),
    .X(_01762_));
 sky130_fd_sc_hd__xor2_2 _21984_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][17] ),
    .X(_08768_));
 sky130_fd_sc_hd__inv_2 _21985_ (.A(_08768_),
    .Y(_08769_));
 sky130_fd_sc_hd__a21oi_2 _21986_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[3][16] ),
    .B1(_08766_),
    .Y(_08770_));
 sky130_fd_sc_hd__xnor2_2 _21987_ (.A(_08768_),
    .B(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__a22o_2 _21988_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[3][17] ),
    .B1(_11712_),
    .B2(_08771_),
    .X(_01763_));
 sky130_fd_sc_hd__or2_2 _21989_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][18] ),
    .X(_08772_));
 sky130_fd_sc_hd__nand2_2 _21990_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][18] ),
    .Y(_08773_));
 sky130_fd_sc_hd__nand2_2 _21991_ (.A(_08772_),
    .B(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__o21ai_2 _21992_ (.A1(\systolic_inst.acc_wires[3][16] ),
    .A2(\systolic_inst.acc_wires[3][17] ),
    .B1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .Y(_08775_));
 sky130_fd_sc_hd__nand2_2 _21993_ (.A(_08766_),
    .B(_08768_),
    .Y(_08776_));
 sky130_fd_sc_hd__a21o_2 _21994_ (.A1(_08775_),
    .A2(_08776_),
    .B1(_08774_),
    .X(_08777_));
 sky130_fd_sc_hd__nand3_2 _21995_ (.A(_08774_),
    .B(_08775_),
    .C(_08776_),
    .Y(_08778_));
 sky130_fd_sc_hd__a32o_2 _21996_ (.A1(_11712_),
    .A2(_08777_),
    .A3(_08778_),
    .B1(\systolic_inst.acc_wires[3][18] ),
    .B2(_11258_),
    .X(_01764_));
 sky130_fd_sc_hd__xnor2_2 _21997_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][19] ),
    .Y(_08779_));
 sky130_fd_sc_hd__a21oi_2 _21998_ (.A1(_08773_),
    .A2(_08777_),
    .B1(_08779_),
    .Y(_08780_));
 sky130_fd_sc_hd__a31o_2 _21999_ (.A1(_08773_),
    .A2(_08777_),
    .A3(_08779_),
    .B1(_11713_),
    .X(_08781_));
 sky130_fd_sc_hd__a2bb2o_2 _22000_ (.A1_N(_08781_),
    .A2_N(_08780_),
    .B1(\systolic_inst.acc_wires[3][19] ),
    .B2(_11258_),
    .X(_01765_));
 sky130_fd_sc_hd__or2_2 _22001_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][20] ),
    .X(_08782_));
 sky130_fd_sc_hd__nand2_2 _22002_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][20] ),
    .Y(_08783_));
 sky130_fd_sc_hd__and2_2 _22003_ (.A(_08782_),
    .B(_08783_),
    .X(_08784_));
 sky130_fd_sc_hd__or4_2 _22004_ (.A(_08765_),
    .B(_08769_),
    .C(_08774_),
    .D(_08779_),
    .X(_08785_));
 sky130_fd_sc_hd__o21ba_2 _22005_ (.A1(_08759_),
    .A2(_08763_),
    .B1_N(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__o41a_2 _22006_ (.A1(\systolic_inst.acc_wires[3][16] ),
    .A2(\systolic_inst.acc_wires[3][17] ),
    .A3(\systolic_inst.acc_wires[3][18] ),
    .A4(\systolic_inst.acc_wires[3][19] ),
    .B1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .X(_08787_));
 sky130_fd_sc_hd__or3_2 _22007_ (.A(_08784_),
    .B(_08786_),
    .C(_08787_),
    .X(_08788_));
 sky130_fd_sc_hd__o21ai_2 _22008_ (.A1(_08786_),
    .A2(_08787_),
    .B1(_08784_),
    .Y(_08789_));
 sky130_fd_sc_hd__a32o_2 _22009_ (.A1(_11712_),
    .A2(_08788_),
    .A3(_08789_),
    .B1(\systolic_inst.acc_wires[3][20] ),
    .B2(_11258_),
    .X(_01766_));
 sky130_fd_sc_hd__xnor2_2 _22010_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][21] ),
    .Y(_08790_));
 sky130_fd_sc_hd__inv_2 _22011_ (.A(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__a21oi_2 _22012_ (.A1(_08783_),
    .A2(_08789_),
    .B1(_08790_),
    .Y(_08792_));
 sky130_fd_sc_hd__a31o_2 _22013_ (.A1(_08783_),
    .A2(_08789_),
    .A3(_08790_),
    .B1(_11713_),
    .X(_08793_));
 sky130_fd_sc_hd__a2bb2o_2 _22014_ (.A1_N(_08793_),
    .A2_N(_08792_),
    .B1(\systolic_inst.acc_wires[3][21] ),
    .B2(_11258_),
    .X(_01767_));
 sky130_fd_sc_hd__nor2_2 _22015_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][22] ),
    .Y(_08794_));
 sky130_fd_sc_hd__and2_2 _22016_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][22] ),
    .X(_08795_));
 sky130_fd_sc_hd__nor2_2 _22017_ (.A(_08794_),
    .B(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__o21a_2 _22018_ (.A1(\systolic_inst.acc_wires[3][20] ),
    .A2(\systolic_inst.acc_wires[3][21] ),
    .B1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .X(_08797_));
 sky130_fd_sc_hd__o21bai_2 _22019_ (.A1(_08789_),
    .A2(_08790_),
    .B1_N(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__xor2_2 _22020_ (.A(_08796_),
    .B(_08798_),
    .X(_08799_));
 sky130_fd_sc_hd__a22o_2 _22021_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[3][22] ),
    .B1(_11712_),
    .B2(_08799_),
    .X(_01768_));
 sky130_fd_sc_hd__xor2_2 _22022_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][23] ),
    .X(_08800_));
 sky130_fd_sc_hd__a21o_2 _22023_ (.A1(_08796_),
    .A2(_08798_),
    .B1(_08795_),
    .X(_08801_));
 sky130_fd_sc_hd__xor2_2 _22024_ (.A(_08800_),
    .B(_08801_),
    .X(_08802_));
 sky130_fd_sc_hd__a22o_2 _22025_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[3][23] ),
    .B1(_11712_),
    .B2(_08802_),
    .X(_01769_));
 sky130_fd_sc_hd__and4_2 _22026_ (.A(_08784_),
    .B(_08791_),
    .C(_08796_),
    .D(_08800_),
    .X(_08803_));
 sky130_fd_sc_hd__a2111o_2 _22027_ (.A1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[3][23] ),
    .B1(_08787_),
    .C1(_08795_),
    .D1(_08797_),
    .X(_08804_));
 sky130_fd_sc_hd__a21oi_2 _22028_ (.A1(_08786_),
    .A2(_08803_),
    .B1(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__nor2_2 _22029_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][24] ),
    .Y(_08806_));
 sky130_fd_sc_hd__and2_2 _22030_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][24] ),
    .X(_08807_));
 sky130_fd_sc_hd__or2_2 _22031_ (.A(_08806_),
    .B(_08807_),
    .X(_08808_));
 sky130_fd_sc_hd__nor2_2 _22032_ (.A(_08805_),
    .B(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__a21o_2 _22033_ (.A1(_08805_),
    .A2(_08808_),
    .B1(_11713_),
    .X(_08810_));
 sky130_fd_sc_hd__a2bb2o_2 _22034_ (.A1_N(_08810_),
    .A2_N(_08809_),
    .B1(\systolic_inst.acc_wires[3][24] ),
    .B2(_11258_),
    .X(_01770_));
 sky130_fd_sc_hd__xor2_2 _22035_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][25] ),
    .X(_08811_));
 sky130_fd_sc_hd__or3_2 _22036_ (.A(_08807_),
    .B(_08809_),
    .C(_08811_),
    .X(_08812_));
 sky130_fd_sc_hd__o21ai_2 _22037_ (.A1(_08807_),
    .A2(_08809_),
    .B1(_08811_),
    .Y(_08813_));
 sky130_fd_sc_hd__a32o_2 _22038_ (.A1(_11712_),
    .A2(_08812_),
    .A3(_08813_),
    .B1(\systolic_inst.acc_wires[3][25] ),
    .B2(_11258_),
    .X(_01771_));
 sky130_fd_sc_hd__or2_2 _22039_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][26] ),
    .X(_08814_));
 sky130_fd_sc_hd__nand2_2 _22040_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][26] ),
    .Y(_08815_));
 sky130_fd_sc_hd__and2_2 _22041_ (.A(_08814_),
    .B(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__o21a_2 _22042_ (.A1(\systolic_inst.acc_wires[3][24] ),
    .A2(\systolic_inst.acc_wires[3][25] ),
    .B1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .X(_08817_));
 sky130_fd_sc_hd__and2_2 _22043_ (.A(_08809_),
    .B(_08811_),
    .X(_08818_));
 sky130_fd_sc_hd__o21ai_2 _22044_ (.A1(_08817_),
    .A2(_08818_),
    .B1(_08816_),
    .Y(_08819_));
 sky130_fd_sc_hd__or3_2 _22045_ (.A(_08816_),
    .B(_08817_),
    .C(_08818_),
    .X(_08820_));
 sky130_fd_sc_hd__a32o_2 _22046_ (.A1(_11712_),
    .A2(_08819_),
    .A3(_08820_),
    .B1(\systolic_inst.acc_wires[3][26] ),
    .B2(_11258_),
    .X(_01772_));
 sky130_fd_sc_hd__xnor2_2 _22047_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][27] ),
    .Y(_08821_));
 sky130_fd_sc_hd__a21oi_2 _22048_ (.A1(_08815_),
    .A2(_08819_),
    .B1(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__a31o_2 _22049_ (.A1(_08815_),
    .A2(_08819_),
    .A3(_08821_),
    .B1(_11713_),
    .X(_08823_));
 sky130_fd_sc_hd__a2bb2o_2 _22050_ (.A1_N(_08823_),
    .A2_N(_08822_),
    .B1(\systolic_inst.acc_wires[3][27] ),
    .B2(_11258_),
    .X(_01773_));
 sky130_fd_sc_hd__nand2_2 _22051_ (.A(_08811_),
    .B(_08816_),
    .Y(_08824_));
 sky130_fd_sc_hd__or4_2 _22052_ (.A(_08805_),
    .B(_08808_),
    .C(_08821_),
    .D(_08824_),
    .X(_08825_));
 sky130_fd_sc_hd__o21a_2 _22053_ (.A1(\systolic_inst.acc_wires[3][26] ),
    .A2(\systolic_inst.acc_wires[3][27] ),
    .B1(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .X(_08826_));
 sky130_fd_sc_hd__nor2_2 _22054_ (.A(_08817_),
    .B(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__nor2_2 _22055_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][28] ),
    .Y(_08828_));
 sky130_fd_sc_hd__and2_2 _22056_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][28] ),
    .X(_08829_));
 sky130_fd_sc_hd__or2_2 _22057_ (.A(_08828_),
    .B(_08829_),
    .X(_08830_));
 sky130_fd_sc_hd__and3_2 _22058_ (.A(_08825_),
    .B(_08827_),
    .C(_08830_),
    .X(_08831_));
 sky130_fd_sc_hd__a21oi_2 _22059_ (.A1(_08825_),
    .A2(_08827_),
    .B1(_08830_),
    .Y(_08832_));
 sky130_fd_sc_hd__or2_2 _22060_ (.A(_08831_),
    .B(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__a2bb2o_2 _22061_ (.A1_N(_11713_),
    .A2_N(_08833_),
    .B1(_11258_),
    .B2(\systolic_inst.acc_wires[3][28] ),
    .X(_01774_));
 sky130_fd_sc_hd__nor2_2 _22062_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][29] ),
    .Y(_08834_));
 sky130_fd_sc_hd__and2_2 _22063_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][29] ),
    .X(_08835_));
 sky130_fd_sc_hd__nor2_2 _22064_ (.A(_08834_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__o21ai_2 _22065_ (.A1(_08829_),
    .A2(_08832_),
    .B1(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__or3_2 _22066_ (.A(_08829_),
    .B(_08832_),
    .C(_08836_),
    .X(_08838_));
 sky130_fd_sc_hd__a32o_2 _22067_ (.A1(_11712_),
    .A2(_08837_),
    .A3(_08838_),
    .B1(\systolic_inst.acc_wires[3][29] ),
    .B2(_11258_),
    .X(_01775_));
 sky130_fd_sc_hd__and2_2 _22068_ (.A(_08832_),
    .B(_08836_),
    .X(_08839_));
 sky130_fd_sc_hd__nand2_2 _22069_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][30] ),
    .Y(_08840_));
 sky130_fd_sc_hd__or2_2 _22070_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][30] ),
    .X(_08841_));
 sky130_fd_sc_hd__a2111o_2 _22071_ (.A1(_08840_),
    .A2(_08841_),
    .B1(_08829_),
    .C1(_08835_),
    .D1(_08839_),
    .X(_08842_));
 sky130_fd_sc_hd__o311ai_2 _22072_ (.A1(_08829_),
    .A2(_08835_),
    .A3(_08839_),
    .B1(_08840_),
    .C1(_08841_),
    .Y(_08843_));
 sky130_fd_sc_hd__a32o_2 _22073_ (.A1(_11712_),
    .A2(_08842_),
    .A3(_08843_),
    .B1(\systolic_inst.acc_wires[3][30] ),
    .B2(_11258_),
    .X(_01776_));
 sky130_fd_sc_hd__xnor2_2 _22074_ (.A(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[3][31] ),
    .Y(_08844_));
 sky130_fd_sc_hd__a21oi_2 _22075_ (.A1(_08840_),
    .A2(_08843_),
    .B1(_08844_),
    .Y(_08845_));
 sky130_fd_sc_hd__a31o_2 _22076_ (.A1(_08840_),
    .A2(_08843_),
    .A3(_08844_),
    .B1(_11713_),
    .X(_08846_));
 sky130_fd_sc_hd__a2bb2o_2 _22077_ (.A1_N(_08846_),
    .A2_N(_08845_),
    .B1(\systolic_inst.acc_wires[3][31] ),
    .B2(_11258_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _22078_ (.A0(\systolic_inst.A_outs[2][0] ),
    .A1(\systolic_inst.A_outs[1][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _22079_ (.A0(\systolic_inst.A_outs[2][1] ),
    .A1(\systolic_inst.A_outs[1][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _22080_ (.A0(\systolic_inst.A_outs[2][2] ),
    .A1(\systolic_inst.A_outs[1][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _22081_ (.A0(\systolic_inst.A_outs[2][3] ),
    .A1(\systolic_inst.A_outs[1][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _22082_ (.A0(\systolic_inst.A_outs[2][4] ),
    .A1(\systolic_inst.A_outs[1][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _22083_ (.A0(\systolic_inst.A_outs[2][5] ),
    .A1(\systolic_inst.A_outs[1][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _22084_ (.A0(\systolic_inst.A_outs[2][6] ),
    .A1(\systolic_inst.A_outs[1][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _22085_ (.A0(\systolic_inst.A_outs[2][7] ),
    .A1(\systolic_inst.A_outs[1][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _22086_ (.A0(\systolic_inst.B_outs[1][0] ),
    .A1(\systolic_inst.B_shift[1][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _22087_ (.A0(\systolic_inst.B_outs[1][1] ),
    .A1(\systolic_inst.B_shift[1][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _22088_ (.A0(\systolic_inst.B_outs[1][2] ),
    .A1(\systolic_inst.B_shift[1][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _22089_ (.A0(\systolic_inst.B_outs[1][3] ),
    .A1(\systolic_inst.B_shift[1][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _22090_ (.A0(\systolic_inst.B_outs[1][4] ),
    .A1(\systolic_inst.B_shift[1][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _22091_ (.A0(\systolic_inst.B_outs[1][5] ),
    .A1(\systolic_inst.B_shift[1][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _22092_ (.A0(\systolic_inst.B_outs[1][6] ),
    .A1(\systolic_inst.B_shift[1][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _22093_ (.A0(\systolic_inst.B_outs[1][7] ),
    .A1(\systolic_inst.B_shift[1][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01793_));
 sky130_fd_sc_hd__and3_2 _22094_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[2][0] ),
    .C(\systolic_inst.A_outs[2][0] ),
    .X(_08847_));
 sky130_fd_sc_hd__a21o_2 _22095_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[0] ),
    .B1(_08847_),
    .X(_01794_));
 sky130_fd_sc_hd__and4_2 _22096_ (.A(\systolic_inst.B_outs[2][0] ),
    .B(\systolic_inst.A_outs[2][0] ),
    .C(\systolic_inst.B_outs[2][1] ),
    .D(\systolic_inst.A_outs[2][1] ),
    .X(_08848_));
 sky130_fd_sc_hd__a22o_2 _22097_ (.A1(\systolic_inst.A_outs[2][0] ),
    .A2(\systolic_inst.B_outs[2][1] ),
    .B1(\systolic_inst.A_outs[2][1] ),
    .B2(\systolic_inst.B_outs[2][0] ),
    .X(_08849_));
 sky130_fd_sc_hd__nand2_2 _22098_ (.A(\systolic_inst.ce_local ),
    .B(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__a2bb2o_2 _22099_ (.A1_N(_08850_),
    .A2_N(_08848_),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01795_));
 sky130_fd_sc_hd__and2_2 _22100_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[2] ),
    .X(_08851_));
 sky130_fd_sc_hd__a22oi_2 _22101_ (.A1(\systolic_inst.B_outs[2][1] ),
    .A2(\systolic_inst.A_outs[2][1] ),
    .B1(\systolic_inst.A_outs[2][2] ),
    .B2(\systolic_inst.B_outs[2][0] ),
    .Y(_08852_));
 sky130_fd_sc_hd__and4_2 _22102_ (.A(\systolic_inst.B_outs[2][0] ),
    .B(\systolic_inst.B_outs[2][1] ),
    .C(\systolic_inst.A_outs[2][1] ),
    .D(\systolic_inst.A_outs[2][2] ),
    .X(_08853_));
 sky130_fd_sc_hd__or2_2 _22103_ (.A(_08852_),
    .B(_08853_),
    .X(_08854_));
 sky130_fd_sc_hd__or3b_2 _22104_ (.A(_08852_),
    .B(_08853_),
    .C_N(_08848_),
    .X(_08855_));
 sky130_fd_sc_hd__xnor2_2 _22105_ (.A(_08848_),
    .B(_08854_),
    .Y(_08856_));
 sky130_fd_sc_hd__nand3_2 _22106_ (.A(\systolic_inst.A_outs[2][0] ),
    .B(\systolic_inst.B_outs[2][2] ),
    .C(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__a21o_2 _22107_ (.A1(\systolic_inst.A_outs[2][0] ),
    .A2(\systolic_inst.B_outs[2][2] ),
    .B1(_08856_),
    .X(_08858_));
 sky130_fd_sc_hd__a31o_2 _22108_ (.A1(\systolic_inst.ce_local ),
    .A2(_08857_),
    .A3(_08858_),
    .B1(_08851_),
    .X(_01796_));
 sky130_fd_sc_hd__a22oi_2 _22109_ (.A1(\systolic_inst.A_outs[2][1] ),
    .A2(\systolic_inst.B_outs[2][2] ),
    .B1(\systolic_inst.B_outs[2][3] ),
    .B2(\systolic_inst.A_outs[2][0] ),
    .Y(_08859_));
 sky130_fd_sc_hd__and4_2 _22110_ (.A(\systolic_inst.A_outs[2][0] ),
    .B(\systolic_inst.A_outs[2][1] ),
    .C(\systolic_inst.B_outs[2][2] ),
    .D(\systolic_inst.B_outs[2][3] ),
    .X(_08860_));
 sky130_fd_sc_hd__nor2_2 _22111_ (.A(_08859_),
    .B(_08860_),
    .Y(_08861_));
 sky130_fd_sc_hd__nand4_2 _22112_ (.A(\systolic_inst.B_outs[2][0] ),
    .B(\systolic_inst.B_outs[2][1] ),
    .C(\systolic_inst.A_outs[2][2] ),
    .D(\systolic_inst.A_outs[2][3] ),
    .Y(_08862_));
 sky130_fd_sc_hd__a22o_2 _22113_ (.A1(\systolic_inst.B_outs[2][1] ),
    .A2(\systolic_inst.A_outs[2][2] ),
    .B1(\systolic_inst.A_outs[2][3] ),
    .B2(\systolic_inst.B_outs[2][0] ),
    .X(_08863_));
 sky130_fd_sc_hd__nand3_2 _22114_ (.A(_08853_),
    .B(_08862_),
    .C(_08863_),
    .Y(_08864_));
 sky130_fd_sc_hd__a21o_2 _22115_ (.A1(_08862_),
    .A2(_08863_),
    .B1(_08853_),
    .X(_08865_));
 sky130_fd_sc_hd__and2_2 _22116_ (.A(_08864_),
    .B(_08865_),
    .X(_08866_));
 sky130_fd_sc_hd__nand2_2 _22117_ (.A(_08861_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__xnor2_2 _22118_ (.A(_08861_),
    .B(_08866_),
    .Y(_08868_));
 sky130_fd_sc_hd__and3_2 _22119_ (.A(_08855_),
    .B(_08857_),
    .C(_08868_),
    .X(_08869_));
 sky130_fd_sc_hd__a21oi_2 _22120_ (.A1(_08855_),
    .A2(_08857_),
    .B1(_08868_),
    .Y(_08870_));
 sky130_fd_sc_hd__nand2_2 _22121_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[3] ),
    .Y(_08871_));
 sky130_fd_sc_hd__o31ai_2 _22122_ (.A1(_11258_),
    .A2(_08869_),
    .A3(_08870_),
    .B1(_08871_),
    .Y(_01797_));
 sky130_fd_sc_hd__and2_2 _22123_ (.A(\systolic_inst.B_outs[2][2] ),
    .B(\systolic_inst.A_outs[2][2] ),
    .X(_08872_));
 sky130_fd_sc_hd__nand4_2 _22124_ (.A(\systolic_inst.A_outs[2][0] ),
    .B(\systolic_inst.A_outs[2][1] ),
    .C(\systolic_inst.B_outs[2][3] ),
    .D(\systolic_inst.B_outs[2][4] ),
    .Y(_08873_));
 sky130_fd_sc_hd__a22o_2 _22125_ (.A1(\systolic_inst.A_outs[2][1] ),
    .A2(\systolic_inst.B_outs[2][3] ),
    .B1(\systolic_inst.B_outs[2][4] ),
    .B2(\systolic_inst.A_outs[2][0] ),
    .X(_08874_));
 sky130_fd_sc_hd__nand2_2 _22126_ (.A(_08873_),
    .B(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__xnor2_2 _22127_ (.A(_08872_),
    .B(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__a22o_2 _22128_ (.A1(\systolic_inst.B_outs[2][1] ),
    .A2(\systolic_inst.A_outs[2][3] ),
    .B1(\systolic_inst.A_outs[2][4] ),
    .B2(\systolic_inst.B_outs[2][0] ),
    .X(_08877_));
 sky130_fd_sc_hd__and3_2 _22129_ (.A(\systolic_inst.B_outs[2][0] ),
    .B(\systolic_inst.B_outs[2][1] ),
    .C(\systolic_inst.A_outs[2][3] ),
    .X(_08878_));
 sky130_fd_sc_hd__nand2_2 _22130_ (.A(\systolic_inst.A_outs[2][4] ),
    .B(_08878_),
    .Y(_08879_));
 sky130_fd_sc_hd__and3_2 _22131_ (.A(_08860_),
    .B(_08877_),
    .C(_08879_),
    .X(_08880_));
 sky130_fd_sc_hd__a21oi_2 _22132_ (.A1(_08877_),
    .A2(_08879_),
    .B1(_08860_),
    .Y(_08881_));
 sky130_fd_sc_hd__o21ai_2 _22133_ (.A1(_08880_),
    .A2(_08881_),
    .B1(_08862_),
    .Y(_08882_));
 sky130_fd_sc_hd__or3_2 _22134_ (.A(_08862_),
    .B(_08880_),
    .C(_08881_),
    .X(_08883_));
 sky130_fd_sc_hd__and3_2 _22135_ (.A(_08876_),
    .B(_08882_),
    .C(_08883_),
    .X(_08884_));
 sky130_fd_sc_hd__a21oi_2 _22136_ (.A1(_08882_),
    .A2(_08883_),
    .B1(_08876_),
    .Y(_08885_));
 sky130_fd_sc_hd__a211o_2 _22137_ (.A1(_08864_),
    .A2(_08867_),
    .B1(_08884_),
    .C1(_08885_),
    .X(_08886_));
 sky130_fd_sc_hd__o211ai_2 _22138_ (.A1(_08884_),
    .A2(_08885_),
    .B1(_08864_),
    .C1(_08867_),
    .Y(_08887_));
 sky130_fd_sc_hd__a21oi_2 _22139_ (.A1(_08886_),
    .A2(_08887_),
    .B1(_08870_),
    .Y(_08888_));
 sky130_fd_sc_hd__and3_2 _22140_ (.A(_08870_),
    .B(_08886_),
    .C(_08887_),
    .X(_08889_));
 sky130_fd_sc_hd__or3_2 _22141_ (.A(_11258_),
    .B(_08888_),
    .C(_08889_),
    .X(_08890_));
 sky130_fd_sc_hd__a21bo_2 _22142_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[4] ),
    .B1_N(_08890_),
    .X(_01798_));
 sky130_fd_sc_hd__and2b_2 _22143_ (.A_N(_08880_),
    .B(_08883_),
    .X(_08891_));
 sky130_fd_sc_hd__a21bo_2 _22144_ (.A1(_08872_),
    .A2(_08874_),
    .B1_N(_08873_),
    .X(_08892_));
 sky130_fd_sc_hd__a22oi_2 _22145_ (.A1(\systolic_inst.B_outs[2][1] ),
    .A2(\systolic_inst.A_outs[2][4] ),
    .B1(\systolic_inst.A_outs[2][5] ),
    .B2(\systolic_inst.B_outs[2][0] ),
    .Y(_08893_));
 sky130_fd_sc_hd__and4_2 _22146_ (.A(\systolic_inst.B_outs[2][0] ),
    .B(\systolic_inst.B_outs[2][1] ),
    .C(\systolic_inst.A_outs[2][4] ),
    .D(\systolic_inst.A_outs[2][5] ),
    .X(_08894_));
 sky130_fd_sc_hd__nor2_2 _22147_ (.A(_08893_),
    .B(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__xor2_2 _22148_ (.A(_08892_),
    .B(_08895_),
    .X(_08896_));
 sky130_fd_sc_hd__xor2_2 _22149_ (.A(_08879_),
    .B(_08896_),
    .X(_08897_));
 sky130_fd_sc_hd__and4_2 _22150_ (.A(\systolic_inst.A_outs[2][1] ),
    .B(\systolic_inst.A_outs[2][2] ),
    .C(\systolic_inst.B_outs[2][3] ),
    .D(\systolic_inst.B_outs[2][4] ),
    .X(_08898_));
 sky130_fd_sc_hd__a22oi_2 _22151_ (.A1(\systolic_inst.A_outs[2][2] ),
    .A2(\systolic_inst.B_outs[2][3] ),
    .B1(\systolic_inst.B_outs[2][4] ),
    .B2(\systolic_inst.A_outs[2][1] ),
    .Y(_08899_));
 sky130_fd_sc_hd__a22o_2 _22152_ (.A1(\systolic_inst.A_outs[2][2] ),
    .A2(\systolic_inst.B_outs[2][3] ),
    .B1(\systolic_inst.B_outs[2][4] ),
    .B2(\systolic_inst.A_outs[2][1] ),
    .X(_08900_));
 sky130_fd_sc_hd__and4b_2 _22153_ (.A_N(_08898_),
    .B(_08900_),
    .C(\systolic_inst.B_outs[2][2] ),
    .D(\systolic_inst.A_outs[2][3] ),
    .X(_08901_));
 sky130_fd_sc_hd__o2bb2a_2 _22154_ (.A1_N(\systolic_inst.B_outs[2][2] ),
    .A2_N(\systolic_inst.A_outs[2][3] ),
    .B1(_08898_),
    .B2(_08899_),
    .X(_08902_));
 sky130_fd_sc_hd__and4bb_2 _22155_ (.A_N(_08901_),
    .B_N(_08902_),
    .C(\systolic_inst.A_outs[2][0] ),
    .D(\systolic_inst.B_outs[2][5] ),
    .X(_08903_));
 sky130_fd_sc_hd__o2bb2a_2 _22156_ (.A1_N(\systolic_inst.A_outs[2][0] ),
    .A2_N(\systolic_inst.B_outs[2][5] ),
    .B1(_08901_),
    .B2(_08902_),
    .X(_08904_));
 sky130_fd_sc_hd__or2_2 _22157_ (.A(_08903_),
    .B(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__nor2_2 _22158_ (.A(_08897_),
    .B(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__xor2_2 _22159_ (.A(_08897_),
    .B(_08905_),
    .X(_08907_));
 sky130_fd_sc_hd__nand2_2 _22160_ (.A(_08884_),
    .B(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__xor2_2 _22161_ (.A(_08884_),
    .B(_08907_),
    .X(_08909_));
 sky130_fd_sc_hd__nand2b_2 _22162_ (.A_N(_08891_),
    .B(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__xnor2_2 _22163_ (.A(_08891_),
    .B(_08909_),
    .Y(_08911_));
 sky130_fd_sc_hd__a21bo_2 _22164_ (.A1(_08870_),
    .A2(_08887_),
    .B1_N(_08886_),
    .X(_08912_));
 sky130_fd_sc_hd__nand2_2 _22165_ (.A(_08911_),
    .B(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__o21a_2 _22166_ (.A1(_08911_),
    .A2(_08912_),
    .B1(\systolic_inst.ce_local ),
    .X(_08914_));
 sky130_fd_sc_hd__a22o_2 _22167_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[5] ),
    .B1(_08913_),
    .B2(_08914_),
    .X(_01799_));
 sky130_fd_sc_hd__a32o_2 _22168_ (.A1(\systolic_inst.A_outs[2][4] ),
    .A2(_08878_),
    .A3(_08896_),
    .B1(_08895_),
    .B2(_08892_),
    .X(_08915_));
 sky130_fd_sc_hd__a31o_2 _22169_ (.A1(\systolic_inst.B_outs[2][2] ),
    .A2(\systolic_inst.A_outs[2][3] ),
    .A3(_08900_),
    .B1(_08898_),
    .X(_08916_));
 sky130_fd_sc_hd__a22oi_2 _22170_ (.A1(\systolic_inst.B_outs[2][1] ),
    .A2(\systolic_inst.A_outs[2][5] ),
    .B1(\systolic_inst.A_outs[2][6] ),
    .B2(\systolic_inst.B_outs[2][0] ),
    .Y(_08917_));
 sky130_fd_sc_hd__and4_2 _22171_ (.A(\systolic_inst.B_outs[2][0] ),
    .B(\systolic_inst.B_outs[2][1] ),
    .C(\systolic_inst.A_outs[2][5] ),
    .D(\systolic_inst.A_outs[2][6] ),
    .X(_08918_));
 sky130_fd_sc_hd__or2_2 _22172_ (.A(_08917_),
    .B(_08918_),
    .X(_08919_));
 sky130_fd_sc_hd__and2b_2 _22173_ (.A_N(_08919_),
    .B(_08916_),
    .X(_08920_));
 sky130_fd_sc_hd__xnor2_2 _22174_ (.A(_08916_),
    .B(_08919_),
    .Y(_08921_));
 sky130_fd_sc_hd__xor2_2 _22175_ (.A(_08894_),
    .B(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__nand4_2 _22176_ (.A(\systolic_inst.A_outs[2][2] ),
    .B(\systolic_inst.B_outs[2][3] ),
    .C(\systolic_inst.A_outs[2][3] ),
    .D(\systolic_inst.B_outs[2][4] ),
    .Y(_08923_));
 sky130_fd_sc_hd__a22o_2 _22177_ (.A1(\systolic_inst.B_outs[2][3] ),
    .A2(\systolic_inst.A_outs[2][3] ),
    .B1(\systolic_inst.B_outs[2][4] ),
    .B2(\systolic_inst.A_outs[2][2] ),
    .X(_08924_));
 sky130_fd_sc_hd__nand4_2 _22178_ (.A(\systolic_inst.B_outs[2][2] ),
    .B(\systolic_inst.A_outs[2][4] ),
    .C(_08923_),
    .D(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__a22o_2 _22179_ (.A1(\systolic_inst.B_outs[2][2] ),
    .A2(\systolic_inst.A_outs[2][4] ),
    .B1(_08923_),
    .B2(_08924_),
    .X(_08926_));
 sky130_fd_sc_hd__a22oi_2 _22180_ (.A1(\systolic_inst.A_outs[2][1] ),
    .A2(\systolic_inst.B_outs[2][5] ),
    .B1(\systolic_inst.B_outs[2][6] ),
    .B2(\systolic_inst.A_outs[2][0] ),
    .Y(_08927_));
 sky130_fd_sc_hd__nand2_2 _22181_ (.A(\systolic_inst.A_outs[2][1] ),
    .B(\systolic_inst.B_outs[2][6] ),
    .Y(_08928_));
 sky130_fd_sc_hd__and4_2 _22182_ (.A(\systolic_inst.A_outs[2][0] ),
    .B(\systolic_inst.A_outs[2][1] ),
    .C(\systolic_inst.B_outs[2][5] ),
    .D(\systolic_inst.B_outs[2][6] ),
    .X(_08929_));
 sky130_fd_sc_hd__nor2_2 _22183_ (.A(_08927_),
    .B(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__nand3_2 _22184_ (.A(_08925_),
    .B(_08926_),
    .C(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__a21o_2 _22185_ (.A1(_08925_),
    .A2(_08926_),
    .B1(_08930_),
    .X(_08932_));
 sky130_fd_sc_hd__and3_2 _22186_ (.A(_08903_),
    .B(_08931_),
    .C(_08932_),
    .X(_08933_));
 sky130_fd_sc_hd__a21oi_2 _22187_ (.A1(_08931_),
    .A2(_08932_),
    .B1(_08903_),
    .Y(_08934_));
 sky130_fd_sc_hd__or3b_2 _22188_ (.A(_08933_),
    .B(_08934_),
    .C_N(_08922_),
    .X(_08935_));
 sky130_fd_sc_hd__o21bai_2 _22189_ (.A1(_08933_),
    .A2(_08934_),
    .B1_N(_08922_),
    .Y(_08936_));
 sky130_fd_sc_hd__nand3_2 _22190_ (.A(_08906_),
    .B(_08935_),
    .C(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__a21o_2 _22191_ (.A1(_08935_),
    .A2(_08936_),
    .B1(_08906_),
    .X(_08938_));
 sky130_fd_sc_hd__and3_2 _22192_ (.A(_08915_),
    .B(_08937_),
    .C(_08938_),
    .X(_08939_));
 sky130_fd_sc_hd__a21oi_2 _22193_ (.A1(_08937_),
    .A2(_08938_),
    .B1(_08915_),
    .Y(_08940_));
 sky130_fd_sc_hd__a211oi_2 _22194_ (.A1(_08908_),
    .A2(_08910_),
    .B1(_08939_),
    .C1(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__o211a_2 _22195_ (.A1(_08939_),
    .A2(_08940_),
    .B1(_08908_),
    .C1(_08910_),
    .X(_08942_));
 sky130_fd_sc_hd__nor2_2 _22196_ (.A(_08941_),
    .B(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__xnor2_2 _22197_ (.A(_08913_),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__mux2_1 _22198_ (.A0(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[6] ),
    .A1(_08944_),
    .S(\systolic_inst.ce_local ),
    .X(_01800_));
 sky130_fd_sc_hd__a21boi_2 _22199_ (.A1(_08915_),
    .A2(_08938_),
    .B1_N(_08937_),
    .Y(_08945_));
 sky130_fd_sc_hd__a21oi_2 _22200_ (.A1(_08894_),
    .A2(_08921_),
    .B1(_08920_),
    .Y(_08946_));
 sky130_fd_sc_hd__nand2_2 _22201_ (.A(_08923_),
    .B(_08925_),
    .Y(_08947_));
 sky130_fd_sc_hd__a22o_2 _22202_ (.A1(\systolic_inst.B_outs[2][1] ),
    .A2(\systolic_inst.A_outs[2][6] ),
    .B1(\systolic_inst.A_outs[2][7] ),
    .B2(\systolic_inst.B_outs[2][0] ),
    .X(_08948_));
 sky130_fd_sc_hd__nand4_2 _22203_ (.A(\systolic_inst.B_outs[2][0] ),
    .B(\systolic_inst.B_outs[2][1] ),
    .C(\systolic_inst.A_outs[2][6] ),
    .D(\systolic_inst.A_outs[2][7] ),
    .Y(_08949_));
 sky130_fd_sc_hd__nand2_2 _22204_ (.A(_08948_),
    .B(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__xnor2_2 _22205_ (.A(_11265_),
    .B(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__nand2b_2 _22206_ (.A_N(_08951_),
    .B(_08947_),
    .Y(_08952_));
 sky130_fd_sc_hd__xnor2_2 _22207_ (.A(_08947_),
    .B(_08951_),
    .Y(_08953_));
 sky130_fd_sc_hd__xnor2_2 _22208_ (.A(_08918_),
    .B(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__nand2_2 _22209_ (.A(\systolic_inst.B_outs[2][2] ),
    .B(\systolic_inst.A_outs[2][5] ),
    .Y(_08955_));
 sky130_fd_sc_hd__and4_2 _22210_ (.A(\systolic_inst.B_outs[2][3] ),
    .B(\systolic_inst.A_outs[2][3] ),
    .C(\systolic_inst.B_outs[2][4] ),
    .D(\systolic_inst.A_outs[2][4] ),
    .X(_08956_));
 sky130_fd_sc_hd__a22oi_2 _22211_ (.A1(\systolic_inst.A_outs[2][3] ),
    .A2(\systolic_inst.B_outs[2][4] ),
    .B1(\systolic_inst.A_outs[2][4] ),
    .B2(\systolic_inst.B_outs[2][3] ),
    .Y(_08957_));
 sky130_fd_sc_hd__or2_2 _22212_ (.A(_08956_),
    .B(_08957_),
    .X(_08958_));
 sky130_fd_sc_hd__xnor2_2 _22213_ (.A(_08955_),
    .B(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__nand2_2 _22214_ (.A(\systolic_inst.A_outs[2][2] ),
    .B(\systolic_inst.B_outs[2][5] ),
    .Y(_08960_));
 sky130_fd_sc_hd__and2b_2 _22215_ (.A_N(\systolic_inst.A_outs[2][0] ),
    .B(\systolic_inst.B_outs[2][7] ),
    .X(_08961_));
 sky130_fd_sc_hd__and3_2 _22216_ (.A(\systolic_inst.A_outs[2][1] ),
    .B(\systolic_inst.B_outs[2][6] ),
    .C(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__xnor2_2 _22217_ (.A(_08928_),
    .B(_08961_),
    .Y(_08963_));
 sky130_fd_sc_hd__xnor2_2 _22218_ (.A(_08960_),
    .B(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__xnor2_2 _22219_ (.A(_08929_),
    .B(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__nor2_2 _22220_ (.A(_08959_),
    .B(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__xnor2_2 _22221_ (.A(_08959_),
    .B(_08965_),
    .Y(_08967_));
 sky130_fd_sc_hd__or2_2 _22222_ (.A(_08931_),
    .B(_08967_),
    .X(_08968_));
 sky130_fd_sc_hd__and2_2 _22223_ (.A(_08931_),
    .B(_08967_),
    .X(_08969_));
 sky130_fd_sc_hd__xor2_2 _22224_ (.A(_08931_),
    .B(_08967_),
    .X(_08970_));
 sky130_fd_sc_hd__xnor2_2 _22225_ (.A(_08954_),
    .B(_08970_),
    .Y(_08971_));
 sky130_fd_sc_hd__and2b_2 _22226_ (.A_N(_08933_),
    .B(_08935_),
    .X(_08972_));
 sky130_fd_sc_hd__nand2b_2 _22227_ (.A_N(_08972_),
    .B(_08971_),
    .Y(_08973_));
 sky130_fd_sc_hd__xnor2_2 _22228_ (.A(_08971_),
    .B(_08972_),
    .Y(_08974_));
 sky130_fd_sc_hd__nand2b_2 _22229_ (.A_N(_08946_),
    .B(_08974_),
    .Y(_08975_));
 sky130_fd_sc_hd__xnor2_2 _22230_ (.A(_08946_),
    .B(_08974_),
    .Y(_08976_));
 sky130_fd_sc_hd__and2b_2 _22231_ (.A_N(_08945_),
    .B(_08976_),
    .X(_08977_));
 sky130_fd_sc_hd__xnor2_2 _22232_ (.A(_08945_),
    .B(_08976_),
    .Y(_08978_));
 sky130_fd_sc_hd__a31o_2 _22233_ (.A1(_08911_),
    .A2(_08912_),
    .A3(_08943_),
    .B1(_08941_),
    .X(_08979_));
 sky130_fd_sc_hd__xor2_2 _22234_ (.A(_08978_),
    .B(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__mux2_1 _22235_ (.A0(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[7] ),
    .A1(_08980_),
    .S(\systolic_inst.ce_local ),
    .X(_01801_));
 sky130_fd_sc_hd__a21bo_2 _22236_ (.A1(_08918_),
    .A2(_08953_),
    .B1_N(_08952_),
    .X(_08981_));
 sky130_fd_sc_hd__a21bo_2 _22237_ (.A1(\systolic_inst.B_outs[2][7] ),
    .A2(_08948_),
    .B1_N(_08949_),
    .X(_08982_));
 sky130_fd_sc_hd__o21bai_2 _22238_ (.A1(_08955_),
    .A2(_08957_),
    .B1_N(_08956_),
    .Y(_08983_));
 sky130_fd_sc_hd__o21a_2 _22239_ (.A1(\systolic_inst.B_outs[2][0] ),
    .A2(\systolic_inst.B_outs[2][1] ),
    .B1(\systolic_inst.A_outs[2][7] ),
    .X(_08984_));
 sky130_fd_sc_hd__o21ai_2 _22240_ (.A1(\systolic_inst.B_outs[2][0] ),
    .A2(\systolic_inst.B_outs[2][1] ),
    .B1(\systolic_inst.A_outs[2][7] ),
    .Y(_08985_));
 sky130_fd_sc_hd__a21o_2 _22241_ (.A1(\systolic_inst.B_outs[2][0] ),
    .A2(\systolic_inst.B_outs[2][1] ),
    .B1(_08985_),
    .X(_08986_));
 sky130_fd_sc_hd__and2b_2 _22242_ (.A_N(_08986_),
    .B(_08983_),
    .X(_08987_));
 sky130_fd_sc_hd__xnor2_2 _22243_ (.A(_08983_),
    .B(_08986_),
    .Y(_08988_));
 sky130_fd_sc_hd__xnor2_2 _22244_ (.A(_08982_),
    .B(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__and4_2 _22245_ (.A(\systolic_inst.B_outs[2][3] ),
    .B(\systolic_inst.B_outs[2][4] ),
    .C(\systolic_inst.A_outs[2][4] ),
    .D(\systolic_inst.A_outs[2][5] ),
    .X(_08990_));
 sky130_fd_sc_hd__a22oi_2 _22246_ (.A1(\systolic_inst.B_outs[2][4] ),
    .A2(\systolic_inst.A_outs[2][4] ),
    .B1(\systolic_inst.A_outs[2][5] ),
    .B2(\systolic_inst.B_outs[2][3] ),
    .Y(_08991_));
 sky130_fd_sc_hd__nor2_2 _22247_ (.A(_08990_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__nand2_2 _22248_ (.A(\systolic_inst.B_outs[2][2] ),
    .B(\systolic_inst.A_outs[2][6] ),
    .Y(_08993_));
 sky130_fd_sc_hd__xnor2_2 _22249_ (.A(_08992_),
    .B(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__nand2_2 _22250_ (.A(\systolic_inst.A_outs[2][3] ),
    .B(\systolic_inst.B_outs[2][5] ),
    .Y(_08995_));
 sky130_fd_sc_hd__and4b_2 _22251_ (.A_N(\systolic_inst.A_outs[2][1] ),
    .B(\systolic_inst.A_outs[2][2] ),
    .C(\systolic_inst.B_outs[2][6] ),
    .D(\systolic_inst.B_outs[2][7] ),
    .X(_08996_));
 sky130_fd_sc_hd__o2bb2a_2 _22252_ (.A1_N(\systolic_inst.A_outs[2][2] ),
    .A2_N(\systolic_inst.B_outs[2][6] ),
    .B1(_11265_),
    .B2(\systolic_inst.A_outs[2][1] ),
    .X(_08997_));
 sky130_fd_sc_hd__nor2_2 _22253_ (.A(_08996_),
    .B(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__xnor2_2 _22254_ (.A(_08995_),
    .B(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__a31oi_2 _22255_ (.A1(\systolic_inst.A_outs[2][2] ),
    .A2(\systolic_inst.B_outs[2][5] ),
    .A3(_08963_),
    .B1(_08962_),
    .Y(_09000_));
 sky130_fd_sc_hd__nand2b_2 _22256_ (.A_N(_09000_),
    .B(_08999_),
    .Y(_09001_));
 sky130_fd_sc_hd__xnor2_2 _22257_ (.A(_08999_),
    .B(_09000_),
    .Y(_09002_));
 sky130_fd_sc_hd__nand2_2 _22258_ (.A(_08994_),
    .B(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__xnor2_2 _22259_ (.A(_08994_),
    .B(_09002_),
    .Y(_09004_));
 sky130_fd_sc_hd__a21oi_2 _22260_ (.A1(_08929_),
    .A2(_08964_),
    .B1(_08966_),
    .Y(_09005_));
 sky130_fd_sc_hd__xnor2_2 _22261_ (.A(_09004_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__or2_2 _22262_ (.A(_08989_),
    .B(_09006_),
    .X(_09007_));
 sky130_fd_sc_hd__xor2_2 _22263_ (.A(_08989_),
    .B(_09006_),
    .X(_09008_));
 sky130_fd_sc_hd__o21a_2 _22264_ (.A1(_08954_),
    .A2(_08969_),
    .B1(_08968_),
    .X(_09009_));
 sky130_fd_sc_hd__nand2b_2 _22265_ (.A_N(_09009_),
    .B(_09008_),
    .Y(_09010_));
 sky130_fd_sc_hd__xor2_2 _22266_ (.A(_09008_),
    .B(_09009_),
    .X(_09011_));
 sky130_fd_sc_hd__nand2b_2 _22267_ (.A_N(_09011_),
    .B(_08981_),
    .Y(_09012_));
 sky130_fd_sc_hd__xor2_2 _22268_ (.A(_08981_),
    .B(_09011_),
    .X(_09013_));
 sky130_fd_sc_hd__and2_2 _22269_ (.A(_08973_),
    .B(_08975_),
    .X(_09014_));
 sky130_fd_sc_hd__xor2_2 _22270_ (.A(_09013_),
    .B(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__a21oi_2 _22271_ (.A1(_08978_),
    .A2(_08979_),
    .B1(_08977_),
    .Y(_09016_));
 sky130_fd_sc_hd__nand2b_2 _22272_ (.A_N(_09016_),
    .B(_09015_),
    .Y(_09017_));
 sky130_fd_sc_hd__nand2b_2 _22273_ (.A_N(_09015_),
    .B(_09016_),
    .Y(_09018_));
 sky130_fd_sc_hd__and2_2 _22274_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[8] ),
    .X(_09019_));
 sky130_fd_sc_hd__a31o_2 _22275_ (.A1(\systolic_inst.ce_local ),
    .A2(_09017_),
    .A3(_09018_),
    .B1(_09019_),
    .X(_01802_));
 sky130_fd_sc_hd__a21o_2 _22276_ (.A1(_08982_),
    .A2(_08988_),
    .B1(_08987_),
    .X(_09020_));
 sky130_fd_sc_hd__o21ba_2 _22277_ (.A1(_08991_),
    .A2(_08993_),
    .B1_N(_08990_),
    .X(_09021_));
 sky130_fd_sc_hd__nor2_2 _22278_ (.A(_08985_),
    .B(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__and2_2 _22279_ (.A(_08985_),
    .B(_09021_),
    .X(_09023_));
 sky130_fd_sc_hd__or2_2 _22280_ (.A(_09022_),
    .B(_09023_),
    .X(_09024_));
 sky130_fd_sc_hd__nand2_2 _22281_ (.A(\systolic_inst.B_outs[2][2] ),
    .B(\systolic_inst.A_outs[2][7] ),
    .Y(_09025_));
 sky130_fd_sc_hd__a22oi_2 _22282_ (.A1(\systolic_inst.B_outs[2][4] ),
    .A2(\systolic_inst.A_outs[2][5] ),
    .B1(\systolic_inst.A_outs[2][6] ),
    .B2(\systolic_inst.B_outs[2][3] ),
    .Y(_09026_));
 sky130_fd_sc_hd__and4_2 _22283_ (.A(\systolic_inst.B_outs[2][3] ),
    .B(\systolic_inst.B_outs[2][4] ),
    .C(\systolic_inst.A_outs[2][5] ),
    .D(\systolic_inst.A_outs[2][6] ),
    .X(_09027_));
 sky130_fd_sc_hd__nor2_2 _22284_ (.A(_09026_),
    .B(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__xnor2_2 _22285_ (.A(_09025_),
    .B(_09028_),
    .Y(_09029_));
 sky130_fd_sc_hd__nand2_2 _22286_ (.A(\systolic_inst.A_outs[2][4] ),
    .B(\systolic_inst.B_outs[2][5] ),
    .Y(_09030_));
 sky130_fd_sc_hd__and4b_2 _22287_ (.A_N(\systolic_inst.A_outs[2][2] ),
    .B(\systolic_inst.A_outs[2][3] ),
    .C(\systolic_inst.B_outs[2][6] ),
    .D(\systolic_inst.B_outs[2][7] ),
    .X(_09031_));
 sky130_fd_sc_hd__o2bb2a_2 _22288_ (.A1_N(\systolic_inst.A_outs[2][3] ),
    .A2_N(\systolic_inst.B_outs[2][6] ),
    .B1(_11265_),
    .B2(\systolic_inst.A_outs[2][2] ),
    .X(_09032_));
 sky130_fd_sc_hd__nor2_2 _22289_ (.A(_09031_),
    .B(_09032_),
    .Y(_09033_));
 sky130_fd_sc_hd__xnor2_2 _22290_ (.A(_09030_),
    .B(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__o21ba_2 _22291_ (.A1(_08995_),
    .A2(_08997_),
    .B1_N(_08996_),
    .X(_09035_));
 sky130_fd_sc_hd__nand2b_2 _22292_ (.A_N(_09035_),
    .B(_09034_),
    .Y(_09036_));
 sky130_fd_sc_hd__xnor2_2 _22293_ (.A(_09034_),
    .B(_09035_),
    .Y(_09037_));
 sky130_fd_sc_hd__xnor2_2 _22294_ (.A(_09029_),
    .B(_09037_),
    .Y(_09038_));
 sky130_fd_sc_hd__a21o_2 _22295_ (.A1(_09001_),
    .A2(_09003_),
    .B1(_09038_),
    .X(_09039_));
 sky130_fd_sc_hd__nand3_2 _22296_ (.A(_09001_),
    .B(_09003_),
    .C(_09038_),
    .Y(_09040_));
 sky130_fd_sc_hd__nand2_2 _22297_ (.A(_09039_),
    .B(_09040_),
    .Y(_09041_));
 sky130_fd_sc_hd__xor2_2 _22298_ (.A(_09024_),
    .B(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__o21a_2 _22299_ (.A1(_09004_),
    .A2(_09005_),
    .B1(_09007_),
    .X(_09043_));
 sky130_fd_sc_hd__nand2b_2 _22300_ (.A_N(_09043_),
    .B(_09042_),
    .Y(_09044_));
 sky130_fd_sc_hd__xnor2_2 _22301_ (.A(_09042_),
    .B(_09043_),
    .Y(_09045_));
 sky130_fd_sc_hd__xnor2_2 _22302_ (.A(_09020_),
    .B(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__nand3_2 _22303_ (.A(_09010_),
    .B(_09012_),
    .C(_09046_),
    .Y(_09047_));
 sky130_fd_sc_hd__inv_2 _22304_ (.A(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__a21oi_2 _22305_ (.A1(_09010_),
    .A2(_09012_),
    .B1(_09046_),
    .Y(_09049_));
 sky130_fd_sc_hd__inv_2 _22306_ (.A(_09049_),
    .Y(_09050_));
 sky130_fd_sc_hd__o21a_2 _22307_ (.A1(_09013_),
    .A2(_09014_),
    .B1(_09017_),
    .X(_09051_));
 sky130_fd_sc_hd__nor2_2 _22308_ (.A(_09048_),
    .B(_09049_),
    .Y(_09052_));
 sky130_fd_sc_hd__and3_2 _22309_ (.A(_09047_),
    .B(_09050_),
    .C(_09051_),
    .X(_09053_));
 sky130_fd_sc_hd__o21ai_2 _22310_ (.A1(_09051_),
    .A2(_09052_),
    .B1(\systolic_inst.ce_local ),
    .Y(_09054_));
 sky130_fd_sc_hd__o22a_2 _22311_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[9] ),
    .B1(_09053_),
    .B2(_09054_),
    .X(_01803_));
 sky130_fd_sc_hd__o21ba_2 _22312_ (.A1(_09025_),
    .A2(_09026_),
    .B1_N(_09027_),
    .X(_09055_));
 sky130_fd_sc_hd__nor2_2 _22313_ (.A(_08985_),
    .B(_09055_),
    .Y(_09056_));
 sky130_fd_sc_hd__and2_2 _22314_ (.A(_08985_),
    .B(_09055_),
    .X(_09057_));
 sky130_fd_sc_hd__or2_2 _22315_ (.A(_09056_),
    .B(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__a22o_2 _22316_ (.A1(\systolic_inst.B_outs[2][4] ),
    .A2(\systolic_inst.A_outs[2][6] ),
    .B1(\systolic_inst.A_outs[2][7] ),
    .B2(\systolic_inst.B_outs[2][3] ),
    .X(_09059_));
 sky130_fd_sc_hd__and3_2 _22317_ (.A(\systolic_inst.B_outs[2][3] ),
    .B(\systolic_inst.B_outs[2][4] ),
    .C(\systolic_inst.A_outs[2][7] ),
    .X(_09060_));
 sky130_fd_sc_hd__a21bo_2 _22318_ (.A1(\systolic_inst.A_outs[2][6] ),
    .A2(_09060_),
    .B1_N(_09059_),
    .X(_09061_));
 sky130_fd_sc_hd__xor2_2 _22319_ (.A(_09025_),
    .B(_09061_),
    .X(_09062_));
 sky130_fd_sc_hd__nand2_2 _22320_ (.A(\systolic_inst.B_outs[2][5] ),
    .B(\systolic_inst.A_outs[2][5] ),
    .Y(_09063_));
 sky130_fd_sc_hd__and4b_2 _22321_ (.A_N(\systolic_inst.A_outs[2][3] ),
    .B(\systolic_inst.A_outs[2][4] ),
    .C(\systolic_inst.B_outs[2][6] ),
    .D(\systolic_inst.B_outs[2][7] ),
    .X(_09064_));
 sky130_fd_sc_hd__o2bb2a_2 _22322_ (.A1_N(\systolic_inst.A_outs[2][4] ),
    .A2_N(\systolic_inst.B_outs[2][6] ),
    .B1(_11265_),
    .B2(\systolic_inst.A_outs[2][3] ),
    .X(_09065_));
 sky130_fd_sc_hd__nor2_2 _22323_ (.A(_09064_),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__xnor2_2 _22324_ (.A(_09063_),
    .B(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__o21ba_2 _22325_ (.A1(_09030_),
    .A2(_09032_),
    .B1_N(_09031_),
    .X(_09068_));
 sky130_fd_sc_hd__nand2b_2 _22326_ (.A_N(_09068_),
    .B(_09067_),
    .Y(_09069_));
 sky130_fd_sc_hd__xnor2_2 _22327_ (.A(_09067_),
    .B(_09068_),
    .Y(_09070_));
 sky130_fd_sc_hd__nand2_2 _22328_ (.A(_09062_),
    .B(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__or2_2 _22329_ (.A(_09062_),
    .B(_09070_),
    .X(_09072_));
 sky130_fd_sc_hd__nand2_2 _22330_ (.A(_09071_),
    .B(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__a21bo_2 _22331_ (.A1(_09029_),
    .A2(_09037_),
    .B1_N(_09036_),
    .X(_09074_));
 sky130_fd_sc_hd__nand2b_2 _22332_ (.A_N(_09073_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__xor2_2 _22333_ (.A(_09073_),
    .B(_09074_),
    .X(_09076_));
 sky130_fd_sc_hd__xor2_2 _22334_ (.A(_09058_),
    .B(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__o21a_2 _22335_ (.A1(_09024_),
    .A2(_09041_),
    .B1(_09039_),
    .X(_09078_));
 sky130_fd_sc_hd__nand2b_2 _22336_ (.A_N(_09078_),
    .B(_09077_),
    .Y(_09079_));
 sky130_fd_sc_hd__xnor2_2 _22337_ (.A(_09077_),
    .B(_09078_),
    .Y(_09080_));
 sky130_fd_sc_hd__nand2_2 _22338_ (.A(_09022_),
    .B(_09080_),
    .Y(_09081_));
 sky130_fd_sc_hd__or2_2 _22339_ (.A(_09022_),
    .B(_09080_),
    .X(_09082_));
 sky130_fd_sc_hd__nand2_2 _22340_ (.A(_09081_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__a21boi_2 _22341_ (.A1(_09020_),
    .A2(_09045_),
    .B1_N(_09044_),
    .Y(_09084_));
 sky130_fd_sc_hd__nor2_2 _22342_ (.A(_09083_),
    .B(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__xnor2_2 _22343_ (.A(_09083_),
    .B(_09084_),
    .Y(_09086_));
 sky130_fd_sc_hd__a21o_2 _22344_ (.A1(_09050_),
    .A2(_09051_),
    .B1(_09048_),
    .X(_09087_));
 sky130_fd_sc_hd__a211oi_2 _22345_ (.A1(_09050_),
    .A2(_09051_),
    .B1(_09086_),
    .C1(_09048_),
    .Y(_09088_));
 sky130_fd_sc_hd__xor2_2 _22346_ (.A(_09086_),
    .B(_09087_),
    .X(_09089_));
 sky130_fd_sc_hd__mux2_1 _22347_ (.A0(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[10] ),
    .A1(_09089_),
    .S(\systolic_inst.ce_local ),
    .X(_01804_));
 sky130_fd_sc_hd__o2bb2a_2 _22348_ (.A1_N(\systolic_inst.A_outs[2][6] ),
    .A2_N(_09060_),
    .B1(_09061_),
    .B2(_09025_),
    .X(_09090_));
 sky130_fd_sc_hd__or2_2 _22349_ (.A(_08985_),
    .B(_09090_),
    .X(_09091_));
 sky130_fd_sc_hd__nand2_2 _22350_ (.A(_08985_),
    .B(_09090_),
    .Y(_09092_));
 sky130_fd_sc_hd__nand2_2 _22351_ (.A(_09091_),
    .B(_09092_),
    .Y(_09093_));
 sky130_fd_sc_hd__or2_2 _22352_ (.A(\systolic_inst.B_outs[2][3] ),
    .B(\systolic_inst.B_outs[2][4] ),
    .X(_09094_));
 sky130_fd_sc_hd__and3b_2 _22353_ (.A_N(_09060_),
    .B(_09094_),
    .C(\systolic_inst.A_outs[2][7] ),
    .X(_09095_));
 sky130_fd_sc_hd__xnor2_2 _22354_ (.A(_09025_),
    .B(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__nand2_2 _22355_ (.A(\systolic_inst.B_outs[2][5] ),
    .B(\systolic_inst.A_outs[2][6] ),
    .Y(_09097_));
 sky130_fd_sc_hd__and4b_2 _22356_ (.A_N(\systolic_inst.A_outs[2][4] ),
    .B(\systolic_inst.A_outs[2][5] ),
    .C(\systolic_inst.B_outs[2][6] ),
    .D(\systolic_inst.B_outs[2][7] ),
    .X(_09098_));
 sky130_fd_sc_hd__o2bb2a_2 _22357_ (.A1_N(\systolic_inst.A_outs[2][5] ),
    .A2_N(\systolic_inst.B_outs[2][6] ),
    .B1(_11265_),
    .B2(\systolic_inst.A_outs[2][4] ),
    .X(_09099_));
 sky130_fd_sc_hd__or2_2 _22358_ (.A(_09098_),
    .B(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__xor2_2 _22359_ (.A(_09097_),
    .B(_09100_),
    .X(_09101_));
 sky130_fd_sc_hd__o21ba_2 _22360_ (.A1(_09063_),
    .A2(_09065_),
    .B1_N(_09064_),
    .X(_09102_));
 sky130_fd_sc_hd__nand2b_2 _22361_ (.A_N(_09102_),
    .B(_09101_),
    .Y(_09103_));
 sky130_fd_sc_hd__xnor2_2 _22362_ (.A(_09101_),
    .B(_09102_),
    .Y(_09104_));
 sky130_fd_sc_hd__nand2_2 _22363_ (.A(_09096_),
    .B(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__xnor2_2 _22364_ (.A(_09096_),
    .B(_09104_),
    .Y(_09106_));
 sky130_fd_sc_hd__a21o_2 _22365_ (.A1(_09069_),
    .A2(_09071_),
    .B1(_09106_),
    .X(_09107_));
 sky130_fd_sc_hd__nand3_2 _22366_ (.A(_09069_),
    .B(_09071_),
    .C(_09106_),
    .Y(_09108_));
 sky130_fd_sc_hd__nand2_2 _22367_ (.A(_09107_),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__xor2_2 _22368_ (.A(_09093_),
    .B(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__o21a_2 _22369_ (.A1(_09058_),
    .A2(_09076_),
    .B1(_09075_),
    .X(_09111_));
 sky130_fd_sc_hd__and2b_2 _22370_ (.A_N(_09111_),
    .B(_09110_),
    .X(_09112_));
 sky130_fd_sc_hd__and2b_2 _22371_ (.A_N(_09110_),
    .B(_09111_),
    .X(_09113_));
 sky130_fd_sc_hd__nor2_2 _22372_ (.A(_09112_),
    .B(_09113_),
    .Y(_09114_));
 sky130_fd_sc_hd__xnor2_2 _22373_ (.A(_09056_),
    .B(_09114_),
    .Y(_09115_));
 sky130_fd_sc_hd__nand3_2 _22374_ (.A(_09079_),
    .B(_09081_),
    .C(_09115_),
    .Y(_09116_));
 sky130_fd_sc_hd__inv_2 _22375_ (.A(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__a21oi_2 _22376_ (.A1(_09079_),
    .A2(_09081_),
    .B1(_09115_),
    .Y(_09118_));
 sky130_fd_sc_hd__o22a_2 _22377_ (.A1(_09085_),
    .A2(_09088_),
    .B1(_09117_),
    .B2(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__or4_2 _22378_ (.A(_09085_),
    .B(_09088_),
    .C(_09117_),
    .D(_09118_),
    .X(_09120_));
 sky130_fd_sc_hd__nand2_2 _22379_ (.A(\systolic_inst.ce_local ),
    .B(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__o22a_2 _22380_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[11] ),
    .B1(_09119_),
    .B2(_09121_),
    .X(_01805_));
 sky130_fd_sc_hd__a31o_2 _22381_ (.A1(\systolic_inst.B_outs[2][2] ),
    .A2(\systolic_inst.A_outs[2][7] ),
    .A3(_09094_),
    .B1(_09060_),
    .X(_09122_));
 sky130_fd_sc_hd__or2_2 _22382_ (.A(_08984_),
    .B(_09122_),
    .X(_09123_));
 sky130_fd_sc_hd__nand2_2 _22383_ (.A(_08984_),
    .B(_09122_),
    .Y(_09124_));
 sky130_fd_sc_hd__nand2_2 _22384_ (.A(_09123_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__inv_2 _22385_ (.A(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__o2bb2a_2 _22386_ (.A1_N(\systolic_inst.B_outs[2][6] ),
    .A2_N(\systolic_inst.A_outs[2][6] ),
    .B1(_11265_),
    .B2(\systolic_inst.A_outs[2][5] ),
    .X(_09127_));
 sky130_fd_sc_hd__and4b_2 _22387_ (.A_N(\systolic_inst.A_outs[2][5] ),
    .B(\systolic_inst.B_outs[2][6] ),
    .C(\systolic_inst.A_outs[2][6] ),
    .D(\systolic_inst.B_outs[2][7] ),
    .X(_09128_));
 sky130_fd_sc_hd__nor2_2 _22388_ (.A(_09127_),
    .B(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__nand2_2 _22389_ (.A(\systolic_inst.B_outs[2][5] ),
    .B(\systolic_inst.A_outs[2][7] ),
    .Y(_09130_));
 sky130_fd_sc_hd__and3_2 _22390_ (.A(\systolic_inst.B_outs[2][5] ),
    .B(\systolic_inst.A_outs[2][7] ),
    .C(_09129_),
    .X(_09131_));
 sky130_fd_sc_hd__xnor2_2 _22391_ (.A(_09129_),
    .B(_09130_),
    .Y(_09132_));
 sky130_fd_sc_hd__o21ba_2 _22392_ (.A1(_09097_),
    .A2(_09099_),
    .B1_N(_09098_),
    .X(_09133_));
 sky130_fd_sc_hd__nand2b_2 _22393_ (.A_N(_09133_),
    .B(_09132_),
    .Y(_09134_));
 sky130_fd_sc_hd__xnor2_2 _22394_ (.A(_09132_),
    .B(_09133_),
    .Y(_09135_));
 sky130_fd_sc_hd__xnor2_2 _22395_ (.A(_09096_),
    .B(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__a21o_2 _22396_ (.A1(_09103_),
    .A2(_09105_),
    .B1(_09136_),
    .X(_09137_));
 sky130_fd_sc_hd__nand3_2 _22397_ (.A(_09103_),
    .B(_09105_),
    .C(_09136_),
    .Y(_09138_));
 sky130_fd_sc_hd__nand2_2 _22398_ (.A(_09137_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__xnor2_2 _22399_ (.A(_09126_),
    .B(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__o21a_2 _22400_ (.A1(_09093_),
    .A2(_09109_),
    .B1(_09107_),
    .X(_09141_));
 sky130_fd_sc_hd__and2b_2 _22401_ (.A_N(_09141_),
    .B(_09140_),
    .X(_09142_));
 sky130_fd_sc_hd__and2b_2 _22402_ (.A_N(_09140_),
    .B(_09141_),
    .X(_09143_));
 sky130_fd_sc_hd__nor2_2 _22403_ (.A(_09142_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__and2b_2 _22404_ (.A_N(_09091_),
    .B(_09144_),
    .X(_09145_));
 sky130_fd_sc_hd__xor2_2 _22405_ (.A(_09091_),
    .B(_09144_),
    .X(_09146_));
 sky130_fd_sc_hd__a21oi_2 _22406_ (.A1(_09056_),
    .A2(_09114_),
    .B1(_09112_),
    .Y(_09147_));
 sky130_fd_sc_hd__nor2_2 _22407_ (.A(_09146_),
    .B(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__and2_2 _22408_ (.A(_09146_),
    .B(_09147_),
    .X(_09149_));
 sky130_fd_sc_hd__nor2_2 _22409_ (.A(_09148_),
    .B(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__o31a_2 _22410_ (.A1(_09085_),
    .A2(_09088_),
    .A3(_09118_),
    .B1(_09116_),
    .X(_09151_));
 sky130_fd_sc_hd__o311a_2 _22411_ (.A1(_09085_),
    .A2(_09088_),
    .A3(_09118_),
    .B1(_09150_),
    .C1(_09116_),
    .X(_09152_));
 sky130_fd_sc_hd__xor2_2 _22412_ (.A(_09150_),
    .B(_09151_),
    .X(_09153_));
 sky130_fd_sc_hd__mux2_1 _22413_ (.A0(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[12] ),
    .A1(_09153_),
    .S(\systolic_inst.ce_local ),
    .X(_01806_));
 sky130_fd_sc_hd__nand2_2 _22414_ (.A(\systolic_inst.B_outs[2][6] ),
    .B(\systolic_inst.A_outs[2][7] ),
    .Y(_09154_));
 sky130_fd_sc_hd__nor2_2 _22415_ (.A(\systolic_inst.A_outs[2][6] ),
    .B(_11265_),
    .Y(_09155_));
 sky130_fd_sc_hd__xnor2_2 _22416_ (.A(_09154_),
    .B(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__nand2b_2 _22417_ (.A_N(_09130_),
    .B(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__xnor2_2 _22418_ (.A(_09130_),
    .B(_09156_),
    .Y(_09158_));
 sky130_fd_sc_hd__o21ai_2 _22419_ (.A1(_09128_),
    .A2(_09131_),
    .B1(_09158_),
    .Y(_09159_));
 sky130_fd_sc_hd__or3_2 _22420_ (.A(_09128_),
    .B(_09131_),
    .C(_09158_),
    .X(_09160_));
 sky130_fd_sc_hd__and2_2 _22421_ (.A(_09159_),
    .B(_09160_),
    .X(_09161_));
 sky130_fd_sc_hd__nand2_2 _22422_ (.A(_09096_),
    .B(_09161_),
    .Y(_09162_));
 sky130_fd_sc_hd__or2_2 _22423_ (.A(_09096_),
    .B(_09161_),
    .X(_09163_));
 sky130_fd_sc_hd__nand2_2 _22424_ (.A(_09162_),
    .B(_09163_),
    .Y(_09164_));
 sky130_fd_sc_hd__a21bo_2 _22425_ (.A1(_09096_),
    .A2(_09135_),
    .B1_N(_09134_),
    .X(_09165_));
 sky130_fd_sc_hd__nand2b_2 _22426_ (.A_N(_09164_),
    .B(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__xor2_2 _22427_ (.A(_09164_),
    .B(_09165_),
    .X(_09167_));
 sky130_fd_sc_hd__xnor2_2 _22428_ (.A(_09126_),
    .B(_09167_),
    .Y(_09168_));
 sky130_fd_sc_hd__o21a_2 _22429_ (.A1(_09125_),
    .A2(_09139_),
    .B1(_09137_),
    .X(_09169_));
 sky130_fd_sc_hd__and2b_2 _22430_ (.A_N(_09169_),
    .B(_09168_),
    .X(_09170_));
 sky130_fd_sc_hd__and2b_2 _22431_ (.A_N(_09168_),
    .B(_09169_),
    .X(_09171_));
 sky130_fd_sc_hd__nor2_2 _22432_ (.A(_09170_),
    .B(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__xnor2_2 _22433_ (.A(_09124_),
    .B(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__o21a_2 _22434_ (.A1(_09142_),
    .A2(_09145_),
    .B1(_09173_),
    .X(_09174_));
 sky130_fd_sc_hd__or3_2 _22435_ (.A(_09142_),
    .B(_09145_),
    .C(_09173_),
    .X(_09175_));
 sky130_fd_sc_hd__and2b_2 _22436_ (.A_N(_09174_),
    .B(_09175_),
    .X(_09176_));
 sky130_fd_sc_hd__nor2_2 _22437_ (.A(_09148_),
    .B(_09152_),
    .Y(_09177_));
 sky130_fd_sc_hd__xnor2_2 _22438_ (.A(_09176_),
    .B(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__mux2_1 _22439_ (.A0(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[13] ),
    .A1(_09178_),
    .S(\systolic_inst.ce_local ),
    .X(_01807_));
 sky130_fd_sc_hd__o211ai_2 _22440_ (.A1(_11265_),
    .A2(\systolic_inst.A_outs[2][7] ),
    .B1(_09130_),
    .C1(_09154_),
    .Y(_09179_));
 sky130_fd_sc_hd__o311a_2 _22441_ (.A1(\systolic_inst.A_outs[2][6] ),
    .A2(_11265_),
    .A3(_09154_),
    .B1(_09157_),
    .C1(_09179_),
    .X(_09180_));
 sky130_fd_sc_hd__a31o_2 _22442_ (.A1(\systolic_inst.B_outs[2][5] ),
    .A2(\systolic_inst.B_outs[2][6] ),
    .A3(\systolic_inst.A_outs[2][7] ),
    .B1(_09180_),
    .X(_09181_));
 sky130_fd_sc_hd__or2_2 _22443_ (.A(_09096_),
    .B(_09181_),
    .X(_09182_));
 sky130_fd_sc_hd__nand2_2 _22444_ (.A(_09096_),
    .B(_09181_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand2_2 _22445_ (.A(_09182_),
    .B(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__a21oi_2 _22446_ (.A1(_09159_),
    .A2(_09162_),
    .B1(_09184_),
    .Y(_09185_));
 sky130_fd_sc_hd__and3_2 _22447_ (.A(_09159_),
    .B(_09162_),
    .C(_09184_),
    .X(_09186_));
 sky130_fd_sc_hd__nor2_2 _22448_ (.A(_09185_),
    .B(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__xnor2_2 _22449_ (.A(_09125_),
    .B(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__o21a_2 _22450_ (.A1(_09125_),
    .A2(_09167_),
    .B1(_09166_),
    .X(_09189_));
 sky130_fd_sc_hd__and2b_2 _22451_ (.A_N(_09189_),
    .B(_09188_),
    .X(_09190_));
 sky130_fd_sc_hd__and2b_2 _22452_ (.A_N(_09188_),
    .B(_09189_),
    .X(_09191_));
 sky130_fd_sc_hd__nor2_2 _22453_ (.A(_09190_),
    .B(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__xnor2_2 _22454_ (.A(_09124_),
    .B(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__o21ba_2 _22455_ (.A1(_09124_),
    .A2(_09171_),
    .B1_N(_09170_),
    .X(_09194_));
 sky130_fd_sc_hd__and2b_2 _22456_ (.A_N(_09194_),
    .B(_09193_),
    .X(_09195_));
 sky130_fd_sc_hd__xnor2_2 _22457_ (.A(_09193_),
    .B(_09194_),
    .Y(_09196_));
 sky130_fd_sc_hd__o31a_2 _22458_ (.A1(_09148_),
    .A2(_09152_),
    .A3(_09174_),
    .B1(_09175_),
    .X(_09197_));
 sky130_fd_sc_hd__xor2_2 _22459_ (.A(_09196_),
    .B(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__mux2_1 _22460_ (.A0(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[14] ),
    .A1(_09198_),
    .S(\systolic_inst.ce_local ),
    .X(_01808_));
 sky130_fd_sc_hd__a31oi_2 _22461_ (.A1(_08984_),
    .A2(_09122_),
    .A3(_09192_),
    .B1(_09190_),
    .Y(_09199_));
 sky130_fd_sc_hd__a21oi_2 _22462_ (.A1(_09126_),
    .A2(_09187_),
    .B1(_09185_),
    .Y(_09200_));
 sky130_fd_sc_hd__xnor2_2 _22463_ (.A(_09123_),
    .B(_09182_),
    .Y(_09201_));
 sky130_fd_sc_hd__xnor2_2 _22464_ (.A(_09200_),
    .B(_09201_),
    .Y(_09202_));
 sky130_fd_sc_hd__xnor2_2 _22465_ (.A(_09199_),
    .B(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__a211o_2 _22466_ (.A1(_09196_),
    .A2(_09197_),
    .B1(_11258_),
    .C1(_09195_),
    .X(_09204_));
 sky130_fd_sc_hd__a2bb2o_2 _22467_ (.A1_N(_09204_),
    .A2_N(_09203_),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B2(_11258_),
    .X(_01809_));
 sky130_fd_sc_hd__a21o_2 _22468_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[2][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_09205_));
 sky130_fd_sc_hd__a21oi_2 _22469_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[2][0] ),
    .Y(_09206_));
 sky130_fd_sc_hd__a21oi_2 _22470_ (.A1(\systolic_inst.ce_local ),
    .A2(_09205_),
    .B1(_09206_),
    .Y(_01810_));
 sky130_fd_sc_hd__and2_2 _22471_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[2][1] ),
    .X(_09207_));
 sky130_fd_sc_hd__nand2_2 _22472_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[2][1] ),
    .Y(_09208_));
 sky130_fd_sc_hd__or2_2 _22473_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[2][1] ),
    .X(_09209_));
 sky130_fd_sc_hd__and4_2 _22474_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[2][0] ),
    .C(_09208_),
    .D(_09209_),
    .X(_09210_));
 sky130_fd_sc_hd__inv_2 _22475_ (.A(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__a22o_2 _22476_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[2][0] ),
    .B1(_09208_),
    .B2(_09209_),
    .X(_09212_));
 sky130_fd_sc_hd__a32o_2 _22477_ (.A1(_11712_),
    .A2(_09211_),
    .A3(_09212_),
    .B1(\systolic_inst.acc_wires[2][1] ),
    .B2(_11258_),
    .X(_01811_));
 sky130_fd_sc_hd__nand2_2 _22478_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[2][2] ),
    .Y(_09213_));
 sky130_fd_sc_hd__or2_2 _22479_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[2][2] ),
    .X(_09214_));
 sky130_fd_sc_hd__a31o_2 _22480_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[2][0] ),
    .A3(_09209_),
    .B1(_09207_),
    .X(_09215_));
 sky130_fd_sc_hd__a21o_2 _22481_ (.A1(_09213_),
    .A2(_09214_),
    .B1(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__and3_2 _22482_ (.A(_09213_),
    .B(_09214_),
    .C(_09215_),
    .X(_09217_));
 sky130_fd_sc_hd__inv_2 _22483_ (.A(_09217_),
    .Y(_09218_));
 sky130_fd_sc_hd__a32o_2 _22484_ (.A1(_11712_),
    .A2(_09216_),
    .A3(_09218_),
    .B1(\systolic_inst.acc_wires[2][2] ),
    .B2(_11258_),
    .X(_01812_));
 sky130_fd_sc_hd__nand2_2 _22485_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[2][3] ),
    .Y(_09219_));
 sky130_fd_sc_hd__or2_2 _22486_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[2][3] ),
    .X(_09220_));
 sky130_fd_sc_hd__a21bo_2 _22487_ (.A1(_09214_),
    .A2(_09215_),
    .B1_N(_09213_),
    .X(_09221_));
 sky130_fd_sc_hd__a21o_2 _22488_ (.A1(_09219_),
    .A2(_09220_),
    .B1(_09221_),
    .X(_09222_));
 sky130_fd_sc_hd__and3_2 _22489_ (.A(_09219_),
    .B(_09220_),
    .C(_09221_),
    .X(_09223_));
 sky130_fd_sc_hd__inv_2 _22490_ (.A(_09223_),
    .Y(_09224_));
 sky130_fd_sc_hd__a32o_2 _22491_ (.A1(_11712_),
    .A2(_09222_),
    .A3(_09224_),
    .B1(\systolic_inst.acc_wires[2][3] ),
    .B2(_11258_),
    .X(_01813_));
 sky130_fd_sc_hd__nand2_2 _22492_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[2][4] ),
    .Y(_09225_));
 sky130_fd_sc_hd__or2_2 _22493_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[2][4] ),
    .X(_09226_));
 sky130_fd_sc_hd__a21bo_2 _22494_ (.A1(_09220_),
    .A2(_09221_),
    .B1_N(_09219_),
    .X(_09227_));
 sky130_fd_sc_hd__a21o_2 _22495_ (.A1(_09225_),
    .A2(_09226_),
    .B1(_09227_),
    .X(_09228_));
 sky130_fd_sc_hd__and3_2 _22496_ (.A(_09225_),
    .B(_09226_),
    .C(_09227_),
    .X(_09229_));
 sky130_fd_sc_hd__inv_2 _22497_ (.A(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__a32o_2 _22498_ (.A1(_11712_),
    .A2(_09228_),
    .A3(_09230_),
    .B1(\systolic_inst.acc_wires[2][4] ),
    .B2(_11258_),
    .X(_01814_));
 sky130_fd_sc_hd__nand2_2 _22499_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[2][5] ),
    .Y(_09231_));
 sky130_fd_sc_hd__or2_2 _22500_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[2][5] ),
    .X(_09232_));
 sky130_fd_sc_hd__a21bo_2 _22501_ (.A1(_09226_),
    .A2(_09227_),
    .B1_N(_09225_),
    .X(_09233_));
 sky130_fd_sc_hd__a21o_2 _22502_ (.A1(_09231_),
    .A2(_09232_),
    .B1(_09233_),
    .X(_09234_));
 sky130_fd_sc_hd__and3_2 _22503_ (.A(_09231_),
    .B(_09232_),
    .C(_09233_),
    .X(_09235_));
 sky130_fd_sc_hd__inv_2 _22504_ (.A(_09235_),
    .Y(_09236_));
 sky130_fd_sc_hd__a32o_2 _22505_ (.A1(_11712_),
    .A2(_09234_),
    .A3(_09236_),
    .B1(\systolic_inst.acc_wires[2][5] ),
    .B2(_11258_),
    .X(_01815_));
 sky130_fd_sc_hd__nand2_2 _22506_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[2][6] ),
    .Y(_09237_));
 sky130_fd_sc_hd__or2_2 _22507_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[2][6] ),
    .X(_09238_));
 sky130_fd_sc_hd__a21bo_2 _22508_ (.A1(_09232_),
    .A2(_09233_),
    .B1_N(_09231_),
    .X(_09239_));
 sky130_fd_sc_hd__a21o_2 _22509_ (.A1(_09237_),
    .A2(_09238_),
    .B1(_09239_),
    .X(_09240_));
 sky130_fd_sc_hd__and3_2 _22510_ (.A(_09237_),
    .B(_09238_),
    .C(_09239_),
    .X(_09241_));
 sky130_fd_sc_hd__inv_2 _22511_ (.A(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__a32o_2 _22512_ (.A1(_11712_),
    .A2(_09240_),
    .A3(_09242_),
    .B1(\systolic_inst.acc_wires[2][6] ),
    .B2(_11258_),
    .X(_01816_));
 sky130_fd_sc_hd__nand2_2 _22513_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[2][7] ),
    .Y(_09243_));
 sky130_fd_sc_hd__or2_2 _22514_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[2][7] ),
    .X(_09244_));
 sky130_fd_sc_hd__a21bo_2 _22515_ (.A1(_09238_),
    .A2(_09239_),
    .B1_N(_09237_),
    .X(_09245_));
 sky130_fd_sc_hd__a21o_2 _22516_ (.A1(_09243_),
    .A2(_09244_),
    .B1(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__nand3_2 _22517_ (.A(_09243_),
    .B(_09244_),
    .C(_09245_),
    .Y(_09247_));
 sky130_fd_sc_hd__a32o_2 _22518_ (.A1(_11712_),
    .A2(_09246_),
    .A3(_09247_),
    .B1(\systolic_inst.acc_wires[2][7] ),
    .B2(_11258_),
    .X(_01817_));
 sky130_fd_sc_hd__a21bo_2 _22519_ (.A1(_09244_),
    .A2(_09245_),
    .B1_N(_09243_),
    .X(_09248_));
 sky130_fd_sc_hd__xor2_2 _22520_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[2][8] ),
    .X(_09249_));
 sky130_fd_sc_hd__and2_2 _22521_ (.A(_09248_),
    .B(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__o21ai_2 _22522_ (.A1(_09248_),
    .A2(_09249_),
    .B1(_11712_),
    .Y(_09251_));
 sky130_fd_sc_hd__a2bb2o_2 _22523_ (.A1_N(_09251_),
    .A2_N(_09250_),
    .B1(\systolic_inst.acc_wires[2][8] ),
    .B2(_11258_),
    .X(_01818_));
 sky130_fd_sc_hd__xor2_2 _22524_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[2][9] ),
    .X(_09252_));
 sky130_fd_sc_hd__a211o_2 _22525_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[2][8] ),
    .B1(_09250_),
    .C1(_09252_),
    .X(_09253_));
 sky130_fd_sc_hd__nand2_2 _22526_ (.A(_09249_),
    .B(_09252_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand2_2 _22527_ (.A(_09250_),
    .B(_09252_),
    .Y(_09255_));
 sky130_fd_sc_hd__and3_2 _22528_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[2][8] ),
    .C(_09252_),
    .X(_09256_));
 sky130_fd_sc_hd__nor2_2 _22529_ (.A(_11713_),
    .B(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__a32o_2 _22530_ (.A1(_09253_),
    .A2(_09255_),
    .A3(_09257_),
    .B1(\systolic_inst.acc_wires[2][9] ),
    .B2(_11258_),
    .X(_01819_));
 sky130_fd_sc_hd__nand2_2 _22531_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[2][10] ),
    .Y(_09258_));
 sky130_fd_sc_hd__or2_2 _22532_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[2][10] ),
    .X(_09259_));
 sky130_fd_sc_hd__and2_2 _22533_ (.A(_09258_),
    .B(_09259_),
    .X(_09260_));
 sky130_fd_sc_hd__a21oi_2 _22534_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[2][9] ),
    .B1(_09256_),
    .Y(_09261_));
 sky130_fd_sc_hd__nand2_2 _22535_ (.A(_09255_),
    .B(_09261_),
    .Y(_09262_));
 sky130_fd_sc_hd__xor2_2 _22536_ (.A(_09260_),
    .B(_09262_),
    .X(_09263_));
 sky130_fd_sc_hd__a22o_2 _22537_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][10] ),
    .B1(_11712_),
    .B2(_09263_),
    .X(_01820_));
 sky130_fd_sc_hd__nor2_2 _22538_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[2][11] ),
    .Y(_09264_));
 sky130_fd_sc_hd__or2_2 _22539_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[2][11] ),
    .X(_09265_));
 sky130_fd_sc_hd__nand2_2 _22540_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[2][11] ),
    .Y(_09266_));
 sky130_fd_sc_hd__nand2_2 _22541_ (.A(_09265_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__a21bo_2 _22542_ (.A1(_09260_),
    .A2(_09262_),
    .B1_N(_09258_),
    .X(_09268_));
 sky130_fd_sc_hd__xnor2_2 _22543_ (.A(_09267_),
    .B(_09268_),
    .Y(_09269_));
 sky130_fd_sc_hd__a22o_2 _22544_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][11] ),
    .B1(_11712_),
    .B2(_09269_),
    .X(_01821_));
 sky130_fd_sc_hd__nand3_2 _22545_ (.A(_09260_),
    .B(_09265_),
    .C(_09266_),
    .Y(_09270_));
 sky130_fd_sc_hd__nor2_2 _22546_ (.A(_09254_),
    .B(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__o2bb2a_2 _22547_ (.A1_N(_09248_),
    .A2_N(_09271_),
    .B1(_09261_),
    .B2(_09270_),
    .X(_09272_));
 sky130_fd_sc_hd__o21a_2 _22548_ (.A1(_09258_),
    .A2(_09264_),
    .B1(_09266_),
    .X(_09273_));
 sky130_fd_sc_hd__xnor2_2 _22549_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[2][12] ),
    .Y(_09274_));
 sky130_fd_sc_hd__and3_2 _22550_ (.A(_09272_),
    .B(_09273_),
    .C(_09274_),
    .X(_09275_));
 sky130_fd_sc_hd__a21oi_2 _22551_ (.A1(_09272_),
    .A2(_09273_),
    .B1(_09274_),
    .Y(_09276_));
 sky130_fd_sc_hd__nor2_2 _22552_ (.A(_09275_),
    .B(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__a22o_2 _22553_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][12] ),
    .B1(_11712_),
    .B2(_09277_),
    .X(_01822_));
 sky130_fd_sc_hd__xor2_2 _22554_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[2][13] ),
    .X(_09278_));
 sky130_fd_sc_hd__a211o_2 _22555_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[2][12] ),
    .B1(_09276_),
    .C1(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__nand2b_2 _22556_ (.A_N(_09274_),
    .B(_09278_),
    .Y(_09280_));
 sky130_fd_sc_hd__a21o_2 _22557_ (.A1(_09272_),
    .A2(_09273_),
    .B1(_09280_),
    .X(_09281_));
 sky130_fd_sc_hd__and3_2 _22558_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[2][12] ),
    .C(_09278_),
    .X(_09282_));
 sky130_fd_sc_hd__nor2_2 _22559_ (.A(_11713_),
    .B(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__a32o_2 _22560_ (.A1(_09279_),
    .A2(_09281_),
    .A3(_09283_),
    .B1(\systolic_inst.acc_wires[2][13] ),
    .B2(_11258_),
    .X(_01823_));
 sky130_fd_sc_hd__or2_2 _22561_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[2][14] ),
    .X(_09284_));
 sky130_fd_sc_hd__nand2_2 _22562_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[2][14] ),
    .Y(_09285_));
 sky130_fd_sc_hd__and2_2 _22563_ (.A(_09284_),
    .B(_09285_),
    .X(_09286_));
 sky130_fd_sc_hd__a21oi_2 _22564_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[2][13] ),
    .B1(_09282_),
    .Y(_09287_));
 sky130_fd_sc_hd__nand2_2 _22565_ (.A(_09281_),
    .B(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__or2_2 _22566_ (.A(_09286_),
    .B(_09288_),
    .X(_09289_));
 sky130_fd_sc_hd__nand2_2 _22567_ (.A(_09286_),
    .B(_09288_),
    .Y(_09290_));
 sky130_fd_sc_hd__a32o_2 _22568_ (.A1(_11712_),
    .A2(_09289_),
    .A3(_09290_),
    .B1(\systolic_inst.acc_wires[2][14] ),
    .B2(_11258_),
    .X(_01824_));
 sky130_fd_sc_hd__nor2_2 _22569_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][15] ),
    .Y(_09291_));
 sky130_fd_sc_hd__and2_2 _22570_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][15] ),
    .X(_09292_));
 sky130_fd_sc_hd__a211o_2 _22571_ (.A1(_09285_),
    .A2(_09290_),
    .B1(_09291_),
    .C1(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__o211ai_2 _22572_ (.A1(_09291_),
    .A2(_09292_),
    .B1(_09285_),
    .C1(_09290_),
    .Y(_09294_));
 sky130_fd_sc_hd__a32o_2 _22573_ (.A1(_11712_),
    .A2(_09293_),
    .A3(_09294_),
    .B1(\systolic_inst.acc_wires[2][15] ),
    .B2(_11258_),
    .X(_01825_));
 sky130_fd_sc_hd__or3b_2 _22574_ (.A(_09291_),
    .B(_09292_),
    .C_N(_09286_),
    .X(_09295_));
 sky130_fd_sc_hd__a21o_2 _22575_ (.A1(_09281_),
    .A2(_09287_),
    .B1(_09295_),
    .X(_09296_));
 sky130_fd_sc_hd__o21ba_2 _22576_ (.A1(_09285_),
    .A2(_09291_),
    .B1_N(_09292_),
    .X(_09297_));
 sky130_fd_sc_hd__and2_2 _22577_ (.A(_09296_),
    .B(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__xnor2_2 _22578_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][16] ),
    .Y(_09299_));
 sky130_fd_sc_hd__nand2_2 _22579_ (.A(_09298_),
    .B(_09299_),
    .Y(_09300_));
 sky130_fd_sc_hd__nor2_2 _22580_ (.A(_09298_),
    .B(_09299_),
    .Y(_09301_));
 sky130_fd_sc_hd__nor2_2 _22581_ (.A(_11713_),
    .B(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__a22o_2 _22582_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][16] ),
    .B1(_09300_),
    .B2(_09302_),
    .X(_01826_));
 sky130_fd_sc_hd__xor2_2 _22583_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][17] ),
    .X(_09303_));
 sky130_fd_sc_hd__inv_2 _22584_ (.A(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__a21oi_2 _22585_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[2][16] ),
    .B1(_09301_),
    .Y(_09305_));
 sky130_fd_sc_hd__xnor2_2 _22586_ (.A(_09303_),
    .B(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__a22o_2 _22587_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][17] ),
    .B1(_11712_),
    .B2(_09306_),
    .X(_01827_));
 sky130_fd_sc_hd__or2_2 _22588_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][18] ),
    .X(_09307_));
 sky130_fd_sc_hd__nand2_2 _22589_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][18] ),
    .Y(_09308_));
 sky130_fd_sc_hd__nand2_2 _22590_ (.A(_09307_),
    .B(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__o21a_2 _22591_ (.A1(\systolic_inst.acc_wires[2][16] ),
    .A2(\systolic_inst.acc_wires[2][17] ),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .X(_09310_));
 sky130_fd_sc_hd__a21oi_2 _22592_ (.A1(_09301_),
    .A2(_09303_),
    .B1(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__xor2_2 _22593_ (.A(_09309_),
    .B(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__a22o_2 _22594_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][18] ),
    .B1(_11712_),
    .B2(_09312_),
    .X(_01828_));
 sky130_fd_sc_hd__xnor2_2 _22595_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][19] ),
    .Y(_09313_));
 sky130_fd_sc_hd__o21ai_2 _22596_ (.A1(_09309_),
    .A2(_09311_),
    .B1(_09308_),
    .Y(_09314_));
 sky130_fd_sc_hd__xnor2_2 _22597_ (.A(_09313_),
    .B(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__a22o_2 _22598_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][19] ),
    .B1(_11712_),
    .B2(_09315_),
    .X(_01829_));
 sky130_fd_sc_hd__xor2_2 _22599_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][20] ),
    .X(_09316_));
 sky130_fd_sc_hd__or4_2 _22600_ (.A(_09299_),
    .B(_09304_),
    .C(_09309_),
    .D(_09313_),
    .X(_09317_));
 sky130_fd_sc_hd__nor2_2 _22601_ (.A(_09298_),
    .B(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__o41a_2 _22602_ (.A1(\systolic_inst.acc_wires[2][16] ),
    .A2(\systolic_inst.acc_wires[2][17] ),
    .A3(\systolic_inst.acc_wires[2][18] ),
    .A4(\systolic_inst.acc_wires[2][19] ),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .X(_09319_));
 sky130_fd_sc_hd__or3_2 _22603_ (.A(_09316_),
    .B(_09318_),
    .C(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__o21ai_2 _22604_ (.A1(_09318_),
    .A2(_09319_),
    .B1(_09316_),
    .Y(_09321_));
 sky130_fd_sc_hd__a32o_2 _22605_ (.A1(_11712_),
    .A2(_09320_),
    .A3(_09321_),
    .B1(\systolic_inst.acc_wires[2][20] ),
    .B2(_11258_),
    .X(_01830_));
 sky130_fd_sc_hd__xor2_2 _22606_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][21] ),
    .X(_09322_));
 sky130_fd_sc_hd__a21bo_2 _22607_ (.A1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[2][20] ),
    .B1_N(_09321_),
    .X(_09323_));
 sky130_fd_sc_hd__xor2_2 _22608_ (.A(_09322_),
    .B(_09323_),
    .X(_09324_));
 sky130_fd_sc_hd__a22o_2 _22609_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][21] ),
    .B1(_11712_),
    .B2(_09324_),
    .X(_01831_));
 sky130_fd_sc_hd__or2_2 _22610_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][22] ),
    .X(_09325_));
 sky130_fd_sc_hd__nand2_2 _22611_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][22] ),
    .Y(_09326_));
 sky130_fd_sc_hd__and2_2 _22612_ (.A(_09325_),
    .B(_09326_),
    .X(_09327_));
 sky130_fd_sc_hd__o21a_2 _22613_ (.A1(\systolic_inst.acc_wires[2][20] ),
    .A2(\systolic_inst.acc_wires[2][21] ),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .X(_09328_));
 sky130_fd_sc_hd__and2b_2 _22614_ (.A_N(_09321_),
    .B(_09322_),
    .X(_09329_));
 sky130_fd_sc_hd__o21ai_2 _22615_ (.A1(_09328_),
    .A2(_09329_),
    .B1(_09327_),
    .Y(_09330_));
 sky130_fd_sc_hd__or3_2 _22616_ (.A(_09327_),
    .B(_09328_),
    .C(_09329_),
    .X(_09331_));
 sky130_fd_sc_hd__a32o_2 _22617_ (.A1(_11712_),
    .A2(_09330_),
    .A3(_09331_),
    .B1(\systolic_inst.acc_wires[2][22] ),
    .B2(_11258_),
    .X(_01832_));
 sky130_fd_sc_hd__xnor2_2 _22618_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][23] ),
    .Y(_09332_));
 sky130_fd_sc_hd__inv_2 _22619_ (.A(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__a21oi_2 _22620_ (.A1(_09326_),
    .A2(_09330_),
    .B1(_09332_),
    .Y(_09334_));
 sky130_fd_sc_hd__a31o_2 _22621_ (.A1(_09326_),
    .A2(_09330_),
    .A3(_09332_),
    .B1(_11713_),
    .X(_09335_));
 sky130_fd_sc_hd__a2bb2o_2 _22622_ (.A1_N(_09335_),
    .A2_N(_09334_),
    .B1(\systolic_inst.acc_wires[2][23] ),
    .B2(_11258_),
    .X(_01833_));
 sky130_fd_sc_hd__nand4_2 _22623_ (.A(_09316_),
    .B(_09322_),
    .C(_09327_),
    .D(_09333_),
    .Y(_09336_));
 sky130_fd_sc_hd__a211o_2 _22624_ (.A1(_09296_),
    .A2(_09297_),
    .B1(_09317_),
    .C1(_09336_),
    .X(_09337_));
 sky130_fd_sc_hd__o41a_2 _22625_ (.A1(\systolic_inst.acc_wires[2][20] ),
    .A2(\systolic_inst.acc_wires[2][21] ),
    .A3(\systolic_inst.acc_wires[2][22] ),
    .A4(\systolic_inst.acc_wires[2][23] ),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .X(_09338_));
 sky130_fd_sc_hd__nor2_2 _22626_ (.A(_09319_),
    .B(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__nor2_2 _22627_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][24] ),
    .Y(_09340_));
 sky130_fd_sc_hd__and2_2 _22628_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][24] ),
    .X(_09341_));
 sky130_fd_sc_hd__or2_2 _22629_ (.A(_09340_),
    .B(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__a21oi_2 _22630_ (.A1(_09337_),
    .A2(_09339_),
    .B1(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__a31o_2 _22631_ (.A1(_09337_),
    .A2(_09339_),
    .A3(_09342_),
    .B1(_11713_),
    .X(_09344_));
 sky130_fd_sc_hd__a2bb2o_2 _22632_ (.A1_N(_09344_),
    .A2_N(_09343_),
    .B1(\systolic_inst.acc_wires[2][24] ),
    .B2(_11258_),
    .X(_01834_));
 sky130_fd_sc_hd__xor2_2 _22633_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][25] ),
    .X(_09345_));
 sky130_fd_sc_hd__or3_2 _22634_ (.A(_09341_),
    .B(_09343_),
    .C(_09345_),
    .X(_09346_));
 sky130_fd_sc_hd__o21ai_2 _22635_ (.A1(_09341_),
    .A2(_09343_),
    .B1(_09345_),
    .Y(_09347_));
 sky130_fd_sc_hd__a32o_2 _22636_ (.A1(_11712_),
    .A2(_09346_),
    .A3(_09347_),
    .B1(\systolic_inst.acc_wires[2][25] ),
    .B2(_11258_),
    .X(_01835_));
 sky130_fd_sc_hd__or2_2 _22637_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][26] ),
    .X(_09348_));
 sky130_fd_sc_hd__nand2_2 _22638_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][26] ),
    .Y(_09349_));
 sky130_fd_sc_hd__nand2_2 _22639_ (.A(_09348_),
    .B(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__o21a_2 _22640_ (.A1(\systolic_inst.acc_wires[2][24] ),
    .A2(\systolic_inst.acc_wires[2][25] ),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .X(_09351_));
 sky130_fd_sc_hd__a21o_2 _22641_ (.A1(_09343_),
    .A2(_09345_),
    .B1(_09351_),
    .X(_09352_));
 sky130_fd_sc_hd__xnor2_2 _22642_ (.A(_09350_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__a22o_2 _22643_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][26] ),
    .B1(_11712_),
    .B2(_09353_),
    .X(_01836_));
 sky130_fd_sc_hd__xnor2_2 _22644_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][27] ),
    .Y(_09354_));
 sky130_fd_sc_hd__a21bo_2 _22645_ (.A1(_09348_),
    .A2(_09352_),
    .B1_N(_09349_),
    .X(_09355_));
 sky130_fd_sc_hd__xnor2_2 _22646_ (.A(_09354_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__a22o_2 _22647_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][27] ),
    .B1(_11712_),
    .B2(_09356_),
    .X(_01837_));
 sky130_fd_sc_hd__nor2_2 _22648_ (.A(_09350_),
    .B(_09354_),
    .Y(_09357_));
 sky130_fd_sc_hd__o21a_2 _22649_ (.A1(\systolic_inst.acc_wires[2][26] ),
    .A2(\systolic_inst.acc_wires[2][27] ),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .X(_09358_));
 sky130_fd_sc_hd__a311oi_2 _22650_ (.A1(_09343_),
    .A2(_09345_),
    .A3(_09357_),
    .B1(_09358_),
    .C1(_09351_),
    .Y(_09359_));
 sky130_fd_sc_hd__or2_2 _22651_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][28] ),
    .X(_09360_));
 sky130_fd_sc_hd__nand2_2 _22652_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][28] ),
    .Y(_09361_));
 sky130_fd_sc_hd__nand2_2 _22653_ (.A(_09360_),
    .B(_09361_),
    .Y(_09362_));
 sky130_fd_sc_hd__xor2_2 _22654_ (.A(_09359_),
    .B(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__a22o_2 _22655_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][28] ),
    .B1(_11712_),
    .B2(_09363_),
    .X(_01838_));
 sky130_fd_sc_hd__xor2_2 _22656_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][29] ),
    .X(_09364_));
 sky130_fd_sc_hd__inv_2 _22657_ (.A(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__o21a_2 _22658_ (.A1(_09359_),
    .A2(_09362_),
    .B1(_09361_),
    .X(_09366_));
 sky130_fd_sc_hd__xnor2_2 _22659_ (.A(_09364_),
    .B(_09366_),
    .Y(_09367_));
 sky130_fd_sc_hd__a22o_2 _22660_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[2][29] ),
    .B1(_11712_),
    .B2(_09367_),
    .X(_01839_));
 sky130_fd_sc_hd__o21ai_2 _22661_ (.A1(\systolic_inst.acc_wires[2][28] ),
    .A2(\systolic_inst.acc_wires[2][29] ),
    .B1(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .Y(_09368_));
 sky130_fd_sc_hd__o31a_2 _22662_ (.A1(_09359_),
    .A2(_09362_),
    .A3(_09365_),
    .B1(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__nand2_2 _22663_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][30] ),
    .Y(_09370_));
 sky130_fd_sc_hd__or2_2 _22664_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][30] ),
    .X(_09371_));
 sky130_fd_sc_hd__nand2_2 _22665_ (.A(_09370_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__nand2_2 _22666_ (.A(_09369_),
    .B(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__or2_2 _22667_ (.A(_09369_),
    .B(_09372_),
    .X(_09374_));
 sky130_fd_sc_hd__a32o_2 _22668_ (.A1(_11712_),
    .A2(_09373_),
    .A3(_09374_),
    .B1(\systolic_inst.acc_wires[2][30] ),
    .B2(_11258_),
    .X(_01840_));
 sky130_fd_sc_hd__xnor2_2 _22669_ (.A(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[2][31] ),
    .Y(_09375_));
 sky130_fd_sc_hd__a21oi_2 _22670_ (.A1(_09370_),
    .A2(_09374_),
    .B1(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__a31o_2 _22671_ (.A1(_09370_),
    .A2(_09374_),
    .A3(_09375_),
    .B1(_11713_),
    .X(_09377_));
 sky130_fd_sc_hd__a2bb2o_2 _22672_ (.A1_N(_09377_),
    .A2_N(_09376_),
    .B1(\systolic_inst.acc_wires[2][31] ),
    .B2(_11258_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _22673_ (.A0(\systolic_inst.A_outs[1][0] ),
    .A1(\systolic_inst.A_outs[0][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _22674_ (.A0(\systolic_inst.A_outs[1][1] ),
    .A1(\systolic_inst.A_outs[0][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _22675_ (.A0(\systolic_inst.A_outs[1][2] ),
    .A1(\systolic_inst.A_outs[0][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _22676_ (.A0(\systolic_inst.A_outs[1][3] ),
    .A1(\systolic_inst.A_outs[0][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _22677_ (.A0(\systolic_inst.A_outs[1][4] ),
    .A1(\systolic_inst.A_outs[0][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _22678_ (.A0(\systolic_inst.A_outs[1][5] ),
    .A1(\systolic_inst.A_outs[0][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _22679_ (.A0(\systolic_inst.A_outs[1][6] ),
    .A1(\systolic_inst.A_outs[0][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _22680_ (.A0(\systolic_inst.A_outs[1][7] ),
    .A1(\systolic_inst.A_outs[0][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _22681_ (.A0(\systolic_inst.B_outs[0][0] ),
    .A1(\systolic_inst.B_shift[0][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _22682_ (.A0(\systolic_inst.B_outs[0][1] ),
    .A1(\systolic_inst.B_shift[0][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _22683_ (.A0(\systolic_inst.B_outs[0][2] ),
    .A1(\systolic_inst.B_shift[0][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _22684_ (.A0(\systolic_inst.B_outs[0][3] ),
    .A1(\systolic_inst.B_shift[0][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _22685_ (.A0(\systolic_inst.B_outs[0][4] ),
    .A1(\systolic_inst.B_shift[0][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _22686_ (.A0(\systolic_inst.B_outs[0][5] ),
    .A1(\systolic_inst.B_shift[0][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _22687_ (.A0(\systolic_inst.B_outs[0][6] ),
    .A1(\systolic_inst.B_shift[0][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _22688_ (.A0(\systolic_inst.B_outs[0][7] ),
    .A1(\systolic_inst.B_shift[0][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01857_));
 sky130_fd_sc_hd__and3_2 _22689_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[1][0] ),
    .C(\systolic_inst.A_outs[1][0] ),
    .X(_09378_));
 sky130_fd_sc_hd__a21o_2 _22690_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[0] ),
    .B1(_09378_),
    .X(_01858_));
 sky130_fd_sc_hd__and4_2 _22691_ (.A(\systolic_inst.B_outs[1][0] ),
    .B(\systolic_inst.A_outs[1][0] ),
    .C(\systolic_inst.B_outs[1][1] ),
    .D(\systolic_inst.A_outs[1][1] ),
    .X(_09379_));
 sky130_fd_sc_hd__a22o_2 _22692_ (.A1(\systolic_inst.A_outs[1][0] ),
    .A2(\systolic_inst.B_outs[1][1] ),
    .B1(\systolic_inst.A_outs[1][1] ),
    .B2(\systolic_inst.B_outs[1][0] ),
    .X(_09380_));
 sky130_fd_sc_hd__nand2_2 _22693_ (.A(\systolic_inst.ce_local ),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__a2bb2o_2 _22694_ (.A1_N(_09381_),
    .A2_N(_09379_),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01859_));
 sky130_fd_sc_hd__and2_2 _22695_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[2] ),
    .X(_09382_));
 sky130_fd_sc_hd__a22oi_2 _22696_ (.A1(\systolic_inst.B_outs[1][1] ),
    .A2(\systolic_inst.A_outs[1][1] ),
    .B1(\systolic_inst.A_outs[1][2] ),
    .B2(\systolic_inst.B_outs[1][0] ),
    .Y(_09383_));
 sky130_fd_sc_hd__and4_2 _22697_ (.A(\systolic_inst.B_outs[1][0] ),
    .B(\systolic_inst.B_outs[1][1] ),
    .C(\systolic_inst.A_outs[1][1] ),
    .D(\systolic_inst.A_outs[1][2] ),
    .X(_09384_));
 sky130_fd_sc_hd__or2_2 _22698_ (.A(_09383_),
    .B(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__or3b_2 _22699_ (.A(_09383_),
    .B(_09384_),
    .C_N(_09379_),
    .X(_09386_));
 sky130_fd_sc_hd__xnor2_2 _22700_ (.A(_09379_),
    .B(_09385_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand3_2 _22701_ (.A(\systolic_inst.A_outs[1][0] ),
    .B(\systolic_inst.B_outs[1][2] ),
    .C(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__a21o_2 _22702_ (.A1(\systolic_inst.A_outs[1][0] ),
    .A2(\systolic_inst.B_outs[1][2] ),
    .B1(_09387_),
    .X(_09389_));
 sky130_fd_sc_hd__a31o_2 _22703_ (.A1(\systolic_inst.ce_local ),
    .A2(_09388_),
    .A3(_09389_),
    .B1(_09382_),
    .X(_01860_));
 sky130_fd_sc_hd__a22oi_2 _22704_ (.A1(\systolic_inst.A_outs[1][1] ),
    .A2(\systolic_inst.B_outs[1][2] ),
    .B1(\systolic_inst.B_outs[1][3] ),
    .B2(\systolic_inst.A_outs[1][0] ),
    .Y(_09390_));
 sky130_fd_sc_hd__and4_2 _22705_ (.A(\systolic_inst.A_outs[1][0] ),
    .B(\systolic_inst.A_outs[1][1] ),
    .C(\systolic_inst.B_outs[1][2] ),
    .D(\systolic_inst.B_outs[1][3] ),
    .X(_09391_));
 sky130_fd_sc_hd__nor2_2 _22706_ (.A(_09390_),
    .B(_09391_),
    .Y(_09392_));
 sky130_fd_sc_hd__nand4_2 _22707_ (.A(\systolic_inst.B_outs[1][0] ),
    .B(\systolic_inst.B_outs[1][1] ),
    .C(\systolic_inst.A_outs[1][2] ),
    .D(\systolic_inst.A_outs[1][3] ),
    .Y(_09393_));
 sky130_fd_sc_hd__a22o_2 _22708_ (.A1(\systolic_inst.B_outs[1][1] ),
    .A2(\systolic_inst.A_outs[1][2] ),
    .B1(\systolic_inst.A_outs[1][3] ),
    .B2(\systolic_inst.B_outs[1][0] ),
    .X(_09394_));
 sky130_fd_sc_hd__nand3_2 _22709_ (.A(_09384_),
    .B(_09393_),
    .C(_09394_),
    .Y(_09395_));
 sky130_fd_sc_hd__a21o_2 _22710_ (.A1(_09393_),
    .A2(_09394_),
    .B1(_09384_),
    .X(_09396_));
 sky130_fd_sc_hd__and2_2 _22711_ (.A(_09395_),
    .B(_09396_),
    .X(_09397_));
 sky130_fd_sc_hd__nand2_2 _22712_ (.A(_09392_),
    .B(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__xnor2_2 _22713_ (.A(_09392_),
    .B(_09397_),
    .Y(_09399_));
 sky130_fd_sc_hd__and3_2 _22714_ (.A(_09386_),
    .B(_09388_),
    .C(_09399_),
    .X(_09400_));
 sky130_fd_sc_hd__a21oi_2 _22715_ (.A1(_09386_),
    .A2(_09388_),
    .B1(_09399_),
    .Y(_09401_));
 sky130_fd_sc_hd__nand2_2 _22716_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[3] ),
    .Y(_09402_));
 sky130_fd_sc_hd__o31ai_2 _22717_ (.A1(_11258_),
    .A2(_09400_),
    .A3(_09401_),
    .B1(_09402_),
    .Y(_01861_));
 sky130_fd_sc_hd__and2_2 _22718_ (.A(\systolic_inst.B_outs[1][2] ),
    .B(\systolic_inst.A_outs[1][2] ),
    .X(_09403_));
 sky130_fd_sc_hd__nand4_2 _22719_ (.A(\systolic_inst.A_outs[1][0] ),
    .B(\systolic_inst.A_outs[1][1] ),
    .C(\systolic_inst.B_outs[1][3] ),
    .D(\systolic_inst.B_outs[1][4] ),
    .Y(_09404_));
 sky130_fd_sc_hd__a22o_2 _22720_ (.A1(\systolic_inst.A_outs[1][1] ),
    .A2(\systolic_inst.B_outs[1][3] ),
    .B1(\systolic_inst.B_outs[1][4] ),
    .B2(\systolic_inst.A_outs[1][0] ),
    .X(_09405_));
 sky130_fd_sc_hd__nand2_2 _22721_ (.A(_09404_),
    .B(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__xnor2_2 _22722_ (.A(_09403_),
    .B(_09406_),
    .Y(_09407_));
 sky130_fd_sc_hd__a22o_2 _22723_ (.A1(\systolic_inst.B_outs[1][1] ),
    .A2(\systolic_inst.A_outs[1][3] ),
    .B1(\systolic_inst.A_outs[1][4] ),
    .B2(\systolic_inst.B_outs[1][0] ),
    .X(_09408_));
 sky130_fd_sc_hd__and3_2 _22724_ (.A(\systolic_inst.B_outs[1][0] ),
    .B(\systolic_inst.B_outs[1][1] ),
    .C(\systolic_inst.A_outs[1][3] ),
    .X(_09409_));
 sky130_fd_sc_hd__nand2_2 _22725_ (.A(\systolic_inst.A_outs[1][4] ),
    .B(_09409_),
    .Y(_09410_));
 sky130_fd_sc_hd__and3_2 _22726_ (.A(_09391_),
    .B(_09408_),
    .C(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__a21oi_2 _22727_ (.A1(_09408_),
    .A2(_09410_),
    .B1(_09391_),
    .Y(_09412_));
 sky130_fd_sc_hd__o21ai_2 _22728_ (.A1(_09411_),
    .A2(_09412_),
    .B1(_09393_),
    .Y(_09413_));
 sky130_fd_sc_hd__nor3_2 _22729_ (.A(_09393_),
    .B(_09411_),
    .C(_09412_),
    .Y(_09414_));
 sky130_fd_sc_hd__or3_2 _22730_ (.A(_09393_),
    .B(_09411_),
    .C(_09412_),
    .X(_09415_));
 sky130_fd_sc_hd__and3_2 _22731_ (.A(_09407_),
    .B(_09413_),
    .C(_09415_),
    .X(_09416_));
 sky130_fd_sc_hd__a21oi_2 _22732_ (.A1(_09413_),
    .A2(_09415_),
    .B1(_09407_),
    .Y(_09417_));
 sky130_fd_sc_hd__a211o_2 _22733_ (.A1(_09395_),
    .A2(_09398_),
    .B1(_09416_),
    .C1(_09417_),
    .X(_09418_));
 sky130_fd_sc_hd__o211ai_2 _22734_ (.A1(_09416_),
    .A2(_09417_),
    .B1(_09395_),
    .C1(_09398_),
    .Y(_09419_));
 sky130_fd_sc_hd__a21oi_2 _22735_ (.A1(_09418_),
    .A2(_09419_),
    .B1(_09401_),
    .Y(_09420_));
 sky130_fd_sc_hd__a31o_2 _22736_ (.A1(_09401_),
    .A2(_09418_),
    .A3(_09419_),
    .B1(_11258_),
    .X(_09421_));
 sky130_fd_sc_hd__a2bb2o_2 _22737_ (.A1_N(_09421_),
    .A2_N(_09420_),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[4] ),
    .B2(_11258_),
    .X(_01862_));
 sky130_fd_sc_hd__a21bo_2 _22738_ (.A1(_09403_),
    .A2(_09405_),
    .B1_N(_09404_),
    .X(_09422_));
 sky130_fd_sc_hd__a22oi_2 _22739_ (.A1(\systolic_inst.B_outs[1][1] ),
    .A2(\systolic_inst.A_outs[1][4] ),
    .B1(\systolic_inst.A_outs[1][5] ),
    .B2(\systolic_inst.B_outs[1][0] ),
    .Y(_09423_));
 sky130_fd_sc_hd__and4_2 _22740_ (.A(\systolic_inst.B_outs[1][0] ),
    .B(\systolic_inst.B_outs[1][1] ),
    .C(\systolic_inst.A_outs[1][4] ),
    .D(\systolic_inst.A_outs[1][5] ),
    .X(_09424_));
 sky130_fd_sc_hd__nor2_2 _22741_ (.A(_09423_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__xor2_2 _22742_ (.A(_09422_),
    .B(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__xor2_2 _22743_ (.A(_09410_),
    .B(_09426_),
    .X(_09427_));
 sky130_fd_sc_hd__and2_2 _22744_ (.A(\systolic_inst.A_outs[1][0] ),
    .B(\systolic_inst.B_outs[1][5] ),
    .X(_09428_));
 sky130_fd_sc_hd__nand2_2 _22745_ (.A(\systolic_inst.A_outs[1][0] ),
    .B(\systolic_inst.B_outs[1][5] ),
    .Y(_09429_));
 sky130_fd_sc_hd__nand2_2 _22746_ (.A(\systolic_inst.B_outs[1][2] ),
    .B(\systolic_inst.A_outs[1][3] ),
    .Y(_09430_));
 sky130_fd_sc_hd__and4_2 _22747_ (.A(\systolic_inst.A_outs[1][1] ),
    .B(\systolic_inst.A_outs[1][2] ),
    .C(\systolic_inst.B_outs[1][3] ),
    .D(\systolic_inst.B_outs[1][4] ),
    .X(_09431_));
 sky130_fd_sc_hd__a22oi_2 _22748_ (.A1(\systolic_inst.A_outs[1][2] ),
    .A2(\systolic_inst.B_outs[1][3] ),
    .B1(\systolic_inst.B_outs[1][4] ),
    .B2(\systolic_inst.A_outs[1][1] ),
    .Y(_09432_));
 sky130_fd_sc_hd__or3_2 _22749_ (.A(_09430_),
    .B(_09431_),
    .C(_09432_),
    .X(_09433_));
 sky130_fd_sc_hd__o21ai_2 _22750_ (.A1(_09431_),
    .A2(_09432_),
    .B1(_09430_),
    .Y(_09434_));
 sky130_fd_sc_hd__and3_2 _22751_ (.A(_09428_),
    .B(_09433_),
    .C(_09434_),
    .X(_09435_));
 sky130_fd_sc_hd__a21oi_2 _22752_ (.A1(_09433_),
    .A2(_09434_),
    .B1(_09428_),
    .Y(_09436_));
 sky130_fd_sc_hd__or2_2 _22753_ (.A(_09435_),
    .B(_09436_),
    .X(_09437_));
 sky130_fd_sc_hd__nor2_2 _22754_ (.A(_09427_),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__xor2_2 _22755_ (.A(_09427_),
    .B(_09437_),
    .X(_09439_));
 sky130_fd_sc_hd__and2_2 _22756_ (.A(_09416_),
    .B(_09439_),
    .X(_09440_));
 sky130_fd_sc_hd__xor2_2 _22757_ (.A(_09416_),
    .B(_09439_),
    .X(_09441_));
 sky130_fd_sc_hd__o21a_2 _22758_ (.A1(_09411_),
    .A2(_09414_),
    .B1(_09441_),
    .X(_09442_));
 sky130_fd_sc_hd__nor3_2 _22759_ (.A(_09411_),
    .B(_09414_),
    .C(_09441_),
    .Y(_09443_));
 sky130_fd_sc_hd__nor2_2 _22760_ (.A(_09442_),
    .B(_09443_),
    .Y(_09444_));
 sky130_fd_sc_hd__a21bo_2 _22761_ (.A1(_09401_),
    .A2(_09419_),
    .B1_N(_09418_),
    .X(_09445_));
 sky130_fd_sc_hd__nand2_2 _22762_ (.A(_09444_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__o21a_2 _22763_ (.A1(_09444_),
    .A2(_09445_),
    .B1(\systolic_inst.ce_local ),
    .X(_09447_));
 sky130_fd_sc_hd__a22o_2 _22764_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[5] ),
    .B1(_09446_),
    .B2(_09447_),
    .X(_01863_));
 sky130_fd_sc_hd__a32o_2 _22765_ (.A1(\systolic_inst.A_outs[1][4] ),
    .A2(_09409_),
    .A3(_09426_),
    .B1(_09425_),
    .B2(_09422_),
    .X(_09448_));
 sky130_fd_sc_hd__o21bai_2 _22766_ (.A1(_09430_),
    .A2(_09432_),
    .B1_N(_09431_),
    .Y(_09449_));
 sky130_fd_sc_hd__a22oi_2 _22767_ (.A1(\systolic_inst.B_outs[1][1] ),
    .A2(\systolic_inst.A_outs[1][5] ),
    .B1(\systolic_inst.A_outs[1][6] ),
    .B2(\systolic_inst.B_outs[1][0] ),
    .Y(_09450_));
 sky130_fd_sc_hd__and4_2 _22768_ (.A(\systolic_inst.B_outs[1][0] ),
    .B(\systolic_inst.B_outs[1][1] ),
    .C(\systolic_inst.A_outs[1][5] ),
    .D(\systolic_inst.A_outs[1][6] ),
    .X(_09451_));
 sky130_fd_sc_hd__or2_2 _22769_ (.A(_09450_),
    .B(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__nand2b_2 _22770_ (.A_N(_09452_),
    .B(_09449_),
    .Y(_09453_));
 sky130_fd_sc_hd__xnor2_2 _22771_ (.A(_09449_),
    .B(_09452_),
    .Y(_09454_));
 sky130_fd_sc_hd__nand2_2 _22772_ (.A(_09424_),
    .B(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__xor2_2 _22773_ (.A(_09424_),
    .B(_09454_),
    .X(_09456_));
 sky130_fd_sc_hd__nand4_2 _22774_ (.A(\systolic_inst.A_outs[1][2] ),
    .B(\systolic_inst.B_outs[1][3] ),
    .C(\systolic_inst.A_outs[1][3] ),
    .D(\systolic_inst.B_outs[1][4] ),
    .Y(_09457_));
 sky130_fd_sc_hd__a22o_2 _22775_ (.A1(\systolic_inst.B_outs[1][3] ),
    .A2(\systolic_inst.A_outs[1][3] ),
    .B1(\systolic_inst.B_outs[1][4] ),
    .B2(\systolic_inst.A_outs[1][2] ),
    .X(_09458_));
 sky130_fd_sc_hd__nand4_2 _22776_ (.A(\systolic_inst.B_outs[1][2] ),
    .B(\systolic_inst.A_outs[1][4] ),
    .C(_09457_),
    .D(_09458_),
    .Y(_09459_));
 sky130_fd_sc_hd__a22o_2 _22777_ (.A1(\systolic_inst.B_outs[1][2] ),
    .A2(\systolic_inst.A_outs[1][4] ),
    .B1(_09457_),
    .B2(_09458_),
    .X(_09460_));
 sky130_fd_sc_hd__nand2_2 _22778_ (.A(\systolic_inst.A_outs[1][1] ),
    .B(\systolic_inst.B_outs[1][6] ),
    .Y(_09461_));
 sky130_fd_sc_hd__a22o_2 _22779_ (.A1(\systolic_inst.A_outs[1][1] ),
    .A2(\systolic_inst.B_outs[1][5] ),
    .B1(\systolic_inst.B_outs[1][6] ),
    .B2(\systolic_inst.A_outs[1][0] ),
    .X(_09462_));
 sky130_fd_sc_hd__o21a_2 _22780_ (.A1(_09429_),
    .A2(_09461_),
    .B1(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__nand3_2 _22781_ (.A(_09459_),
    .B(_09460_),
    .C(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__a21o_2 _22782_ (.A1(_09459_),
    .A2(_09460_),
    .B1(_09463_),
    .X(_09465_));
 sky130_fd_sc_hd__nand3_2 _22783_ (.A(_09435_),
    .B(_09464_),
    .C(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__a21o_2 _22784_ (.A1(_09464_),
    .A2(_09465_),
    .B1(_09435_),
    .X(_09467_));
 sky130_fd_sc_hd__nand3_2 _22785_ (.A(_09456_),
    .B(_09466_),
    .C(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__a21o_2 _22786_ (.A1(_09466_),
    .A2(_09467_),
    .B1(_09456_),
    .X(_09469_));
 sky130_fd_sc_hd__nand3_2 _22787_ (.A(_09438_),
    .B(_09468_),
    .C(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__a21o_2 _22788_ (.A1(_09468_),
    .A2(_09469_),
    .B1(_09438_),
    .X(_09471_));
 sky130_fd_sc_hd__nand3_2 _22789_ (.A(_09448_),
    .B(_09470_),
    .C(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__a21o_2 _22790_ (.A1(_09470_),
    .A2(_09471_),
    .B1(_09448_),
    .X(_09473_));
 sky130_fd_sc_hd__o211a_2 _22791_ (.A1(_09440_),
    .A2(_09442_),
    .B1(_09472_),
    .C1(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__a211o_2 _22792_ (.A1(_09472_),
    .A2(_09473_),
    .B1(_09440_),
    .C1(_09442_),
    .X(_09475_));
 sky130_fd_sc_hd__and2b_2 _22793_ (.A_N(_09474_),
    .B(_09475_),
    .X(_09476_));
 sky130_fd_sc_hd__xnor2_2 _22794_ (.A(_09446_),
    .B(_09476_),
    .Y(_09477_));
 sky130_fd_sc_hd__mux2_1 _22795_ (.A0(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[6] ),
    .A1(_09477_),
    .S(\systolic_inst.ce_local ),
    .X(_01864_));
 sky130_fd_sc_hd__nand2_2 _22796_ (.A(_09457_),
    .B(_09459_),
    .Y(_09478_));
 sky130_fd_sc_hd__nand2_2 _22797_ (.A(\systolic_inst.B_outs[1][0] ),
    .B(\systolic_inst.A_outs[1][7] ),
    .Y(_09479_));
 sky130_fd_sc_hd__nand2_2 _22798_ (.A(\systolic_inst.B_outs[1][2] ),
    .B(\systolic_inst.A_outs[1][6] ),
    .Y(_09480_));
 sky130_fd_sc_hd__and4_2 _22799_ (.A(\systolic_inst.B_outs[1][1] ),
    .B(\systolic_inst.B_outs[1][2] ),
    .C(\systolic_inst.A_outs[1][5] ),
    .D(\systolic_inst.A_outs[1][6] ),
    .X(_09481_));
 sky130_fd_sc_hd__a22o_2 _22800_ (.A1(\systolic_inst.B_outs[1][2] ),
    .A2(\systolic_inst.A_outs[1][5] ),
    .B1(\systolic_inst.A_outs[1][6] ),
    .B2(\systolic_inst.B_outs[1][1] ),
    .X(_09482_));
 sky130_fd_sc_hd__and2b_2 _22801_ (.A_N(_09481_),
    .B(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__xnor2_2 _22802_ (.A(_09479_),
    .B(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__and2_2 _22803_ (.A(_09478_),
    .B(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__xor2_2 _22804_ (.A(_09478_),
    .B(_09484_),
    .X(_09486_));
 sky130_fd_sc_hd__xnor2_2 _22805_ (.A(_09451_),
    .B(_09486_),
    .Y(_09487_));
 sky130_fd_sc_hd__nand2_2 _22806_ (.A(\systolic_inst.B_outs[1][3] ),
    .B(\systolic_inst.A_outs[1][4] ),
    .Y(_09488_));
 sky130_fd_sc_hd__nand2_2 _22807_ (.A(\systolic_inst.A_outs[1][3] ),
    .B(\systolic_inst.B_outs[1][5] ),
    .Y(_09489_));
 sky130_fd_sc_hd__and4_2 _22808_ (.A(\systolic_inst.A_outs[1][2] ),
    .B(\systolic_inst.A_outs[1][3] ),
    .C(\systolic_inst.B_outs[1][4] ),
    .D(\systolic_inst.B_outs[1][5] ),
    .X(_09490_));
 sky130_fd_sc_hd__a22o_2 _22809_ (.A1(\systolic_inst.A_outs[1][3] ),
    .A2(\systolic_inst.B_outs[1][4] ),
    .B1(\systolic_inst.B_outs[1][5] ),
    .B2(\systolic_inst.A_outs[1][2] ),
    .X(_09491_));
 sky130_fd_sc_hd__and2b_2 _22810_ (.A_N(_09490_),
    .B(_09491_),
    .X(_09492_));
 sky130_fd_sc_hd__xnor2_2 _22811_ (.A(_09488_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__a2bb2o_2 _22812_ (.A1_N(_09428_),
    .A2_N(_09461_),
    .B1(\systolic_inst.A_outs[1][0] ),
    .B2(\systolic_inst.B_outs[1][7] ),
    .X(_09494_));
 sky130_fd_sc_hd__or4b_2 _22813_ (.A(\systolic_inst.B_outs[1][5] ),
    .B(_11277_),
    .C(_09461_),
    .D_N(\systolic_inst.A_outs[1][0] ),
    .X(_09495_));
 sky130_fd_sc_hd__and2_2 _22814_ (.A(_09494_),
    .B(_09495_),
    .X(_09496_));
 sky130_fd_sc_hd__nand2_2 _22815_ (.A(_09493_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__xnor2_2 _22816_ (.A(_09493_),
    .B(_09496_),
    .Y(_09498_));
 sky130_fd_sc_hd__xnor2_2 _22817_ (.A(_09464_),
    .B(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__or2_2 _22818_ (.A(_09487_),
    .B(_09499_),
    .X(_09500_));
 sky130_fd_sc_hd__nand2_2 _22819_ (.A(_09487_),
    .B(_09499_),
    .Y(_09501_));
 sky130_fd_sc_hd__nand2_2 _22820_ (.A(_09466_),
    .B(_09468_),
    .Y(_09502_));
 sky130_fd_sc_hd__and3_2 _22821_ (.A(_09500_),
    .B(_09501_),
    .C(_09502_),
    .X(_09503_));
 sky130_fd_sc_hd__a21oi_2 _22822_ (.A1(_09500_),
    .A2(_09501_),
    .B1(_09502_),
    .Y(_09504_));
 sky130_fd_sc_hd__a211oi_2 _22823_ (.A1(_09453_),
    .A2(_09455_),
    .B1(_09503_),
    .C1(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__o211a_2 _22824_ (.A1(_09503_),
    .A2(_09504_),
    .B1(_09453_),
    .C1(_09455_),
    .X(_09506_));
 sky130_fd_sc_hd__a211oi_2 _22825_ (.A1(_09470_),
    .A2(_09472_),
    .B1(_09505_),
    .C1(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__o211ai_2 _22826_ (.A1(_09505_),
    .A2(_09506_),
    .B1(_09470_),
    .C1(_09472_),
    .Y(_09508_));
 sky130_fd_sc_hd__nand2b_2 _22827_ (.A_N(_09507_),
    .B(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__a31o_2 _22828_ (.A1(_09444_),
    .A2(_09445_),
    .A3(_09475_),
    .B1(_09474_),
    .X(_09510_));
 sky130_fd_sc_hd__xnor2_2 _22829_ (.A(_09509_),
    .B(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__mux2_1 _22830_ (.A0(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[7] ),
    .A1(_09511_),
    .S(\systolic_inst.ce_local ),
    .X(_01865_));
 sky130_fd_sc_hd__a21oi_2 _22831_ (.A1(_09451_),
    .A2(_09486_),
    .B1(_09485_),
    .Y(_09512_));
 sky130_fd_sc_hd__a31o_2 _22832_ (.A1(\systolic_inst.B_outs[1][0] ),
    .A2(\systolic_inst.A_outs[1][7] ),
    .A3(_09482_),
    .B1(_09481_),
    .X(_09513_));
 sky130_fd_sc_hd__a31o_2 _22833_ (.A1(\systolic_inst.B_outs[1][3] ),
    .A2(\systolic_inst.A_outs[1][4] ),
    .A3(_09491_),
    .B1(_09490_),
    .X(_09514_));
 sky130_fd_sc_hd__o21ai_2 _22834_ (.A1(\systolic_inst.B_outs[1][0] ),
    .A2(\systolic_inst.B_outs[1][1] ),
    .B1(\systolic_inst.A_outs[1][7] ),
    .Y(_09515_));
 sky130_fd_sc_hd__o21a_2 _22835_ (.A1(\systolic_inst.B_outs[1][0] ),
    .A2(\systolic_inst.B_outs[1][1] ),
    .B1(\systolic_inst.A_outs[1][7] ),
    .X(_09516_));
 sky130_fd_sc_hd__a21o_2 _22836_ (.A1(\systolic_inst.B_outs[1][0] ),
    .A2(\systolic_inst.B_outs[1][1] ),
    .B1(_09515_),
    .X(_09517_));
 sky130_fd_sc_hd__and2b_2 _22837_ (.A_N(_09517_),
    .B(_09514_),
    .X(_09518_));
 sky130_fd_sc_hd__xnor2_2 _22838_ (.A(_09514_),
    .B(_09517_),
    .Y(_09519_));
 sky130_fd_sc_hd__xnor2_2 _22839_ (.A(_09513_),
    .B(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__and4_2 _22840_ (.A(\systolic_inst.B_outs[1][3] ),
    .B(\systolic_inst.B_outs[1][4] ),
    .C(\systolic_inst.A_outs[1][4] ),
    .D(\systolic_inst.A_outs[1][5] ),
    .X(_09521_));
 sky130_fd_sc_hd__a22oi_2 _22841_ (.A1(\systolic_inst.B_outs[1][4] ),
    .A2(\systolic_inst.A_outs[1][4] ),
    .B1(\systolic_inst.A_outs[1][5] ),
    .B2(\systolic_inst.B_outs[1][3] ),
    .Y(_09522_));
 sky130_fd_sc_hd__nor2_2 _22842_ (.A(_09521_),
    .B(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__xnor2_2 _22843_ (.A(_09480_),
    .B(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__inv_2 _22844_ (.A(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__and2b_2 _22845_ (.A_N(\systolic_inst.A_outs[1][1] ),
    .B(\systolic_inst.B_outs[1][7] ),
    .X(_09526_));
 sky130_fd_sc_hd__nand2_2 _22846_ (.A(\systolic_inst.A_outs[1][2] ),
    .B(\systolic_inst.B_outs[1][6] ),
    .Y(_09527_));
 sky130_fd_sc_hd__and3_2 _22847_ (.A(\systolic_inst.A_outs[1][2] ),
    .B(\systolic_inst.B_outs[1][6] ),
    .C(_09526_),
    .X(_09528_));
 sky130_fd_sc_hd__xnor2_2 _22848_ (.A(_09526_),
    .B(_09527_),
    .Y(_09529_));
 sky130_fd_sc_hd__xnor2_2 _22849_ (.A(_09489_),
    .B(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__nand2_2 _22850_ (.A(\systolic_inst.A_outs[1][0] ),
    .B(_09461_),
    .Y(_09531_));
 sky130_fd_sc_hd__nand2_2 _22851_ (.A(\systolic_inst.B_outs[1][7] ),
    .B(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__and3_2 _22852_ (.A(\systolic_inst.B_outs[1][7] ),
    .B(_09530_),
    .C(_09531_),
    .X(_09533_));
 sky130_fd_sc_hd__xor2_2 _22853_ (.A(_09530_),
    .B(_09532_),
    .X(_09534_));
 sky130_fd_sc_hd__xnor2_2 _22854_ (.A(_09525_),
    .B(_09534_),
    .Y(_09535_));
 sky130_fd_sc_hd__o31a_2 _22855_ (.A1(\systolic_inst.B_outs[1][7] ),
    .A2(_09429_),
    .A3(_09461_),
    .B1(_09497_),
    .X(_09536_));
 sky130_fd_sc_hd__or2_2 _22856_ (.A(_09535_),
    .B(_09536_),
    .X(_09537_));
 sky130_fd_sc_hd__xnor2_2 _22857_ (.A(_09535_),
    .B(_09536_),
    .Y(_09538_));
 sky130_fd_sc_hd__xnor2_2 _22858_ (.A(_09520_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__o21ai_2 _22859_ (.A1(_09464_),
    .A2(_09498_),
    .B1(_09500_),
    .Y(_09540_));
 sky130_fd_sc_hd__nand2b_2 _22860_ (.A_N(_09539_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__xnor2_2 _22861_ (.A(_09539_),
    .B(_09540_),
    .Y(_09542_));
 sky130_fd_sc_hd__nand2b_2 _22862_ (.A_N(_09512_),
    .B(_09542_),
    .Y(_09543_));
 sky130_fd_sc_hd__xnor2_2 _22863_ (.A(_09512_),
    .B(_09542_),
    .Y(_09544_));
 sky130_fd_sc_hd__nor2_2 _22864_ (.A(_09503_),
    .B(_09505_),
    .Y(_09545_));
 sky130_fd_sc_hd__nand2b_2 _22865_ (.A_N(_09545_),
    .B(_09544_),
    .Y(_09546_));
 sky130_fd_sc_hd__xnor2_2 _22866_ (.A(_09544_),
    .B(_09545_),
    .Y(_09547_));
 sky130_fd_sc_hd__a21oi_2 _22867_ (.A1(_09508_),
    .A2(_09510_),
    .B1(_09507_),
    .Y(_09548_));
 sky130_fd_sc_hd__nand2b_2 _22868_ (.A_N(_09548_),
    .B(_09547_),
    .Y(_09549_));
 sky130_fd_sc_hd__nand2b_2 _22869_ (.A_N(_09547_),
    .B(_09548_),
    .Y(_09550_));
 sky130_fd_sc_hd__and2_2 _22870_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[8] ),
    .X(_09551_));
 sky130_fd_sc_hd__a31o_2 _22871_ (.A1(\systolic_inst.ce_local ),
    .A2(_09549_),
    .A3(_09550_),
    .B1(_09551_),
    .X(_01866_));
 sky130_fd_sc_hd__a21o_2 _22872_ (.A1(_09513_),
    .A2(_09519_),
    .B1(_09518_),
    .X(_09552_));
 sky130_fd_sc_hd__o21ba_2 _22873_ (.A1(_09480_),
    .A2(_09522_),
    .B1_N(_09521_),
    .X(_09553_));
 sky130_fd_sc_hd__nor2_2 _22874_ (.A(_09515_),
    .B(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__and2_2 _22875_ (.A(_09515_),
    .B(_09553_),
    .X(_09555_));
 sky130_fd_sc_hd__or2_2 _22876_ (.A(_09554_),
    .B(_09555_),
    .X(_09556_));
 sky130_fd_sc_hd__nand2_2 _22877_ (.A(\systolic_inst.B_outs[1][2] ),
    .B(\systolic_inst.A_outs[1][7] ),
    .Y(_09557_));
 sky130_fd_sc_hd__a22oi_2 _22878_ (.A1(\systolic_inst.B_outs[1][4] ),
    .A2(\systolic_inst.A_outs[1][5] ),
    .B1(\systolic_inst.A_outs[1][6] ),
    .B2(\systolic_inst.B_outs[1][3] ),
    .Y(_09558_));
 sky130_fd_sc_hd__and4_2 _22879_ (.A(\systolic_inst.B_outs[1][3] ),
    .B(\systolic_inst.B_outs[1][4] ),
    .C(\systolic_inst.A_outs[1][5] ),
    .D(\systolic_inst.A_outs[1][6] ),
    .X(_09559_));
 sky130_fd_sc_hd__nor2_2 _22880_ (.A(_09558_),
    .B(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__xnor2_2 _22881_ (.A(_09557_),
    .B(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__nand2_2 _22882_ (.A(\systolic_inst.A_outs[1][4] ),
    .B(\systolic_inst.B_outs[1][5] ),
    .Y(_09562_));
 sky130_fd_sc_hd__and4b_2 _22883_ (.A_N(\systolic_inst.A_outs[1][2] ),
    .B(\systolic_inst.A_outs[1][3] ),
    .C(\systolic_inst.B_outs[1][6] ),
    .D(\systolic_inst.B_outs[1][7] ),
    .X(_09563_));
 sky130_fd_sc_hd__o2bb2a_2 _22884_ (.A1_N(\systolic_inst.A_outs[1][3] ),
    .A2_N(\systolic_inst.B_outs[1][6] ),
    .B1(_11277_),
    .B2(\systolic_inst.A_outs[1][2] ),
    .X(_09564_));
 sky130_fd_sc_hd__nor2_2 _22885_ (.A(_09563_),
    .B(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__xnor2_2 _22886_ (.A(_09562_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__a31oi_2 _22887_ (.A1(\systolic_inst.A_outs[1][3] ),
    .A2(\systolic_inst.B_outs[1][5] ),
    .A3(_09529_),
    .B1(_09528_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand2b_2 _22888_ (.A_N(_09567_),
    .B(_09566_),
    .Y(_09568_));
 sky130_fd_sc_hd__xnor2_2 _22889_ (.A(_09566_),
    .B(_09567_),
    .Y(_09569_));
 sky130_fd_sc_hd__xnor2_2 _22890_ (.A(_09561_),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__o21ba_2 _22891_ (.A1(_09525_),
    .A2(_09534_),
    .B1_N(_09533_),
    .X(_09571_));
 sky130_fd_sc_hd__xnor2_2 _22892_ (.A(_09570_),
    .B(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__or2_2 _22893_ (.A(_09556_),
    .B(_09572_),
    .X(_09573_));
 sky130_fd_sc_hd__nand2_2 _22894_ (.A(_09556_),
    .B(_09572_),
    .Y(_09574_));
 sky130_fd_sc_hd__and2_2 _22895_ (.A(_09573_),
    .B(_09574_),
    .X(_09575_));
 sky130_fd_sc_hd__o21a_2 _22896_ (.A1(_09520_),
    .A2(_09538_),
    .B1(_09537_),
    .X(_09576_));
 sky130_fd_sc_hd__nand2b_2 _22897_ (.A_N(_09576_),
    .B(_09575_),
    .Y(_09577_));
 sky130_fd_sc_hd__xnor2_2 _22898_ (.A(_09575_),
    .B(_09576_),
    .Y(_09578_));
 sky130_fd_sc_hd__xnor2_2 _22899_ (.A(_09552_),
    .B(_09578_),
    .Y(_09579_));
 sky130_fd_sc_hd__a21o_2 _22900_ (.A1(_09541_),
    .A2(_09543_),
    .B1(_09579_),
    .X(_09580_));
 sky130_fd_sc_hd__nand3_2 _22901_ (.A(_09541_),
    .B(_09543_),
    .C(_09579_),
    .Y(_09581_));
 sky130_fd_sc_hd__nand2_2 _22902_ (.A(_09580_),
    .B(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__nand2_2 _22903_ (.A(_09546_),
    .B(_09549_),
    .Y(_09583_));
 sky130_fd_sc_hd__xnor2_2 _22904_ (.A(_09582_),
    .B(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__mux2_1 _22905_ (.A0(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[9] ),
    .A1(_09584_),
    .S(\systolic_inst.ce_local ),
    .X(_01867_));
 sky130_fd_sc_hd__o21ba_2 _22906_ (.A1(_09557_),
    .A2(_09558_),
    .B1_N(_09559_),
    .X(_09585_));
 sky130_fd_sc_hd__nor2_2 _22907_ (.A(_09515_),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__and2_2 _22908_ (.A(_09515_),
    .B(_09585_),
    .X(_09587_));
 sky130_fd_sc_hd__or2_2 _22909_ (.A(_09586_),
    .B(_09587_),
    .X(_09588_));
 sky130_fd_sc_hd__a22o_2 _22910_ (.A1(\systolic_inst.B_outs[1][4] ),
    .A2(\systolic_inst.A_outs[1][6] ),
    .B1(\systolic_inst.A_outs[1][7] ),
    .B2(\systolic_inst.B_outs[1][3] ),
    .X(_09589_));
 sky130_fd_sc_hd__and3_2 _22911_ (.A(\systolic_inst.B_outs[1][3] ),
    .B(\systolic_inst.B_outs[1][4] ),
    .C(\systolic_inst.A_outs[1][7] ),
    .X(_09590_));
 sky130_fd_sc_hd__a21bo_2 _22912_ (.A1(\systolic_inst.A_outs[1][6] ),
    .A2(_09590_),
    .B1_N(_09589_),
    .X(_09591_));
 sky130_fd_sc_hd__xor2_2 _22913_ (.A(_09557_),
    .B(_09591_),
    .X(_09592_));
 sky130_fd_sc_hd__nand2_2 _22914_ (.A(\systolic_inst.B_outs[1][5] ),
    .B(\systolic_inst.A_outs[1][5] ),
    .Y(_09593_));
 sky130_fd_sc_hd__and4b_2 _22915_ (.A_N(\systolic_inst.A_outs[1][3] ),
    .B(\systolic_inst.A_outs[1][4] ),
    .C(\systolic_inst.B_outs[1][6] ),
    .D(\systolic_inst.B_outs[1][7] ),
    .X(_09594_));
 sky130_fd_sc_hd__o2bb2a_2 _22916_ (.A1_N(\systolic_inst.A_outs[1][4] ),
    .A2_N(\systolic_inst.B_outs[1][6] ),
    .B1(_11277_),
    .B2(\systolic_inst.A_outs[1][3] ),
    .X(_09595_));
 sky130_fd_sc_hd__nor2_2 _22917_ (.A(_09594_),
    .B(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__xnor2_2 _22918_ (.A(_09593_),
    .B(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__o21ba_2 _22919_ (.A1(_09562_),
    .A2(_09564_),
    .B1_N(_09563_),
    .X(_09598_));
 sky130_fd_sc_hd__nand2b_2 _22920_ (.A_N(_09598_),
    .B(_09597_),
    .Y(_09599_));
 sky130_fd_sc_hd__xnor2_2 _22921_ (.A(_09597_),
    .B(_09598_),
    .Y(_09600_));
 sky130_fd_sc_hd__nand2_2 _22922_ (.A(_09592_),
    .B(_09600_),
    .Y(_09601_));
 sky130_fd_sc_hd__or2_2 _22923_ (.A(_09592_),
    .B(_09600_),
    .X(_09602_));
 sky130_fd_sc_hd__nand2_2 _22924_ (.A(_09601_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__a21bo_2 _22925_ (.A1(_09561_),
    .A2(_09569_),
    .B1_N(_09568_),
    .X(_09604_));
 sky130_fd_sc_hd__nand2b_2 _22926_ (.A_N(_09603_),
    .B(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__xor2_2 _22927_ (.A(_09603_),
    .B(_09604_),
    .X(_09606_));
 sky130_fd_sc_hd__xor2_2 _22928_ (.A(_09588_),
    .B(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__o21a_2 _22929_ (.A1(_09570_),
    .A2(_09571_),
    .B1(_09573_),
    .X(_09608_));
 sky130_fd_sc_hd__nand2b_2 _22930_ (.A_N(_09608_),
    .B(_09607_),
    .Y(_09609_));
 sky130_fd_sc_hd__xnor2_2 _22931_ (.A(_09607_),
    .B(_09608_),
    .Y(_09610_));
 sky130_fd_sc_hd__nand2_2 _22932_ (.A(_09554_),
    .B(_09610_),
    .Y(_09611_));
 sky130_fd_sc_hd__xnor2_2 _22933_ (.A(_09554_),
    .B(_09610_),
    .Y(_09612_));
 sky130_fd_sc_hd__a21boi_2 _22934_ (.A1(_09552_),
    .A2(_09578_),
    .B1_N(_09577_),
    .Y(_09613_));
 sky130_fd_sc_hd__or2_2 _22935_ (.A(_09612_),
    .B(_09613_),
    .X(_09614_));
 sky130_fd_sc_hd__nand2_2 _22936_ (.A(_09612_),
    .B(_09613_),
    .Y(_09615_));
 sky130_fd_sc_hd__nand2_2 _22937_ (.A(_09614_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__nand2_2 _22938_ (.A(_09581_),
    .B(_09583_),
    .Y(_09617_));
 sky130_fd_sc_hd__and3_2 _22939_ (.A(_09580_),
    .B(_09616_),
    .C(_09617_),
    .X(_09618_));
 sky130_fd_sc_hd__a21o_2 _22940_ (.A1(_09580_),
    .A2(_09617_),
    .B1(_09616_),
    .X(_09619_));
 sky130_fd_sc_hd__nand2_2 _22941_ (.A(\systolic_inst.ce_local ),
    .B(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__a2bb2o_2 _22942_ (.A1_N(_09620_),
    .A2_N(_09618_),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[10] ),
    .B2(_11258_),
    .X(_01868_));
 sky130_fd_sc_hd__o2bb2a_2 _22943_ (.A1_N(\systolic_inst.A_outs[1][6] ),
    .A2_N(_09590_),
    .B1(_09591_),
    .B2(_09557_),
    .X(_09621_));
 sky130_fd_sc_hd__or2_2 _22944_ (.A(_09515_),
    .B(_09621_),
    .X(_09622_));
 sky130_fd_sc_hd__nand2_2 _22945_ (.A(_09515_),
    .B(_09621_),
    .Y(_09623_));
 sky130_fd_sc_hd__nand2_2 _22946_ (.A(_09622_),
    .B(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__or2_2 _22947_ (.A(\systolic_inst.B_outs[1][3] ),
    .B(\systolic_inst.B_outs[1][4] ),
    .X(_09625_));
 sky130_fd_sc_hd__and3b_2 _22948_ (.A_N(_09590_),
    .B(_09625_),
    .C(\systolic_inst.A_outs[1][7] ),
    .X(_09626_));
 sky130_fd_sc_hd__xnor2_2 _22949_ (.A(_09557_),
    .B(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__nand2_2 _22950_ (.A(\systolic_inst.B_outs[1][5] ),
    .B(\systolic_inst.A_outs[1][6] ),
    .Y(_09628_));
 sky130_fd_sc_hd__and4b_2 _22951_ (.A_N(\systolic_inst.A_outs[1][4] ),
    .B(\systolic_inst.A_outs[1][5] ),
    .C(\systolic_inst.B_outs[1][6] ),
    .D(\systolic_inst.B_outs[1][7] ),
    .X(_09629_));
 sky130_fd_sc_hd__o2bb2a_2 _22952_ (.A1_N(\systolic_inst.A_outs[1][5] ),
    .A2_N(\systolic_inst.B_outs[1][6] ),
    .B1(_11277_),
    .B2(\systolic_inst.A_outs[1][4] ),
    .X(_09630_));
 sky130_fd_sc_hd__or2_2 _22953_ (.A(_09629_),
    .B(_09630_),
    .X(_09631_));
 sky130_fd_sc_hd__xor2_2 _22954_ (.A(_09628_),
    .B(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__o21ba_2 _22955_ (.A1(_09593_),
    .A2(_09595_),
    .B1_N(_09594_),
    .X(_09633_));
 sky130_fd_sc_hd__nand2b_2 _22956_ (.A_N(_09633_),
    .B(_09632_),
    .Y(_09634_));
 sky130_fd_sc_hd__xnor2_2 _22957_ (.A(_09632_),
    .B(_09633_),
    .Y(_09635_));
 sky130_fd_sc_hd__nand2_2 _22958_ (.A(_09627_),
    .B(_09635_),
    .Y(_09636_));
 sky130_fd_sc_hd__xnor2_2 _22959_ (.A(_09627_),
    .B(_09635_),
    .Y(_09637_));
 sky130_fd_sc_hd__a21o_2 _22960_ (.A1(_09599_),
    .A2(_09601_),
    .B1(_09637_),
    .X(_09638_));
 sky130_fd_sc_hd__nand3_2 _22961_ (.A(_09599_),
    .B(_09601_),
    .C(_09637_),
    .Y(_09639_));
 sky130_fd_sc_hd__nand2_2 _22962_ (.A(_09638_),
    .B(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__xor2_2 _22963_ (.A(_09624_),
    .B(_09640_),
    .X(_09641_));
 sky130_fd_sc_hd__o21a_2 _22964_ (.A1(_09588_),
    .A2(_09606_),
    .B1(_09605_),
    .X(_09642_));
 sky130_fd_sc_hd__and2b_2 _22965_ (.A_N(_09642_),
    .B(_09641_),
    .X(_09643_));
 sky130_fd_sc_hd__and2b_2 _22966_ (.A_N(_09641_),
    .B(_09642_),
    .X(_09644_));
 sky130_fd_sc_hd__nor2_2 _22967_ (.A(_09643_),
    .B(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__xnor2_2 _22968_ (.A(_09586_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__and3_2 _22969_ (.A(_09609_),
    .B(_09611_),
    .C(_09646_),
    .X(_09647_));
 sky130_fd_sc_hd__a21o_2 _22970_ (.A1(_09609_),
    .A2(_09611_),
    .B1(_09646_),
    .X(_09648_));
 sky130_fd_sc_hd__nand2b_2 _22971_ (.A_N(_09647_),
    .B(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__nand2_2 _22972_ (.A(_09614_),
    .B(_09619_),
    .Y(_09650_));
 sky130_fd_sc_hd__xnor2_2 _22973_ (.A(_09649_),
    .B(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__mux2_1 _22974_ (.A0(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[11] ),
    .A1(_09651_),
    .S(\systolic_inst.ce_local ),
    .X(_01869_));
 sky130_fd_sc_hd__a31o_2 _22975_ (.A1(\systolic_inst.B_outs[1][2] ),
    .A2(\systolic_inst.A_outs[1][7] ),
    .A3(_09625_),
    .B1(_09590_),
    .X(_09652_));
 sky130_fd_sc_hd__or2_2 _22976_ (.A(_09516_),
    .B(_09652_),
    .X(_09653_));
 sky130_fd_sc_hd__nand2_2 _22977_ (.A(_09516_),
    .B(_09652_),
    .Y(_09654_));
 sky130_fd_sc_hd__nand2_2 _22978_ (.A(_09653_),
    .B(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__inv_2 _22979_ (.A(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__o2bb2a_2 _22980_ (.A1_N(\systolic_inst.B_outs[1][6] ),
    .A2_N(\systolic_inst.A_outs[1][6] ),
    .B1(_11277_),
    .B2(\systolic_inst.A_outs[1][5] ),
    .X(_09657_));
 sky130_fd_sc_hd__and4b_2 _22981_ (.A_N(\systolic_inst.A_outs[1][5] ),
    .B(\systolic_inst.B_outs[1][6] ),
    .C(\systolic_inst.A_outs[1][6] ),
    .D(\systolic_inst.B_outs[1][7] ),
    .X(_09658_));
 sky130_fd_sc_hd__nor2_2 _22982_ (.A(_09657_),
    .B(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__nand2_2 _22983_ (.A(\systolic_inst.B_outs[1][5] ),
    .B(\systolic_inst.A_outs[1][7] ),
    .Y(_09660_));
 sky130_fd_sc_hd__and3_2 _22984_ (.A(\systolic_inst.B_outs[1][5] ),
    .B(\systolic_inst.A_outs[1][7] ),
    .C(_09659_),
    .X(_09661_));
 sky130_fd_sc_hd__xnor2_2 _22985_ (.A(_09659_),
    .B(_09660_),
    .Y(_09662_));
 sky130_fd_sc_hd__o21ba_2 _22986_ (.A1(_09628_),
    .A2(_09630_),
    .B1_N(_09629_),
    .X(_09663_));
 sky130_fd_sc_hd__nand2b_2 _22987_ (.A_N(_09663_),
    .B(_09662_),
    .Y(_09664_));
 sky130_fd_sc_hd__xnor2_2 _22988_ (.A(_09662_),
    .B(_09663_),
    .Y(_09665_));
 sky130_fd_sc_hd__xnor2_2 _22989_ (.A(_09627_),
    .B(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__a21o_2 _22990_ (.A1(_09634_),
    .A2(_09636_),
    .B1(_09666_),
    .X(_09667_));
 sky130_fd_sc_hd__nand3_2 _22991_ (.A(_09634_),
    .B(_09636_),
    .C(_09666_),
    .Y(_09668_));
 sky130_fd_sc_hd__nand2_2 _22992_ (.A(_09667_),
    .B(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__xnor2_2 _22993_ (.A(_09656_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__o21a_2 _22994_ (.A1(_09624_),
    .A2(_09640_),
    .B1(_09638_),
    .X(_09671_));
 sky130_fd_sc_hd__and2b_2 _22995_ (.A_N(_09671_),
    .B(_09670_),
    .X(_09672_));
 sky130_fd_sc_hd__and2b_2 _22996_ (.A_N(_09670_),
    .B(_09671_),
    .X(_09673_));
 sky130_fd_sc_hd__nor2_2 _22997_ (.A(_09672_),
    .B(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__and2b_2 _22998_ (.A_N(_09622_),
    .B(_09674_),
    .X(_09675_));
 sky130_fd_sc_hd__xor2_2 _22999_ (.A(_09622_),
    .B(_09674_),
    .X(_09676_));
 sky130_fd_sc_hd__a21oi_2 _23000_ (.A1(_09586_),
    .A2(_09645_),
    .B1(_09643_),
    .Y(_09677_));
 sky130_fd_sc_hd__or2_2 _23001_ (.A(_09676_),
    .B(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__inv_2 _23002_ (.A(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__nand2_2 _23003_ (.A(_09676_),
    .B(_09677_),
    .Y(_09680_));
 sky130_fd_sc_hd__nand2_2 _23004_ (.A(_09678_),
    .B(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__a31o_2 _23005_ (.A1(_09614_),
    .A2(_09619_),
    .A3(_09648_),
    .B1(_09647_),
    .X(_09682_));
 sky130_fd_sc_hd__nand2_2 _23006_ (.A(_09681_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__a311oi_2 _23007_ (.A1(_09614_),
    .A2(_09619_),
    .A3(_09648_),
    .B1(_09681_),
    .C1(_09647_),
    .Y(_09684_));
 sky130_fd_sc_hd__nor2_2 _23008_ (.A(_11258_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__a22o_2 _23009_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[12] ),
    .B1(_09683_),
    .B2(_09685_),
    .X(_01870_));
 sky130_fd_sc_hd__nand2_2 _23010_ (.A(\systolic_inst.B_outs[1][6] ),
    .B(\systolic_inst.A_outs[1][7] ),
    .Y(_09686_));
 sky130_fd_sc_hd__nor2_2 _23011_ (.A(\systolic_inst.A_outs[1][6] ),
    .B(_11277_),
    .Y(_09687_));
 sky130_fd_sc_hd__xnor2_2 _23012_ (.A(_09686_),
    .B(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__nand2b_2 _23013_ (.A_N(_09660_),
    .B(_09688_),
    .Y(_09689_));
 sky130_fd_sc_hd__xnor2_2 _23014_ (.A(_09660_),
    .B(_09688_),
    .Y(_09690_));
 sky130_fd_sc_hd__o21ai_2 _23015_ (.A1(_09658_),
    .A2(_09661_),
    .B1(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__or3_2 _23016_ (.A(_09658_),
    .B(_09661_),
    .C(_09690_),
    .X(_09692_));
 sky130_fd_sc_hd__and2_2 _23017_ (.A(_09691_),
    .B(_09692_),
    .X(_09693_));
 sky130_fd_sc_hd__nand2_2 _23018_ (.A(_09627_),
    .B(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__or2_2 _23019_ (.A(_09627_),
    .B(_09693_),
    .X(_09695_));
 sky130_fd_sc_hd__nand2_2 _23020_ (.A(_09694_),
    .B(_09695_),
    .Y(_09696_));
 sky130_fd_sc_hd__a21bo_2 _23021_ (.A1(_09627_),
    .A2(_09665_),
    .B1_N(_09664_),
    .X(_09697_));
 sky130_fd_sc_hd__nand2b_2 _23022_ (.A_N(_09696_),
    .B(_09697_),
    .Y(_09698_));
 sky130_fd_sc_hd__xor2_2 _23023_ (.A(_09696_),
    .B(_09697_),
    .X(_09699_));
 sky130_fd_sc_hd__xnor2_2 _23024_ (.A(_09656_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__o21a_2 _23025_ (.A1(_09655_),
    .A2(_09669_),
    .B1(_09667_),
    .X(_09701_));
 sky130_fd_sc_hd__and2b_2 _23026_ (.A_N(_09701_),
    .B(_09700_),
    .X(_09702_));
 sky130_fd_sc_hd__and2b_2 _23027_ (.A_N(_09700_),
    .B(_09701_),
    .X(_09703_));
 sky130_fd_sc_hd__nor2_2 _23028_ (.A(_09702_),
    .B(_09703_),
    .Y(_09704_));
 sky130_fd_sc_hd__xnor2_2 _23029_ (.A(_09654_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__o21a_2 _23030_ (.A1(_09672_),
    .A2(_09675_),
    .B1(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__nor3_2 _23031_ (.A(_09672_),
    .B(_09675_),
    .C(_09705_),
    .Y(_09707_));
 sky130_fd_sc_hd__inv_2 _23032_ (.A(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__nor2_2 _23033_ (.A(_09706_),
    .B(_09707_),
    .Y(_09709_));
 sky130_fd_sc_hd__or3_2 _23034_ (.A(_09679_),
    .B(_09684_),
    .C(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__o21ai_2 _23035_ (.A1(_09679_),
    .A2(_09684_),
    .B1(_09709_),
    .Y(_09711_));
 sky130_fd_sc_hd__and2_2 _23036_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[13] ),
    .X(_09712_));
 sky130_fd_sc_hd__a31o_2 _23037_ (.A1(\systolic_inst.ce_local ),
    .A2(_09710_),
    .A3(_09711_),
    .B1(_09712_),
    .X(_01871_));
 sky130_fd_sc_hd__and2_2 _23038_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[14] ),
    .X(_09713_));
 sky130_fd_sc_hd__o211ai_2 _23039_ (.A1(_11277_),
    .A2(\systolic_inst.A_outs[1][7] ),
    .B1(_09660_),
    .C1(_09686_),
    .Y(_09714_));
 sky130_fd_sc_hd__o311a_2 _23040_ (.A1(\systolic_inst.A_outs[1][6] ),
    .A2(_11277_),
    .A3(_09686_),
    .B1(_09689_),
    .C1(_09714_),
    .X(_09715_));
 sky130_fd_sc_hd__a31o_2 _23041_ (.A1(\systolic_inst.B_outs[1][5] ),
    .A2(\systolic_inst.B_outs[1][6] ),
    .A3(\systolic_inst.A_outs[1][7] ),
    .B1(_09715_),
    .X(_09716_));
 sky130_fd_sc_hd__nor2_2 _23042_ (.A(_09627_),
    .B(_09716_),
    .Y(_09717_));
 sky130_fd_sc_hd__and2_2 _23043_ (.A(_09627_),
    .B(_09716_),
    .X(_09718_));
 sky130_fd_sc_hd__or2_2 _23044_ (.A(_09717_),
    .B(_09718_),
    .X(_09719_));
 sky130_fd_sc_hd__a21oi_2 _23045_ (.A1(_09691_),
    .A2(_09694_),
    .B1(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__and3_2 _23046_ (.A(_09691_),
    .B(_09694_),
    .C(_09719_),
    .X(_09721_));
 sky130_fd_sc_hd__nor2_2 _23047_ (.A(_09720_),
    .B(_09721_),
    .Y(_09722_));
 sky130_fd_sc_hd__xnor2_2 _23048_ (.A(_09655_),
    .B(_09722_),
    .Y(_09723_));
 sky130_fd_sc_hd__o21a_2 _23049_ (.A1(_09655_),
    .A2(_09699_),
    .B1(_09698_),
    .X(_09724_));
 sky130_fd_sc_hd__and2b_2 _23050_ (.A_N(_09724_),
    .B(_09723_),
    .X(_09725_));
 sky130_fd_sc_hd__and2b_2 _23051_ (.A_N(_09723_),
    .B(_09724_),
    .X(_09726_));
 sky130_fd_sc_hd__nor2_2 _23052_ (.A(_09725_),
    .B(_09726_),
    .Y(_09727_));
 sky130_fd_sc_hd__xnor2_2 _23053_ (.A(_09654_),
    .B(_09727_),
    .Y(_09728_));
 sky130_fd_sc_hd__o21ba_2 _23054_ (.A1(_09654_),
    .A2(_09703_),
    .B1_N(_09702_),
    .X(_09729_));
 sky130_fd_sc_hd__nand2b_2 _23055_ (.A_N(_09729_),
    .B(_09728_),
    .Y(_09730_));
 sky130_fd_sc_hd__xnor2_2 _23056_ (.A(_09728_),
    .B(_09729_),
    .Y(_09731_));
 sky130_fd_sc_hd__o31a_2 _23057_ (.A1(_09679_),
    .A2(_09684_),
    .A3(_09706_),
    .B1(_09708_),
    .X(_09732_));
 sky130_fd_sc_hd__or2_2 _23058_ (.A(_09731_),
    .B(_09732_),
    .X(_09733_));
 sky130_fd_sc_hd__nand2_2 _23059_ (.A(_09731_),
    .B(_09732_),
    .Y(_09734_));
 sky130_fd_sc_hd__a31o_2 _23060_ (.A1(\systolic_inst.ce_local ),
    .A2(_09733_),
    .A3(_09734_),
    .B1(_09713_),
    .X(_01872_));
 sky130_fd_sc_hd__a31oi_2 _23061_ (.A1(_09516_),
    .A2(_09652_),
    .A3(_09727_),
    .B1(_09725_),
    .Y(_09735_));
 sky130_fd_sc_hd__a21oi_2 _23062_ (.A1(_09656_),
    .A2(_09722_),
    .B1(_09720_),
    .Y(_09736_));
 sky130_fd_sc_hd__xnor2_2 _23063_ (.A(_09653_),
    .B(_09717_),
    .Y(_09737_));
 sky130_fd_sc_hd__xnor2_2 _23064_ (.A(_09736_),
    .B(_09737_),
    .Y(_09738_));
 sky130_fd_sc_hd__xnor2_2 _23065_ (.A(_09735_),
    .B(_09738_),
    .Y(_09739_));
 sky130_fd_sc_hd__and3_2 _23066_ (.A(\systolic_inst.ce_local ),
    .B(_09730_),
    .C(_09739_),
    .X(_09740_));
 sky130_fd_sc_hd__a22o_2 _23067_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B1(_09734_),
    .B2(_09740_),
    .X(_01873_));
 sky130_fd_sc_hd__a21o_2 _23068_ (.A1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[1][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_09741_));
 sky130_fd_sc_hd__a21oi_2 _23069_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[1][0] ),
    .Y(_09742_));
 sky130_fd_sc_hd__a21oi_2 _23070_ (.A1(\systolic_inst.ce_local ),
    .A2(_09741_),
    .B1(_09742_),
    .Y(_01874_));
 sky130_fd_sc_hd__and2_2 _23071_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[1][1] ),
    .X(_09743_));
 sky130_fd_sc_hd__nand2_2 _23072_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[1][1] ),
    .Y(_09744_));
 sky130_fd_sc_hd__or2_2 _23073_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[1][1] ),
    .X(_09745_));
 sky130_fd_sc_hd__and4_2 _23074_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[1][0] ),
    .C(_09744_),
    .D(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__inv_2 _23075_ (.A(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__a22o_2 _23076_ (.A1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[1][0] ),
    .B1(_09744_),
    .B2(_09745_),
    .X(_09748_));
 sky130_fd_sc_hd__a32o_2 _23077_ (.A1(_11712_),
    .A2(_09747_),
    .A3(_09748_),
    .B1(\systolic_inst.acc_wires[1][1] ),
    .B2(_11258_),
    .X(_01875_));
 sky130_fd_sc_hd__nand2_2 _23078_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[1][2] ),
    .Y(_09749_));
 sky130_fd_sc_hd__or2_2 _23079_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[1][2] ),
    .X(_09750_));
 sky130_fd_sc_hd__a31o_2 _23080_ (.A1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[1][0] ),
    .A3(_09745_),
    .B1(_09743_),
    .X(_09751_));
 sky130_fd_sc_hd__a21o_2 _23081_ (.A1(_09749_),
    .A2(_09750_),
    .B1(_09751_),
    .X(_09752_));
 sky130_fd_sc_hd__and3_2 _23082_ (.A(_09749_),
    .B(_09750_),
    .C(_09751_),
    .X(_09753_));
 sky130_fd_sc_hd__inv_2 _23083_ (.A(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__a32o_2 _23084_ (.A1(_11712_),
    .A2(_09752_),
    .A3(_09754_),
    .B1(\systolic_inst.acc_wires[1][2] ),
    .B2(_11258_),
    .X(_01876_));
 sky130_fd_sc_hd__nand2_2 _23085_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[1][3] ),
    .Y(_09755_));
 sky130_fd_sc_hd__or2_2 _23086_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[1][3] ),
    .X(_09756_));
 sky130_fd_sc_hd__a21bo_2 _23087_ (.A1(_09750_),
    .A2(_09751_),
    .B1_N(_09749_),
    .X(_09757_));
 sky130_fd_sc_hd__a21o_2 _23088_ (.A1(_09755_),
    .A2(_09756_),
    .B1(_09757_),
    .X(_09758_));
 sky130_fd_sc_hd__and3_2 _23089_ (.A(_09755_),
    .B(_09756_),
    .C(_09757_),
    .X(_09759_));
 sky130_fd_sc_hd__inv_2 _23090_ (.A(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__a32o_2 _23091_ (.A1(_11712_),
    .A2(_09758_),
    .A3(_09760_),
    .B1(\systolic_inst.acc_wires[1][3] ),
    .B2(_11258_),
    .X(_01877_));
 sky130_fd_sc_hd__nand2_2 _23092_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[1][4] ),
    .Y(_09761_));
 sky130_fd_sc_hd__or2_2 _23093_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[1][4] ),
    .X(_09762_));
 sky130_fd_sc_hd__a21bo_2 _23094_ (.A1(_09756_),
    .A2(_09757_),
    .B1_N(_09755_),
    .X(_09763_));
 sky130_fd_sc_hd__a21o_2 _23095_ (.A1(_09761_),
    .A2(_09762_),
    .B1(_09763_),
    .X(_09764_));
 sky130_fd_sc_hd__and3_2 _23096_ (.A(_09761_),
    .B(_09762_),
    .C(_09763_),
    .X(_09765_));
 sky130_fd_sc_hd__inv_2 _23097_ (.A(_09765_),
    .Y(_09766_));
 sky130_fd_sc_hd__a32o_2 _23098_ (.A1(_11712_),
    .A2(_09764_),
    .A3(_09766_),
    .B1(\systolic_inst.acc_wires[1][4] ),
    .B2(_11258_),
    .X(_01878_));
 sky130_fd_sc_hd__nand2_2 _23099_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[1][5] ),
    .Y(_09767_));
 sky130_fd_sc_hd__or2_2 _23100_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[1][5] ),
    .X(_09768_));
 sky130_fd_sc_hd__a21bo_2 _23101_ (.A1(_09762_),
    .A2(_09763_),
    .B1_N(_09761_),
    .X(_09769_));
 sky130_fd_sc_hd__a21o_2 _23102_ (.A1(_09767_),
    .A2(_09768_),
    .B1(_09769_),
    .X(_09770_));
 sky130_fd_sc_hd__and3_2 _23103_ (.A(_09767_),
    .B(_09768_),
    .C(_09769_),
    .X(_09771_));
 sky130_fd_sc_hd__inv_2 _23104_ (.A(_09771_),
    .Y(_09772_));
 sky130_fd_sc_hd__a32o_2 _23105_ (.A1(_11712_),
    .A2(_09770_),
    .A3(_09772_),
    .B1(\systolic_inst.acc_wires[1][5] ),
    .B2(_11258_),
    .X(_01879_));
 sky130_fd_sc_hd__nand2_2 _23106_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[1][6] ),
    .Y(_09773_));
 sky130_fd_sc_hd__or2_2 _23107_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[1][6] ),
    .X(_09774_));
 sky130_fd_sc_hd__a21bo_2 _23108_ (.A1(_09768_),
    .A2(_09769_),
    .B1_N(_09767_),
    .X(_09775_));
 sky130_fd_sc_hd__a21o_2 _23109_ (.A1(_09773_),
    .A2(_09774_),
    .B1(_09775_),
    .X(_09776_));
 sky130_fd_sc_hd__and3_2 _23110_ (.A(_09773_),
    .B(_09774_),
    .C(_09775_),
    .X(_09777_));
 sky130_fd_sc_hd__inv_2 _23111_ (.A(_09777_),
    .Y(_09778_));
 sky130_fd_sc_hd__a32o_2 _23112_ (.A1(_11712_),
    .A2(_09776_),
    .A3(_09778_),
    .B1(\systolic_inst.acc_wires[1][6] ),
    .B2(_11258_),
    .X(_01880_));
 sky130_fd_sc_hd__nand2_2 _23113_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[1][7] ),
    .Y(_09779_));
 sky130_fd_sc_hd__or2_2 _23114_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[1][7] ),
    .X(_09780_));
 sky130_fd_sc_hd__a21bo_2 _23115_ (.A1(_09774_),
    .A2(_09775_),
    .B1_N(_09773_),
    .X(_09781_));
 sky130_fd_sc_hd__a21o_2 _23116_ (.A1(_09779_),
    .A2(_09780_),
    .B1(_09781_),
    .X(_09782_));
 sky130_fd_sc_hd__nand3_2 _23117_ (.A(_09779_),
    .B(_09780_),
    .C(_09781_),
    .Y(_09783_));
 sky130_fd_sc_hd__a32o_2 _23118_ (.A1(_11712_),
    .A2(_09782_),
    .A3(_09783_),
    .B1(\systolic_inst.acc_wires[1][7] ),
    .B2(_11258_),
    .X(_01881_));
 sky130_fd_sc_hd__a21bo_2 _23119_ (.A1(_09780_),
    .A2(_09781_),
    .B1_N(_09779_),
    .X(_09784_));
 sky130_fd_sc_hd__xor2_2 _23120_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[1][8] ),
    .X(_09785_));
 sky130_fd_sc_hd__and2_2 _23121_ (.A(_09784_),
    .B(_09785_),
    .X(_09786_));
 sky130_fd_sc_hd__o21ai_2 _23122_ (.A1(_09784_),
    .A2(_09785_),
    .B1(_11712_),
    .Y(_09787_));
 sky130_fd_sc_hd__a2bb2o_2 _23123_ (.A1_N(_09787_),
    .A2_N(_09786_),
    .B1(\systolic_inst.acc_wires[1][8] ),
    .B2(_11258_),
    .X(_01882_));
 sky130_fd_sc_hd__xor2_2 _23124_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[1][9] ),
    .X(_09788_));
 sky130_fd_sc_hd__a211o_2 _23125_ (.A1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[1][8] ),
    .B1(_09786_),
    .C1(_09788_),
    .X(_09789_));
 sky130_fd_sc_hd__nand2_2 _23126_ (.A(_09785_),
    .B(_09788_),
    .Y(_09790_));
 sky130_fd_sc_hd__nand2_2 _23127_ (.A(_09786_),
    .B(_09788_),
    .Y(_09791_));
 sky130_fd_sc_hd__and3_2 _23128_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[1][8] ),
    .C(_09788_),
    .X(_09792_));
 sky130_fd_sc_hd__nor2_2 _23129_ (.A(_11713_),
    .B(_09792_),
    .Y(_09793_));
 sky130_fd_sc_hd__a32o_2 _23130_ (.A1(_09789_),
    .A2(_09791_),
    .A3(_09793_),
    .B1(\systolic_inst.acc_wires[1][9] ),
    .B2(_11258_),
    .X(_01883_));
 sky130_fd_sc_hd__nand2_2 _23131_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[1][10] ),
    .Y(_09794_));
 sky130_fd_sc_hd__or2_2 _23132_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[1][10] ),
    .X(_09795_));
 sky130_fd_sc_hd__and2_2 _23133_ (.A(_09794_),
    .B(_09795_),
    .X(_09796_));
 sky130_fd_sc_hd__a21oi_2 _23134_ (.A1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[1][9] ),
    .B1(_09792_),
    .Y(_09797_));
 sky130_fd_sc_hd__nand2_2 _23135_ (.A(_09791_),
    .B(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__xor2_2 _23136_ (.A(_09796_),
    .B(_09798_),
    .X(_09799_));
 sky130_fd_sc_hd__a22o_2 _23137_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][10] ),
    .B1(_11712_),
    .B2(_09799_),
    .X(_01884_));
 sky130_fd_sc_hd__nor2_2 _23138_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[1][11] ),
    .Y(_09800_));
 sky130_fd_sc_hd__or2_2 _23139_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[1][11] ),
    .X(_09801_));
 sky130_fd_sc_hd__nand2_2 _23140_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[1][11] ),
    .Y(_09802_));
 sky130_fd_sc_hd__nand2_2 _23141_ (.A(_09801_),
    .B(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__a21bo_2 _23142_ (.A1(_09796_),
    .A2(_09798_),
    .B1_N(_09794_),
    .X(_09804_));
 sky130_fd_sc_hd__xnor2_2 _23143_ (.A(_09803_),
    .B(_09804_),
    .Y(_09805_));
 sky130_fd_sc_hd__a22o_2 _23144_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][11] ),
    .B1(_11712_),
    .B2(_09805_),
    .X(_01885_));
 sky130_fd_sc_hd__nand3_2 _23145_ (.A(_09796_),
    .B(_09801_),
    .C(_09802_),
    .Y(_09806_));
 sky130_fd_sc_hd__nor2_2 _23146_ (.A(_09790_),
    .B(_09806_),
    .Y(_09807_));
 sky130_fd_sc_hd__o2bb2a_2 _23147_ (.A1_N(_09784_),
    .A2_N(_09807_),
    .B1(_09797_),
    .B2(_09806_),
    .X(_09808_));
 sky130_fd_sc_hd__o21a_2 _23148_ (.A1(_09794_),
    .A2(_09800_),
    .B1(_09802_),
    .X(_09809_));
 sky130_fd_sc_hd__xnor2_2 _23149_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[1][12] ),
    .Y(_09810_));
 sky130_fd_sc_hd__and3_2 _23150_ (.A(_09808_),
    .B(_09809_),
    .C(_09810_),
    .X(_09811_));
 sky130_fd_sc_hd__a21oi_2 _23151_ (.A1(_09808_),
    .A2(_09809_),
    .B1(_09810_),
    .Y(_09812_));
 sky130_fd_sc_hd__nor2_2 _23152_ (.A(_09811_),
    .B(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__a22o_2 _23153_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][12] ),
    .B1(_11712_),
    .B2(_09813_),
    .X(_01886_));
 sky130_fd_sc_hd__xor2_2 _23154_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[1][13] ),
    .X(_09814_));
 sky130_fd_sc_hd__a211o_2 _23155_ (.A1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[1][12] ),
    .B1(_09812_),
    .C1(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__nand2b_2 _23156_ (.A_N(_09810_),
    .B(_09814_),
    .Y(_09816_));
 sky130_fd_sc_hd__a21o_2 _23157_ (.A1(_09808_),
    .A2(_09809_),
    .B1(_09816_),
    .X(_09817_));
 sky130_fd_sc_hd__and3_2 _23158_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[1][12] ),
    .C(_09814_),
    .X(_09818_));
 sky130_fd_sc_hd__nor2_2 _23159_ (.A(_11713_),
    .B(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__a32o_2 _23160_ (.A1(_09815_),
    .A2(_09817_),
    .A3(_09819_),
    .B1(\systolic_inst.acc_wires[1][13] ),
    .B2(_11258_),
    .X(_01887_));
 sky130_fd_sc_hd__or2_2 _23161_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[1][14] ),
    .X(_09820_));
 sky130_fd_sc_hd__nand2_2 _23162_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[1][14] ),
    .Y(_09821_));
 sky130_fd_sc_hd__and2_2 _23163_ (.A(_09820_),
    .B(_09821_),
    .X(_09822_));
 sky130_fd_sc_hd__nand2_2 _23164_ (.A(_09820_),
    .B(_09821_),
    .Y(_09823_));
 sky130_fd_sc_hd__a21oi_2 _23165_ (.A1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[1][13] ),
    .B1(_09818_),
    .Y(_09824_));
 sky130_fd_sc_hd__nand2_2 _23166_ (.A(_09817_),
    .B(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__nand2_2 _23167_ (.A(_09822_),
    .B(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__or2_2 _23168_ (.A(_09822_),
    .B(_09825_),
    .X(_09827_));
 sky130_fd_sc_hd__a32o_2 _23169_ (.A1(_11712_),
    .A2(_09826_),
    .A3(_09827_),
    .B1(\systolic_inst.acc_wires[1][14] ),
    .B2(_11258_),
    .X(_01888_));
 sky130_fd_sc_hd__nor2_2 _23170_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][15] ),
    .Y(_09828_));
 sky130_fd_sc_hd__and2_2 _23171_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][15] ),
    .X(_09829_));
 sky130_fd_sc_hd__or2_2 _23172_ (.A(_09828_),
    .B(_09829_),
    .X(_09830_));
 sky130_fd_sc_hd__a21oi_2 _23173_ (.A1(_09821_),
    .A2(_09826_),
    .B1(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__a31o_2 _23174_ (.A1(_09821_),
    .A2(_09826_),
    .A3(_09830_),
    .B1(_11713_),
    .X(_09832_));
 sky130_fd_sc_hd__a2bb2o_2 _23175_ (.A1_N(_09832_),
    .A2_N(_09831_),
    .B1(\systolic_inst.acc_wires[1][15] ),
    .B2(_11258_),
    .X(_01889_));
 sky130_fd_sc_hd__a211o_2 _23176_ (.A1(_09817_),
    .A2(_09824_),
    .B1(_09830_),
    .C1(_09823_),
    .X(_09833_));
 sky130_fd_sc_hd__o21ba_2 _23177_ (.A1(_09821_),
    .A2(_09828_),
    .B1_N(_09829_),
    .X(_09834_));
 sky130_fd_sc_hd__and2_2 _23178_ (.A(_09833_),
    .B(_09834_),
    .X(_09835_));
 sky130_fd_sc_hd__xnor2_2 _23179_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][16] ),
    .Y(_09836_));
 sky130_fd_sc_hd__nand2_2 _23180_ (.A(_09835_),
    .B(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__nor2_2 _23181_ (.A(_09835_),
    .B(_09836_),
    .Y(_09838_));
 sky130_fd_sc_hd__nor2_2 _23182_ (.A(_11713_),
    .B(_09838_),
    .Y(_09839_));
 sky130_fd_sc_hd__a22o_2 _23183_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][16] ),
    .B1(_09837_),
    .B2(_09839_),
    .X(_01890_));
 sky130_fd_sc_hd__xor2_2 _23184_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][17] ),
    .X(_09840_));
 sky130_fd_sc_hd__inv_2 _23185_ (.A(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__a21oi_2 _23186_ (.A1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[1][16] ),
    .B1(_09838_),
    .Y(_09842_));
 sky130_fd_sc_hd__xnor2_2 _23187_ (.A(_09840_),
    .B(_09842_),
    .Y(_09843_));
 sky130_fd_sc_hd__a22o_2 _23188_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][17] ),
    .B1(_11712_),
    .B2(_09843_),
    .X(_01891_));
 sky130_fd_sc_hd__or2_2 _23189_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][18] ),
    .X(_09844_));
 sky130_fd_sc_hd__nand2_2 _23190_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][18] ),
    .Y(_09845_));
 sky130_fd_sc_hd__nand2_2 _23191_ (.A(_09844_),
    .B(_09845_),
    .Y(_09846_));
 sky130_fd_sc_hd__o21a_2 _23192_ (.A1(\systolic_inst.acc_wires[1][16] ),
    .A2(\systolic_inst.acc_wires[1][17] ),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .X(_09847_));
 sky130_fd_sc_hd__a21oi_2 _23193_ (.A1(_09838_),
    .A2(_09840_),
    .B1(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__xor2_2 _23194_ (.A(_09846_),
    .B(_09848_),
    .X(_09849_));
 sky130_fd_sc_hd__a22o_2 _23195_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][18] ),
    .B1(_11712_),
    .B2(_09849_),
    .X(_01892_));
 sky130_fd_sc_hd__xnor2_2 _23196_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][19] ),
    .Y(_09850_));
 sky130_fd_sc_hd__o21ai_2 _23197_ (.A1(_09846_),
    .A2(_09848_),
    .B1(_09845_),
    .Y(_09851_));
 sky130_fd_sc_hd__xnor2_2 _23198_ (.A(_09850_),
    .B(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__a22o_2 _23199_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][19] ),
    .B1(_11712_),
    .B2(_09852_),
    .X(_01893_));
 sky130_fd_sc_hd__or2_2 _23200_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][20] ),
    .X(_09853_));
 sky130_fd_sc_hd__nand2_2 _23201_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][20] ),
    .Y(_09854_));
 sky130_fd_sc_hd__and2_2 _23202_ (.A(_09853_),
    .B(_09854_),
    .X(_09855_));
 sky130_fd_sc_hd__or4_2 _23203_ (.A(_09836_),
    .B(_09841_),
    .C(_09846_),
    .D(_09850_),
    .X(_09856_));
 sky130_fd_sc_hd__nor2_2 _23204_ (.A(_09835_),
    .B(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__o41a_2 _23205_ (.A1(\systolic_inst.acc_wires[1][16] ),
    .A2(\systolic_inst.acc_wires[1][17] ),
    .A3(\systolic_inst.acc_wires[1][18] ),
    .A4(\systolic_inst.acc_wires[1][19] ),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .X(_09858_));
 sky130_fd_sc_hd__or3_2 _23206_ (.A(_09855_),
    .B(_09857_),
    .C(_09858_),
    .X(_09859_));
 sky130_fd_sc_hd__o21ai_2 _23207_ (.A1(_09857_),
    .A2(_09858_),
    .B1(_09855_),
    .Y(_09860_));
 sky130_fd_sc_hd__a32o_2 _23208_ (.A1(_11712_),
    .A2(_09859_),
    .A3(_09860_),
    .B1(\systolic_inst.acc_wires[1][20] ),
    .B2(_11258_),
    .X(_01894_));
 sky130_fd_sc_hd__xnor2_2 _23209_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][21] ),
    .Y(_09861_));
 sky130_fd_sc_hd__inv_2 _23210_ (.A(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__a21oi_2 _23211_ (.A1(_09854_),
    .A2(_09860_),
    .B1(_09861_),
    .Y(_09863_));
 sky130_fd_sc_hd__a31o_2 _23212_ (.A1(_09854_),
    .A2(_09860_),
    .A3(_09861_),
    .B1(_11713_),
    .X(_09864_));
 sky130_fd_sc_hd__a2bb2o_2 _23213_ (.A1_N(_09864_),
    .A2_N(_09863_),
    .B1(\systolic_inst.acc_wires[1][21] ),
    .B2(_11258_),
    .X(_01895_));
 sky130_fd_sc_hd__or2_2 _23214_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][22] ),
    .X(_09865_));
 sky130_fd_sc_hd__nand2_2 _23215_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][22] ),
    .Y(_09866_));
 sky130_fd_sc_hd__and2_2 _23216_ (.A(_09865_),
    .B(_09866_),
    .X(_09867_));
 sky130_fd_sc_hd__o21a_2 _23217_ (.A1(\systolic_inst.acc_wires[1][20] ),
    .A2(\systolic_inst.acc_wires[1][21] ),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .X(_09868_));
 sky130_fd_sc_hd__nor2_2 _23218_ (.A(_09860_),
    .B(_09861_),
    .Y(_09869_));
 sky130_fd_sc_hd__o21ai_2 _23219_ (.A1(_09868_),
    .A2(_09869_),
    .B1(_09867_),
    .Y(_09870_));
 sky130_fd_sc_hd__or3_2 _23220_ (.A(_09867_),
    .B(_09868_),
    .C(_09869_),
    .X(_09871_));
 sky130_fd_sc_hd__a32o_2 _23221_ (.A1(_11712_),
    .A2(_09870_),
    .A3(_09871_),
    .B1(\systolic_inst.acc_wires[1][22] ),
    .B2(_11258_),
    .X(_01896_));
 sky130_fd_sc_hd__xor2_2 _23222_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][23] ),
    .X(_09872_));
 sky130_fd_sc_hd__inv_2 _23223_ (.A(_09872_),
    .Y(_09873_));
 sky130_fd_sc_hd__nand3_2 _23224_ (.A(_09866_),
    .B(_09870_),
    .C(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__a21o_2 _23225_ (.A1(_09866_),
    .A2(_09870_),
    .B1(_09873_),
    .X(_09875_));
 sky130_fd_sc_hd__a32o_2 _23226_ (.A1(_11712_),
    .A2(_09874_),
    .A3(_09875_),
    .B1(\systolic_inst.acc_wires[1][23] ),
    .B2(_11258_),
    .X(_01897_));
 sky130_fd_sc_hd__nand4_2 _23227_ (.A(_09855_),
    .B(_09862_),
    .C(_09867_),
    .D(_09872_),
    .Y(_09876_));
 sky130_fd_sc_hd__a211o_2 _23228_ (.A1(_09833_),
    .A2(_09834_),
    .B1(_09856_),
    .C1(_09876_),
    .X(_09877_));
 sky130_fd_sc_hd__o41a_2 _23229_ (.A1(\systolic_inst.acc_wires[1][20] ),
    .A2(\systolic_inst.acc_wires[1][21] ),
    .A3(\systolic_inst.acc_wires[1][22] ),
    .A4(\systolic_inst.acc_wires[1][23] ),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .X(_09878_));
 sky130_fd_sc_hd__nor2_2 _23230_ (.A(_09858_),
    .B(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__nor2_2 _23231_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][24] ),
    .Y(_09880_));
 sky130_fd_sc_hd__and2_2 _23232_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][24] ),
    .X(_09881_));
 sky130_fd_sc_hd__or2_2 _23233_ (.A(_09880_),
    .B(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__a21oi_2 _23234_ (.A1(_09877_),
    .A2(_09879_),
    .B1(_09882_),
    .Y(_09883_));
 sky130_fd_sc_hd__a31o_2 _23235_ (.A1(_09877_),
    .A2(_09879_),
    .A3(_09882_),
    .B1(_11713_),
    .X(_09884_));
 sky130_fd_sc_hd__a2bb2o_2 _23236_ (.A1_N(_09884_),
    .A2_N(_09883_),
    .B1(\systolic_inst.acc_wires[1][24] ),
    .B2(_11258_),
    .X(_01898_));
 sky130_fd_sc_hd__xor2_2 _23237_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][25] ),
    .X(_09885_));
 sky130_fd_sc_hd__or3_2 _23238_ (.A(_09881_),
    .B(_09883_),
    .C(_09885_),
    .X(_09886_));
 sky130_fd_sc_hd__o21ai_2 _23239_ (.A1(_09881_),
    .A2(_09883_),
    .B1(_09885_),
    .Y(_09887_));
 sky130_fd_sc_hd__a32o_2 _23240_ (.A1(_11712_),
    .A2(_09886_),
    .A3(_09887_),
    .B1(\systolic_inst.acc_wires[1][25] ),
    .B2(_11258_),
    .X(_01899_));
 sky130_fd_sc_hd__or2_2 _23241_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][26] ),
    .X(_09888_));
 sky130_fd_sc_hd__nand2_2 _23242_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][26] ),
    .Y(_09889_));
 sky130_fd_sc_hd__nand2_2 _23243_ (.A(_09888_),
    .B(_09889_),
    .Y(_09890_));
 sky130_fd_sc_hd__o21a_2 _23244_ (.A1(\systolic_inst.acc_wires[1][24] ),
    .A2(\systolic_inst.acc_wires[1][25] ),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .X(_09891_));
 sky130_fd_sc_hd__a21o_2 _23245_ (.A1(_09883_),
    .A2(_09885_),
    .B1(_09891_),
    .X(_09892_));
 sky130_fd_sc_hd__xnor2_2 _23246_ (.A(_09890_),
    .B(_09892_),
    .Y(_09893_));
 sky130_fd_sc_hd__a22o_2 _23247_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][26] ),
    .B1(_11712_),
    .B2(_09893_),
    .X(_01900_));
 sky130_fd_sc_hd__xnor2_2 _23248_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][27] ),
    .Y(_09894_));
 sky130_fd_sc_hd__a21bo_2 _23249_ (.A1(_09888_),
    .A2(_09892_),
    .B1_N(_09889_),
    .X(_09895_));
 sky130_fd_sc_hd__xnor2_2 _23250_ (.A(_09894_),
    .B(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__a22o_2 _23251_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][27] ),
    .B1(_11712_),
    .B2(_09896_),
    .X(_01901_));
 sky130_fd_sc_hd__nor2_2 _23252_ (.A(_09890_),
    .B(_09894_),
    .Y(_09897_));
 sky130_fd_sc_hd__o21a_2 _23253_ (.A1(\systolic_inst.acc_wires[1][26] ),
    .A2(\systolic_inst.acc_wires[1][27] ),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .X(_09898_));
 sky130_fd_sc_hd__a311oi_2 _23254_ (.A1(_09883_),
    .A2(_09885_),
    .A3(_09897_),
    .B1(_09898_),
    .C1(_09891_),
    .Y(_09899_));
 sky130_fd_sc_hd__or2_2 _23255_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][28] ),
    .X(_09900_));
 sky130_fd_sc_hd__nand2_2 _23256_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][28] ),
    .Y(_09901_));
 sky130_fd_sc_hd__nand2_2 _23257_ (.A(_09900_),
    .B(_09901_),
    .Y(_09902_));
 sky130_fd_sc_hd__xor2_2 _23258_ (.A(_09899_),
    .B(_09902_),
    .X(_09903_));
 sky130_fd_sc_hd__a22o_2 _23259_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][28] ),
    .B1(_11712_),
    .B2(_09903_),
    .X(_01902_));
 sky130_fd_sc_hd__xor2_2 _23260_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][29] ),
    .X(_09904_));
 sky130_fd_sc_hd__inv_2 _23261_ (.A(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__o21a_2 _23262_ (.A1(_09899_),
    .A2(_09902_),
    .B1(_09901_),
    .X(_09906_));
 sky130_fd_sc_hd__xnor2_2 _23263_ (.A(_09904_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__a22o_2 _23264_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[1][29] ),
    .B1(_11712_),
    .B2(_09907_),
    .X(_01903_));
 sky130_fd_sc_hd__o21ai_2 _23265_ (.A1(\systolic_inst.acc_wires[1][28] ),
    .A2(\systolic_inst.acc_wires[1][29] ),
    .B1(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .Y(_09908_));
 sky130_fd_sc_hd__o31a_2 _23266_ (.A1(_09899_),
    .A2(_09902_),
    .A3(_09905_),
    .B1(_09908_),
    .X(_09909_));
 sky130_fd_sc_hd__nand2_2 _23267_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][30] ),
    .Y(_09910_));
 sky130_fd_sc_hd__or2_2 _23268_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][30] ),
    .X(_09911_));
 sky130_fd_sc_hd__nand2_2 _23269_ (.A(_09910_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__nand2_2 _23270_ (.A(_09909_),
    .B(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__or2_2 _23271_ (.A(_09909_),
    .B(_09912_),
    .X(_09914_));
 sky130_fd_sc_hd__a32o_2 _23272_ (.A1(_11712_),
    .A2(_09913_),
    .A3(_09914_),
    .B1(\systolic_inst.acc_wires[1][30] ),
    .B2(_11258_),
    .X(_01904_));
 sky130_fd_sc_hd__xnor2_2 _23273_ (.A(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[1][31] ),
    .Y(_09915_));
 sky130_fd_sc_hd__a21oi_2 _23274_ (.A1(_09910_),
    .A2(_09914_),
    .B1(_09915_),
    .Y(_09916_));
 sky130_fd_sc_hd__a31o_2 _23275_ (.A1(_09910_),
    .A2(_09914_),
    .A3(_09915_),
    .B1(_11713_),
    .X(_09917_));
 sky130_fd_sc_hd__a2bb2o_2 _23276_ (.A1_N(_09917_),
    .A2_N(_09916_),
    .B1(\systolic_inst.acc_wires[1][31] ),
    .B2(_11258_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _23277_ (.A0(\systolic_inst.A_outs[0][0] ),
    .A1(\systolic_inst.A_shift[0][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _23278_ (.A0(\systolic_inst.A_outs[0][1] ),
    .A1(\systolic_inst.A_shift[0][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _23279_ (.A0(\systolic_inst.A_outs[0][2] ),
    .A1(\systolic_inst.A_shift[0][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _23280_ (.A0(\systolic_inst.A_outs[0][3] ),
    .A1(\systolic_inst.A_shift[0][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _23281_ (.A0(\systolic_inst.A_outs[0][4] ),
    .A1(\systolic_inst.A_shift[0][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _23282_ (.A0(\systolic_inst.A_outs[0][5] ),
    .A1(\systolic_inst.A_shift[0][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _23283_ (.A0(\systolic_inst.A_outs[0][6] ),
    .A1(\systolic_inst.A_shift[0][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _23284_ (.A0(\systolic_inst.A_outs[0][7] ),
    .A1(\systolic_inst.A_shift[0][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_01913_));
 sky130_fd_sc_hd__and3_2 _23285_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.B_outs[0][0] ),
    .C(\systolic_inst.A_outs[0][0] ),
    .X(_09918_));
 sky130_fd_sc_hd__a21o_2 _23286_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[0] ),
    .B1(_09918_),
    .X(_01914_));
 sky130_fd_sc_hd__and4_2 _23287_ (.A(\systolic_inst.B_outs[0][0] ),
    .B(\systolic_inst.A_outs[0][0] ),
    .C(\systolic_inst.B_outs[0][1] ),
    .D(\systolic_inst.A_outs[0][1] ),
    .X(_09919_));
 sky130_fd_sc_hd__a22o_2 _23288_ (.A1(\systolic_inst.A_outs[0][0] ),
    .A2(\systolic_inst.B_outs[0][1] ),
    .B1(\systolic_inst.A_outs[0][1] ),
    .B2(\systolic_inst.B_outs[0][0] ),
    .X(_09920_));
 sky130_fd_sc_hd__nand2_2 _23289_ (.A(\systolic_inst.ce_local ),
    .B(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__a2bb2o_2 _23290_ (.A1_N(_09921_),
    .A2_N(_09919_),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[1] ),
    .B2(_11258_),
    .X(_01915_));
 sky130_fd_sc_hd__a22o_2 _23291_ (.A1(\systolic_inst.B_outs[0][1] ),
    .A2(\systolic_inst.A_outs[0][1] ),
    .B1(\systolic_inst.B_outs[0][2] ),
    .B2(\systolic_inst.A_outs[0][0] ),
    .X(_09922_));
 sky130_fd_sc_hd__nand4_2 _23292_ (.A(\systolic_inst.A_outs[0][0] ),
    .B(\systolic_inst.B_outs[0][1] ),
    .C(\systolic_inst.A_outs[0][1] ),
    .D(\systolic_inst.B_outs[0][2] ),
    .Y(_09923_));
 sky130_fd_sc_hd__and4_2 _23293_ (.A(\systolic_inst.B_outs[0][0] ),
    .B(\systolic_inst.A_outs[0][2] ),
    .C(_09922_),
    .D(_09923_),
    .X(_09924_));
 sky130_fd_sc_hd__inv_2 _23294_ (.A(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__a22oi_2 _23295_ (.A1(\systolic_inst.B_outs[0][0] ),
    .A2(\systolic_inst.A_outs[0][2] ),
    .B1(_09922_),
    .B2(_09923_),
    .Y(_09926_));
 sky130_fd_sc_hd__nor2_2 _23296_ (.A(_09924_),
    .B(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__xor2_2 _23297_ (.A(_09919_),
    .B(_09927_),
    .X(_09928_));
 sky130_fd_sc_hd__mux2_1 _23298_ (.A0(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[2] ),
    .A1(_09928_),
    .S(\systolic_inst.ce_local ),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_2 _23299_ (.A(\systolic_inst.A_outs[0][0] ),
    .B(\systolic_inst.B_outs[0][3] ),
    .Y(_09929_));
 sky130_fd_sc_hd__a22o_2 _23300_ (.A1(\systolic_inst.A_outs[0][1] ),
    .A2(\systolic_inst.B_outs[0][2] ),
    .B1(\systolic_inst.A_outs[0][2] ),
    .B2(\systolic_inst.B_outs[0][1] ),
    .X(_09930_));
 sky130_fd_sc_hd__nand4_2 _23301_ (.A(\systolic_inst.B_outs[0][1] ),
    .B(\systolic_inst.A_outs[0][1] ),
    .C(\systolic_inst.B_outs[0][2] ),
    .D(\systolic_inst.A_outs[0][2] ),
    .Y(_09931_));
 sky130_fd_sc_hd__and3b_2 _23302_ (.A_N(_09923_),
    .B(_09930_),
    .C(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__a21bo_2 _23303_ (.A1(_09930_),
    .A2(_09931_),
    .B1_N(_09923_),
    .X(_09933_));
 sky130_fd_sc_hd__and2b_2 _23304_ (.A_N(_09932_),
    .B(_09933_),
    .X(_09934_));
 sky130_fd_sc_hd__xnor2_2 _23305_ (.A(_09929_),
    .B(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_2 _23306_ (.A(\systolic_inst.B_outs[0][0] ),
    .B(\systolic_inst.A_outs[0][3] ),
    .Y(_09936_));
 sky130_fd_sc_hd__and3_2 _23307_ (.A(\systolic_inst.B_outs[0][0] ),
    .B(\systolic_inst.A_outs[0][3] ),
    .C(_09935_),
    .X(_09937_));
 sky130_fd_sc_hd__xor2_2 _23308_ (.A(_09935_),
    .B(_09936_),
    .X(_09938_));
 sky130_fd_sc_hd__or2_2 _23309_ (.A(_09925_),
    .B(_09938_),
    .X(_09939_));
 sky130_fd_sc_hd__nand2_2 _23310_ (.A(_09925_),
    .B(_09938_),
    .Y(_09940_));
 sky130_fd_sc_hd__or4b_2 _23311_ (.A(_09924_),
    .B(_09926_),
    .C(_09938_),
    .D_N(_09919_),
    .X(_09941_));
 sky130_fd_sc_hd__a22o_2 _23312_ (.A1(_09919_),
    .A2(_09927_),
    .B1(_09939_),
    .B2(_09940_),
    .X(_09942_));
 sky130_fd_sc_hd__and2_2 _23313_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[3] ),
    .X(_09943_));
 sky130_fd_sc_hd__a31o_2 _23314_ (.A1(\systolic_inst.ce_local ),
    .A2(_09941_),
    .A3(_09942_),
    .B1(_09943_),
    .X(_01917_));
 sky130_fd_sc_hd__nand2_2 _23315_ (.A(\systolic_inst.B_outs[0][0] ),
    .B(\systolic_inst.A_outs[0][4] ),
    .Y(_09944_));
 sky130_fd_sc_hd__a22o_2 _23316_ (.A1(\systolic_inst.A_outs[0][1] ),
    .A2(\systolic_inst.B_outs[0][3] ),
    .B1(\systolic_inst.B_outs[0][4] ),
    .B2(\systolic_inst.A_outs[0][0] ),
    .X(_09945_));
 sky130_fd_sc_hd__nand2_2 _23317_ (.A(\systolic_inst.A_outs[0][1] ),
    .B(\systolic_inst.B_outs[0][4] ),
    .Y(_09946_));
 sky130_fd_sc_hd__or2_2 _23318_ (.A(_09929_),
    .B(_09946_),
    .X(_09947_));
 sky130_fd_sc_hd__a22o_2 _23319_ (.A1(\systolic_inst.B_outs[0][2] ),
    .A2(\systolic_inst.A_outs[0][2] ),
    .B1(\systolic_inst.A_outs[0][3] ),
    .B2(\systolic_inst.B_outs[0][1] ),
    .X(_09948_));
 sky130_fd_sc_hd__nand4_2 _23320_ (.A(\systolic_inst.B_outs[0][1] ),
    .B(\systolic_inst.B_outs[0][2] ),
    .C(\systolic_inst.A_outs[0][2] ),
    .D(\systolic_inst.A_outs[0][3] ),
    .Y(_09949_));
 sky130_fd_sc_hd__nand3b_2 _23321_ (.A_N(_09931_),
    .B(_09948_),
    .C(_09949_),
    .Y(_09950_));
 sky130_fd_sc_hd__a21bo_2 _23322_ (.A1(_09948_),
    .A2(_09949_),
    .B1_N(_09931_),
    .X(_09951_));
 sky130_fd_sc_hd__nand4_2 _23323_ (.A(_09945_),
    .B(_09947_),
    .C(_09950_),
    .D(_09951_),
    .Y(_09952_));
 sky130_fd_sc_hd__a22o_2 _23324_ (.A1(_09945_),
    .A2(_09947_),
    .B1(_09950_),
    .B2(_09951_),
    .X(_09953_));
 sky130_fd_sc_hd__a31o_2 _23325_ (.A1(\systolic_inst.A_outs[0][0] ),
    .A2(\systolic_inst.B_outs[0][3] ),
    .A3(_09933_),
    .B1(_09932_),
    .X(_09954_));
 sky130_fd_sc_hd__and3_2 _23326_ (.A(_09952_),
    .B(_09953_),
    .C(_09954_),
    .X(_09955_));
 sky130_fd_sc_hd__a21oi_2 _23327_ (.A1(_09952_),
    .A2(_09953_),
    .B1(_09954_),
    .Y(_09956_));
 sky130_fd_sc_hd__or3_2 _23328_ (.A(_09944_),
    .B(_09955_),
    .C(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__o21ai_2 _23329_ (.A1(_09955_),
    .A2(_09956_),
    .B1(_09944_),
    .Y(_09958_));
 sky130_fd_sc_hd__and3_2 _23330_ (.A(_09937_),
    .B(_09957_),
    .C(_09958_),
    .X(_09959_));
 sky130_fd_sc_hd__a21oi_2 _23331_ (.A1(_09957_),
    .A2(_09958_),
    .B1(_09937_),
    .Y(_09960_));
 sky130_fd_sc_hd__nor2_2 _23332_ (.A(_09959_),
    .B(_09960_),
    .Y(_09961_));
 sky130_fd_sc_hd__xor2_2 _23333_ (.A(_09939_),
    .B(_09961_),
    .X(_09962_));
 sky130_fd_sc_hd__mux2_1 _23334_ (.A0(_09961_),
    .A1(_09962_),
    .S(_09941_),
    .X(_09963_));
 sky130_fd_sc_hd__inv_2 _23335_ (.A(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__mux2_1 _23336_ (.A0(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[4] ),
    .A1(_09964_),
    .S(\systolic_inst.ce_local ),
    .X(_01918_));
 sky130_fd_sc_hd__a211o_2 _23337_ (.A1(_09939_),
    .A2(_09941_),
    .B1(_09959_),
    .C1(_09960_),
    .X(_09965_));
 sky130_fd_sc_hd__nand4_2 _23338_ (.A(\systolic_inst.B_outs[0][0] ),
    .B(\systolic_inst.A_outs[0][0] ),
    .C(\systolic_inst.B_outs[0][5] ),
    .D(\systolic_inst.A_outs[0][5] ),
    .Y(_09966_));
 sky130_fd_sc_hd__a22o_2 _23339_ (.A1(\systolic_inst.A_outs[0][0] ),
    .A2(\systolic_inst.B_outs[0][5] ),
    .B1(\systolic_inst.A_outs[0][5] ),
    .B2(\systolic_inst.B_outs[0][0] ),
    .X(_09967_));
 sky130_fd_sc_hd__nand3b_2 _23340_ (.A_N(_09947_),
    .B(_09966_),
    .C(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__a21bo_2 _23341_ (.A1(_09966_),
    .A2(_09967_),
    .B1_N(_09947_),
    .X(_09969_));
 sky130_fd_sc_hd__nand2_2 _23342_ (.A(_09968_),
    .B(_09969_),
    .Y(_09970_));
 sky130_fd_sc_hd__nand2_2 _23343_ (.A(\systolic_inst.A_outs[0][2] ),
    .B(\systolic_inst.B_outs[0][3] ),
    .Y(_09971_));
 sky130_fd_sc_hd__and4_2 _23344_ (.A(\systolic_inst.A_outs[0][1] ),
    .B(\systolic_inst.A_outs[0][2] ),
    .C(\systolic_inst.B_outs[0][3] ),
    .D(\systolic_inst.B_outs[0][4] ),
    .X(_09972_));
 sky130_fd_sc_hd__a21o_2 _23345_ (.A1(_09946_),
    .A2(_09971_),
    .B1(_09972_),
    .X(_09973_));
 sky130_fd_sc_hd__a22oi_2 _23346_ (.A1(\systolic_inst.B_outs[0][2] ),
    .A2(\systolic_inst.A_outs[0][3] ),
    .B1(\systolic_inst.A_outs[0][4] ),
    .B2(\systolic_inst.B_outs[0][1] ),
    .Y(_09974_));
 sky130_fd_sc_hd__and4_2 _23347_ (.A(\systolic_inst.B_outs[0][1] ),
    .B(\systolic_inst.B_outs[0][2] ),
    .C(\systolic_inst.A_outs[0][3] ),
    .D(\systolic_inst.A_outs[0][4] ),
    .X(_09975_));
 sky130_fd_sc_hd__nor3_2 _23348_ (.A(_09949_),
    .B(_09974_),
    .C(_09975_),
    .Y(_09976_));
 sky130_fd_sc_hd__o21a_2 _23349_ (.A1(_09974_),
    .A2(_09975_),
    .B1(_09949_),
    .X(_09977_));
 sky130_fd_sc_hd__nor2_2 _23350_ (.A(_09976_),
    .B(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__xnor2_2 _23351_ (.A(_09973_),
    .B(_09978_),
    .Y(_09979_));
 sky130_fd_sc_hd__nand2_2 _23352_ (.A(_09950_),
    .B(_09952_),
    .Y(_09980_));
 sky130_fd_sc_hd__xor2_2 _23353_ (.A(_09979_),
    .B(_09980_),
    .X(_09981_));
 sky130_fd_sc_hd__xor2_2 _23354_ (.A(_09970_),
    .B(_09981_),
    .X(_09982_));
 sky130_fd_sc_hd__nand2b_2 _23355_ (.A_N(_09955_),
    .B(_09957_),
    .Y(_09983_));
 sky130_fd_sc_hd__nand2b_2 _23356_ (.A_N(_09982_),
    .B(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__xnor2_2 _23357_ (.A(_09982_),
    .B(_09983_),
    .Y(_09985_));
 sky130_fd_sc_hd__nand2b_2 _23358_ (.A_N(_09965_),
    .B(_09985_),
    .Y(_09986_));
 sky130_fd_sc_hd__xnor2_2 _23359_ (.A(_09965_),
    .B(_09985_),
    .Y(_09987_));
 sky130_fd_sc_hd__nand2_2 _23360_ (.A(_09959_),
    .B(_09987_),
    .Y(_09988_));
 sky130_fd_sc_hd__xor2_2 _23361_ (.A(_09959_),
    .B(_09987_),
    .X(_09989_));
 sky130_fd_sc_hd__mux2_1 _23362_ (.A0(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[5] ),
    .A1(_09989_),
    .S(\systolic_inst.ce_local ),
    .X(_01919_));
 sky130_fd_sc_hd__a22oi_2 _23363_ (.A1(\systolic_inst.A_outs[0][1] ),
    .A2(\systolic_inst.B_outs[0][5] ),
    .B1(\systolic_inst.A_outs[0][6] ),
    .B2(\systolic_inst.B_outs[0][0] ),
    .Y(_09990_));
 sky130_fd_sc_hd__and4_2 _23364_ (.A(\systolic_inst.B_outs[0][0] ),
    .B(\systolic_inst.A_outs[0][1] ),
    .C(\systolic_inst.B_outs[0][5] ),
    .D(\systolic_inst.A_outs[0][6] ),
    .X(_09991_));
 sky130_fd_sc_hd__nor2_2 _23365_ (.A(_09990_),
    .B(_09991_),
    .Y(_09992_));
 sky130_fd_sc_hd__nand2_2 _23366_ (.A(_09972_),
    .B(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__xnor2_2 _23367_ (.A(_09972_),
    .B(_09992_),
    .Y(_09994_));
 sky130_fd_sc_hd__nand2_2 _23368_ (.A(_09966_),
    .B(_09994_),
    .Y(_09995_));
 sky130_fd_sc_hd__or2_2 _23369_ (.A(_09966_),
    .B(_09994_),
    .X(_09996_));
 sky130_fd_sc_hd__nand2_2 _23370_ (.A(_09995_),
    .B(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__nand2_2 _23371_ (.A(\systolic_inst.A_outs[0][0] ),
    .B(\systolic_inst.B_outs[0][6] ),
    .Y(_09998_));
 sky130_fd_sc_hd__and4_2 _23372_ (.A(\systolic_inst.A_outs[0][2] ),
    .B(\systolic_inst.B_outs[0][3] ),
    .C(\systolic_inst.A_outs[0][3] ),
    .D(\systolic_inst.B_outs[0][4] ),
    .X(_09999_));
 sky130_fd_sc_hd__a22oi_2 _23373_ (.A1(\systolic_inst.B_outs[0][3] ),
    .A2(\systolic_inst.A_outs[0][3] ),
    .B1(\systolic_inst.B_outs[0][4] ),
    .B2(\systolic_inst.A_outs[0][2] ),
    .Y(_10000_));
 sky130_fd_sc_hd__or2_2 _23374_ (.A(_09999_),
    .B(_10000_),
    .X(_10001_));
 sky130_fd_sc_hd__xor2_2 _23375_ (.A(_09998_),
    .B(_10001_),
    .X(_10002_));
 sky130_fd_sc_hd__a22oi_2 _23376_ (.A1(\systolic_inst.B_outs[0][2] ),
    .A2(\systolic_inst.A_outs[0][4] ),
    .B1(\systolic_inst.A_outs[0][5] ),
    .B2(\systolic_inst.B_outs[0][1] ),
    .Y(_10003_));
 sky130_fd_sc_hd__and4_2 _23377_ (.A(\systolic_inst.B_outs[0][1] ),
    .B(\systolic_inst.B_outs[0][2] ),
    .C(\systolic_inst.A_outs[0][4] ),
    .D(\systolic_inst.A_outs[0][5] ),
    .X(_10004_));
 sky130_fd_sc_hd__or3b_2 _23378_ (.A(_10003_),
    .B(_10004_),
    .C_N(_09975_),
    .X(_10005_));
 sky130_fd_sc_hd__o21bai_2 _23379_ (.A1(_10003_),
    .A2(_10004_),
    .B1_N(_09975_),
    .Y(_10006_));
 sky130_fd_sc_hd__and2_2 _23380_ (.A(_10005_),
    .B(_10006_),
    .X(_10007_));
 sky130_fd_sc_hd__xnor2_2 _23381_ (.A(_10002_),
    .B(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__o21bai_2 _23382_ (.A1(_09973_),
    .A2(_09977_),
    .B1_N(_09976_),
    .Y(_10009_));
 sky130_fd_sc_hd__and2b_2 _23383_ (.A_N(_10008_),
    .B(_10009_),
    .X(_10010_));
 sky130_fd_sc_hd__xor2_2 _23384_ (.A(_10008_),
    .B(_10009_),
    .X(_10011_));
 sky130_fd_sc_hd__nor2_2 _23385_ (.A(_09997_),
    .B(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__xor2_2 _23386_ (.A(_09997_),
    .B(_10011_),
    .X(_10013_));
 sky130_fd_sc_hd__a32o_2 _23387_ (.A1(_09968_),
    .A2(_09969_),
    .A3(_09981_),
    .B1(_09980_),
    .B2(_09979_),
    .X(_10014_));
 sky130_fd_sc_hd__nand2_2 _23388_ (.A(_10013_),
    .B(_10014_),
    .Y(_10015_));
 sky130_fd_sc_hd__xnor2_2 _23389_ (.A(_10013_),
    .B(_10014_),
    .Y(_10016_));
 sky130_fd_sc_hd__or2_2 _23390_ (.A(_09968_),
    .B(_10016_),
    .X(_10017_));
 sky130_fd_sc_hd__xnor2_2 _23391_ (.A(_09968_),
    .B(_10016_),
    .Y(_10018_));
 sky130_fd_sc_hd__nor2_2 _23392_ (.A(_09984_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__xnor2_2 _23393_ (.A(_09984_),
    .B(_10018_),
    .Y(_10020_));
 sky130_fd_sc_hd__a21oi_2 _23394_ (.A1(_09986_),
    .A2(_09988_),
    .B1(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__and3_2 _23395_ (.A(_09986_),
    .B(_09988_),
    .C(_10020_),
    .X(_10022_));
 sky130_fd_sc_hd__nand2_2 _23396_ (.A(_11258_),
    .B(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[6] ),
    .Y(_10023_));
 sky130_fd_sc_hd__o31ai_2 _23397_ (.A1(_11258_),
    .A2(_10021_),
    .A3(_10022_),
    .B1(_10023_),
    .Y(_01920_));
 sky130_fd_sc_hd__o21ba_2 _23398_ (.A1(_09998_),
    .A2(_10001_),
    .B1_N(_09999_),
    .X(_10024_));
 sky130_fd_sc_hd__and2_2 _23399_ (.A(\systolic_inst.B_outs[0][0] ),
    .B(\systolic_inst.A_outs[0][7] ),
    .X(_10025_));
 sky130_fd_sc_hd__a21o_2 _23400_ (.A1(\systolic_inst.A_outs[0][2] ),
    .A2(\systolic_inst.B_outs[0][5] ),
    .B1(_10025_),
    .X(_10026_));
 sky130_fd_sc_hd__nand3_2 _23401_ (.A(\systolic_inst.A_outs[0][2] ),
    .B(\systolic_inst.B_outs[0][5] ),
    .C(_10025_),
    .Y(_10027_));
 sky130_fd_sc_hd__nand2_2 _23402_ (.A(_10026_),
    .B(_10027_),
    .Y(_10028_));
 sky130_fd_sc_hd__xor2_2 _23403_ (.A(\systolic_inst.B_outs[0][7] ),
    .B(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__or2_2 _23404_ (.A(_10024_),
    .B(_10029_),
    .X(_10030_));
 sky130_fd_sc_hd__xor2_2 _23405_ (.A(_10024_),
    .B(_10029_),
    .X(_10031_));
 sky130_fd_sc_hd__nand2_2 _23406_ (.A(_09991_),
    .B(_10031_),
    .Y(_10032_));
 sky130_fd_sc_hd__xnor2_2 _23407_ (.A(_09991_),
    .B(_10031_),
    .Y(_10033_));
 sky130_fd_sc_hd__nand2_2 _23408_ (.A(\systolic_inst.A_outs[0][1] ),
    .B(\systolic_inst.B_outs[0][6] ),
    .Y(_10034_));
 sky130_fd_sc_hd__and4_2 _23409_ (.A(\systolic_inst.B_outs[0][3] ),
    .B(\systolic_inst.A_outs[0][3] ),
    .C(\systolic_inst.B_outs[0][4] ),
    .D(\systolic_inst.A_outs[0][4] ),
    .X(_10035_));
 sky130_fd_sc_hd__a22oi_2 _23410_ (.A1(\systolic_inst.A_outs[0][3] ),
    .A2(\systolic_inst.B_outs[0][4] ),
    .B1(\systolic_inst.A_outs[0][4] ),
    .B2(\systolic_inst.B_outs[0][3] ),
    .Y(_10036_));
 sky130_fd_sc_hd__nor2_2 _23411_ (.A(_10035_),
    .B(_10036_),
    .Y(_10037_));
 sky130_fd_sc_hd__xnor2_2 _23412_ (.A(_10034_),
    .B(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__and2b_2 _23413_ (.A_N(\systolic_inst.A_outs[0][0] ),
    .B(\systolic_inst.B_outs[0][7] ),
    .X(_10039_));
 sky130_fd_sc_hd__and4_2 _23414_ (.A(\systolic_inst.B_outs[0][1] ),
    .B(\systolic_inst.B_outs[0][2] ),
    .C(\systolic_inst.A_outs[0][5] ),
    .D(\systolic_inst.A_outs[0][6] ),
    .X(_10040_));
 sky130_fd_sc_hd__a22oi_2 _23415_ (.A1(\systolic_inst.B_outs[0][2] ),
    .A2(\systolic_inst.A_outs[0][5] ),
    .B1(\systolic_inst.A_outs[0][6] ),
    .B2(\systolic_inst.B_outs[0][1] ),
    .Y(_10041_));
 sky130_fd_sc_hd__nor2_2 _23416_ (.A(_10040_),
    .B(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__xor2_2 _23417_ (.A(_10039_),
    .B(_10042_),
    .X(_10043_));
 sky130_fd_sc_hd__nand2_2 _23418_ (.A(_10004_),
    .B(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__xnor2_2 _23419_ (.A(_10004_),
    .B(_10043_),
    .Y(_10045_));
 sky130_fd_sc_hd__inv_2 _23420_ (.A(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__nand2_2 _23421_ (.A(_10038_),
    .B(_10046_),
    .Y(_10047_));
 sky130_fd_sc_hd__xor2_2 _23422_ (.A(_10038_),
    .B(_10045_),
    .X(_10048_));
 sky130_fd_sc_hd__a21bo_2 _23423_ (.A1(_10002_),
    .A2(_10007_),
    .B1_N(_10005_),
    .X(_10049_));
 sky130_fd_sc_hd__nand2b_2 _23424_ (.A_N(_10048_),
    .B(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__xor2_2 _23425_ (.A(_10048_),
    .B(_10049_),
    .X(_10051_));
 sky130_fd_sc_hd__or2_2 _23426_ (.A(_10033_),
    .B(_10051_),
    .X(_10052_));
 sky130_fd_sc_hd__nand2_2 _23427_ (.A(_10033_),
    .B(_10051_),
    .Y(_10053_));
 sky130_fd_sc_hd__o211a_2 _23428_ (.A1(_10010_),
    .A2(_10012_),
    .B1(_10052_),
    .C1(_10053_),
    .X(_10054_));
 sky130_fd_sc_hd__a211oi_2 _23429_ (.A1(_10052_),
    .A2(_10053_),
    .B1(_10010_),
    .C1(_10012_),
    .Y(_10055_));
 sky130_fd_sc_hd__a211oi_2 _23430_ (.A1(_09993_),
    .A2(_09996_),
    .B1(_10054_),
    .C1(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__o211a_2 _23431_ (.A1(_10054_),
    .A2(_10055_),
    .B1(_09993_),
    .C1(_09996_),
    .X(_10057_));
 sky130_fd_sc_hd__a211oi_2 _23432_ (.A1(_10015_),
    .A2(_10017_),
    .B1(_10056_),
    .C1(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__a211o_2 _23433_ (.A1(_10015_),
    .A2(_10017_),
    .B1(_10056_),
    .C1(_10057_),
    .X(_10059_));
 sky130_fd_sc_hd__o211ai_2 _23434_ (.A1(_10056_),
    .A2(_10057_),
    .B1(_10015_),
    .C1(_10017_),
    .Y(_10060_));
 sky130_fd_sc_hd__o211a_2 _23435_ (.A1(_10019_),
    .A2(_10021_),
    .B1(_10059_),
    .C1(_10060_),
    .X(_10061_));
 sky130_fd_sc_hd__a211o_2 _23436_ (.A1(_10059_),
    .A2(_10060_),
    .B1(_10019_),
    .C1(_10021_),
    .X(_10062_));
 sky130_fd_sc_hd__nand2_2 _23437_ (.A(\systolic_inst.ce_local ),
    .B(_10062_),
    .Y(_10063_));
 sky130_fd_sc_hd__a2bb2o_2 _23438_ (.A1_N(_10063_),
    .A2_N(_10061_),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[7] ),
    .B2(_11258_),
    .X(_01921_));
 sky130_fd_sc_hd__a21boi_2 _23439_ (.A1(\systolic_inst.B_outs[0][7] ),
    .A2(_10026_),
    .B1_N(_10027_),
    .Y(_10064_));
 sky130_fd_sc_hd__o21ba_2 _23440_ (.A1(_10034_),
    .A2(_10036_),
    .B1_N(_10035_),
    .X(_10065_));
 sky130_fd_sc_hd__and3_2 _23441_ (.A(\systolic_inst.A_outs[0][3] ),
    .B(\systolic_inst.B_outs[0][5] ),
    .C(_10025_),
    .X(_10066_));
 sky130_fd_sc_hd__a21oi_2 _23442_ (.A1(\systolic_inst.A_outs[0][3] ),
    .A2(\systolic_inst.B_outs[0][5] ),
    .B1(_10025_),
    .Y(_10067_));
 sky130_fd_sc_hd__nor3_2 _23443_ (.A(_10065_),
    .B(_10066_),
    .C(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__o21a_2 _23444_ (.A1(_10066_),
    .A2(_10067_),
    .B1(_10065_),
    .X(_10069_));
 sky130_fd_sc_hd__nor2_2 _23445_ (.A(_10068_),
    .B(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__and2b_2 _23446_ (.A_N(_10064_),
    .B(_10070_),
    .X(_10071_));
 sky130_fd_sc_hd__xnor2_2 _23447_ (.A(_10064_),
    .B(_10070_),
    .Y(_10072_));
 sky130_fd_sc_hd__nand2_2 _23448_ (.A(\systolic_inst.A_outs[0][2] ),
    .B(\systolic_inst.B_outs[0][6] ),
    .Y(_10073_));
 sky130_fd_sc_hd__and4_2 _23449_ (.A(\systolic_inst.B_outs[0][3] ),
    .B(\systolic_inst.B_outs[0][4] ),
    .C(\systolic_inst.A_outs[0][4] ),
    .D(\systolic_inst.A_outs[0][5] ),
    .X(_10074_));
 sky130_fd_sc_hd__a22oi_2 _23450_ (.A1(\systolic_inst.B_outs[0][4] ),
    .A2(\systolic_inst.A_outs[0][4] ),
    .B1(\systolic_inst.A_outs[0][5] ),
    .B2(\systolic_inst.B_outs[0][3] ),
    .Y(_10075_));
 sky130_fd_sc_hd__nor2_2 _23451_ (.A(_10074_),
    .B(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__xnor2_2 _23452_ (.A(_10073_),
    .B(_10076_),
    .Y(_10077_));
 sky130_fd_sc_hd__nand2b_2 _23453_ (.A_N(\systolic_inst.A_outs[0][1] ),
    .B(\systolic_inst.B_outs[0][7] ),
    .Y(_10078_));
 sky130_fd_sc_hd__a22oi_2 _23454_ (.A1(\systolic_inst.B_outs[0][2] ),
    .A2(\systolic_inst.A_outs[0][6] ),
    .B1(\systolic_inst.A_outs[0][7] ),
    .B2(\systolic_inst.B_outs[0][1] ),
    .Y(_10079_));
 sky130_fd_sc_hd__and3_2 _23455_ (.A(\systolic_inst.B_outs[0][1] ),
    .B(\systolic_inst.B_outs[0][2] ),
    .C(\systolic_inst.A_outs[0][7] ),
    .X(_10080_));
 sky130_fd_sc_hd__a21oi_2 _23456_ (.A1(\systolic_inst.A_outs[0][6] ),
    .A2(_10080_),
    .B1(_10079_),
    .Y(_10081_));
 sky130_fd_sc_hd__xnor2_2 _23457_ (.A(_10078_),
    .B(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__a21oi_2 _23458_ (.A1(_10039_),
    .A2(_10042_),
    .B1(_10040_),
    .Y(_10083_));
 sky130_fd_sc_hd__nand2b_2 _23459_ (.A_N(_10083_),
    .B(_10082_),
    .Y(_10084_));
 sky130_fd_sc_hd__xnor2_2 _23460_ (.A(_10082_),
    .B(_10083_),
    .Y(_10085_));
 sky130_fd_sc_hd__nand2_2 _23461_ (.A(_10077_),
    .B(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__or2_2 _23462_ (.A(_10077_),
    .B(_10085_),
    .X(_10087_));
 sky130_fd_sc_hd__nand2_2 _23463_ (.A(_10086_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__a21o_2 _23464_ (.A1(_10044_),
    .A2(_10047_),
    .B1(_10088_),
    .X(_10089_));
 sky130_fd_sc_hd__nand3_2 _23465_ (.A(_10044_),
    .B(_10047_),
    .C(_10088_),
    .Y(_10090_));
 sky130_fd_sc_hd__and3_2 _23466_ (.A(_10072_),
    .B(_10089_),
    .C(_10090_),
    .X(_10091_));
 sky130_fd_sc_hd__nand3_2 _23467_ (.A(_10072_),
    .B(_10089_),
    .C(_10090_),
    .Y(_10092_));
 sky130_fd_sc_hd__a21oi_2 _23468_ (.A1(_10089_),
    .A2(_10090_),
    .B1(_10072_),
    .Y(_10093_));
 sky130_fd_sc_hd__a211oi_2 _23469_ (.A1(_10050_),
    .A2(_10052_),
    .B1(_10091_),
    .C1(_10093_),
    .Y(_10094_));
 sky130_fd_sc_hd__o211a_2 _23470_ (.A1(_10091_),
    .A2(_10093_),
    .B1(_10050_),
    .C1(_10052_),
    .X(_10095_));
 sky130_fd_sc_hd__a211oi_2 _23471_ (.A1(_10030_),
    .A2(_10032_),
    .B1(_10094_),
    .C1(_10095_),
    .Y(_10096_));
 sky130_fd_sc_hd__a211o_2 _23472_ (.A1(_10030_),
    .A2(_10032_),
    .B1(_10094_),
    .C1(_10095_),
    .X(_10097_));
 sky130_fd_sc_hd__o211ai_2 _23473_ (.A1(_10094_),
    .A2(_10095_),
    .B1(_10030_),
    .C1(_10032_),
    .Y(_10098_));
 sky130_fd_sc_hd__o211a_2 _23474_ (.A1(_10054_),
    .A2(_10056_),
    .B1(_10097_),
    .C1(_10098_),
    .X(_10099_));
 sky130_fd_sc_hd__o211ai_2 _23475_ (.A1(_10054_),
    .A2(_10056_),
    .B1(_10097_),
    .C1(_10098_),
    .Y(_10100_));
 sky130_fd_sc_hd__a211o_2 _23476_ (.A1(_10097_),
    .A2(_10098_),
    .B1(_10054_),
    .C1(_10056_),
    .X(_10101_));
 sky130_fd_sc_hd__o211a_2 _23477_ (.A1(_10058_),
    .A2(_10061_),
    .B1(_10100_),
    .C1(_10101_),
    .X(_10102_));
 sky130_fd_sc_hd__a211o_2 _23478_ (.A1(_10100_),
    .A2(_10101_),
    .B1(_10058_),
    .C1(_10061_),
    .X(_10103_));
 sky130_fd_sc_hd__and3b_2 _23479_ (.A_N(_10102_),
    .B(_10103_),
    .C(\systolic_inst.ce_local ),
    .X(_10104_));
 sky130_fd_sc_hd__a21o_2 _23480_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[8] ),
    .B1(_10104_),
    .X(_01922_));
 sky130_fd_sc_hd__o21ba_2 _23481_ (.A1(_10073_),
    .A2(_10075_),
    .B1_N(_10074_),
    .X(_10105_));
 sky130_fd_sc_hd__and3_2 _23482_ (.A(\systolic_inst.A_outs[0][4] ),
    .B(\systolic_inst.B_outs[0][5] ),
    .C(_10025_),
    .X(_10106_));
 sky130_fd_sc_hd__a21oi_2 _23483_ (.A1(\systolic_inst.A_outs[0][4] ),
    .A2(\systolic_inst.B_outs[0][5] ),
    .B1(_10025_),
    .Y(_10107_));
 sky130_fd_sc_hd__nor2_2 _23484_ (.A(_10106_),
    .B(_10107_),
    .Y(_10108_));
 sky130_fd_sc_hd__or3_2 _23485_ (.A(_10105_),
    .B(_10106_),
    .C(_10107_),
    .X(_10109_));
 sky130_fd_sc_hd__xnor2_2 _23486_ (.A(_10105_),
    .B(_10108_),
    .Y(_10110_));
 sky130_fd_sc_hd__nand2_2 _23487_ (.A(_10066_),
    .B(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__or2_2 _23488_ (.A(_10066_),
    .B(_10110_),
    .X(_10112_));
 sky130_fd_sc_hd__nand2_2 _23489_ (.A(_10111_),
    .B(_10112_),
    .Y(_10113_));
 sky130_fd_sc_hd__nand2_2 _23490_ (.A(\systolic_inst.A_outs[0][3] ),
    .B(\systolic_inst.B_outs[0][6] ),
    .Y(_10114_));
 sky130_fd_sc_hd__and4_2 _23491_ (.A(\systolic_inst.B_outs[0][3] ),
    .B(\systolic_inst.B_outs[0][4] ),
    .C(\systolic_inst.A_outs[0][5] ),
    .D(\systolic_inst.A_outs[0][6] ),
    .X(_10115_));
 sky130_fd_sc_hd__a22oi_2 _23492_ (.A1(\systolic_inst.B_outs[0][4] ),
    .A2(\systolic_inst.A_outs[0][5] ),
    .B1(\systolic_inst.A_outs[0][6] ),
    .B2(\systolic_inst.B_outs[0][3] ),
    .Y(_10116_));
 sky130_fd_sc_hd__or2_2 _23493_ (.A(_10115_),
    .B(_10116_),
    .X(_10117_));
 sky130_fd_sc_hd__xor2_2 _23494_ (.A(_10114_),
    .B(_10117_),
    .X(_10118_));
 sky130_fd_sc_hd__o21ai_2 _23495_ (.A1(\systolic_inst.B_outs[0][1] ),
    .A2(\systolic_inst.B_outs[0][2] ),
    .B1(\systolic_inst.A_outs[0][7] ),
    .Y(_10119_));
 sky130_fd_sc_hd__nor2_2 _23496_ (.A(_10080_),
    .B(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__a21oi_2 _23497_ (.A1(_11266_),
    .A2(\systolic_inst.B_outs[0][7] ),
    .B1(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__and3_2 _23498_ (.A(_11266_),
    .B(\systolic_inst.B_outs[0][7] ),
    .C(_10120_),
    .X(_10122_));
 sky130_fd_sc_hd__or2_2 _23499_ (.A(_10121_),
    .B(_10122_),
    .X(_10123_));
 sky130_fd_sc_hd__o2bb2a_2 _23500_ (.A1_N(\systolic_inst.A_outs[0][6] ),
    .A2_N(_10080_),
    .B1(_10079_),
    .B2(_10078_),
    .X(_10124_));
 sky130_fd_sc_hd__or2_2 _23501_ (.A(_10123_),
    .B(_10124_),
    .X(_10125_));
 sky130_fd_sc_hd__xnor2_2 _23502_ (.A(_10123_),
    .B(_10124_),
    .Y(_10126_));
 sky130_fd_sc_hd__inv_2 _23503_ (.A(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__nand2_2 _23504_ (.A(_10118_),
    .B(_10127_),
    .Y(_10128_));
 sky130_fd_sc_hd__xor2_2 _23505_ (.A(_10118_),
    .B(_10126_),
    .X(_10129_));
 sky130_fd_sc_hd__a21oi_2 _23506_ (.A1(_10084_),
    .A2(_10086_),
    .B1(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__and3_2 _23507_ (.A(_10084_),
    .B(_10086_),
    .C(_10129_),
    .X(_10131_));
 sky130_fd_sc_hd__nor3_2 _23508_ (.A(_10113_),
    .B(_10130_),
    .C(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__o21a_2 _23509_ (.A1(_10130_),
    .A2(_10131_),
    .B1(_10113_),
    .X(_10133_));
 sky130_fd_sc_hd__a211o_2 _23510_ (.A1(_10089_),
    .A2(_10092_),
    .B1(_10132_),
    .C1(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__o211ai_2 _23511_ (.A1(_10132_),
    .A2(_10133_),
    .B1(_10089_),
    .C1(_10092_),
    .Y(_10135_));
 sky130_fd_sc_hd__o211ai_2 _23512_ (.A1(_10068_),
    .A2(_10071_),
    .B1(_10134_),
    .C1(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__a211o_2 _23513_ (.A1(_10134_),
    .A2(_10135_),
    .B1(_10068_),
    .C1(_10071_),
    .X(_10137_));
 sky130_fd_sc_hd__o211a_2 _23514_ (.A1(_10094_),
    .A2(_10096_),
    .B1(_10136_),
    .C1(_10137_),
    .X(_10138_));
 sky130_fd_sc_hd__a211o_2 _23515_ (.A1(_10136_),
    .A2(_10137_),
    .B1(_10094_),
    .C1(_10096_),
    .X(_10139_));
 sky130_fd_sc_hd__and2b_2 _23516_ (.A_N(_10138_),
    .B(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__nor2_2 _23517_ (.A(_10099_),
    .B(_10102_),
    .Y(_10141_));
 sky130_fd_sc_hd__and2_2 _23518_ (.A(_10140_),
    .B(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__o21ai_2 _23519_ (.A1(_10140_),
    .A2(_10141_),
    .B1(\systolic_inst.ce_local ),
    .Y(_10143_));
 sky130_fd_sc_hd__o22a_2 _23520_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[9] ),
    .B1(_10142_),
    .B2(_10143_),
    .X(_01923_));
 sky130_fd_sc_hd__o21ba_2 _23521_ (.A1(_10114_),
    .A2(_10116_),
    .B1_N(_10115_),
    .X(_10144_));
 sky130_fd_sc_hd__and3_2 _23522_ (.A(\systolic_inst.B_outs[0][5] ),
    .B(\systolic_inst.A_outs[0][5] ),
    .C(_10025_),
    .X(_10145_));
 sky130_fd_sc_hd__a21oi_2 _23523_ (.A1(\systolic_inst.B_outs[0][5] ),
    .A2(\systolic_inst.A_outs[0][5] ),
    .B1(_10025_),
    .Y(_10146_));
 sky130_fd_sc_hd__or2_2 _23524_ (.A(_10145_),
    .B(_10146_),
    .X(_10147_));
 sky130_fd_sc_hd__or2_2 _23525_ (.A(_10144_),
    .B(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__xor2_2 _23526_ (.A(_10144_),
    .B(_10147_),
    .X(_10149_));
 sky130_fd_sc_hd__or2_2 _23527_ (.A(_10106_),
    .B(_10149_),
    .X(_10150_));
 sky130_fd_sc_hd__nand2_2 _23528_ (.A(_10106_),
    .B(_10149_),
    .Y(_10151_));
 sky130_fd_sc_hd__nand2_2 _23529_ (.A(_10150_),
    .B(_10151_),
    .Y(_10152_));
 sky130_fd_sc_hd__a22oi_2 _23530_ (.A1(\systolic_inst.B_outs[0][4] ),
    .A2(\systolic_inst.A_outs[0][6] ),
    .B1(\systolic_inst.A_outs[0][7] ),
    .B2(\systolic_inst.B_outs[0][3] ),
    .Y(_10153_));
 sky130_fd_sc_hd__and3_2 _23531_ (.A(\systolic_inst.B_outs[0][3] ),
    .B(\systolic_inst.B_outs[0][4] ),
    .C(\systolic_inst.A_outs[0][7] ),
    .X(_10154_));
 sky130_fd_sc_hd__a21oi_2 _23532_ (.A1(\systolic_inst.A_outs[0][6] ),
    .A2(_10154_),
    .B1(_10153_),
    .Y(_10155_));
 sky130_fd_sc_hd__and3_2 _23533_ (.A(\systolic_inst.A_outs[0][4] ),
    .B(\systolic_inst.B_outs[0][6] ),
    .C(_10155_),
    .X(_10156_));
 sky130_fd_sc_hd__a21oi_2 _23534_ (.A1(\systolic_inst.A_outs[0][4] ),
    .A2(\systolic_inst.B_outs[0][6] ),
    .B1(_10155_),
    .Y(_10157_));
 sky130_fd_sc_hd__or2_2 _23535_ (.A(_10156_),
    .B(_10157_),
    .X(_10158_));
 sky130_fd_sc_hd__nand2b_2 _23536_ (.A_N(\systolic_inst.A_outs[0][3] ),
    .B(\systolic_inst.B_outs[0][7] ),
    .Y(_10159_));
 sky130_fd_sc_hd__xnor2_2 _23537_ (.A(_10120_),
    .B(_10159_),
    .Y(_10160_));
 sky130_fd_sc_hd__o21a_2 _23538_ (.A1(_10080_),
    .A2(_10122_),
    .B1(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__nor3_2 _23539_ (.A(_10080_),
    .B(_10122_),
    .C(_10160_),
    .Y(_10162_));
 sky130_fd_sc_hd__or2_2 _23540_ (.A(_10161_),
    .B(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__nor2_2 _23541_ (.A(_10158_),
    .B(_10163_),
    .Y(_10164_));
 sky130_fd_sc_hd__and2_2 _23542_ (.A(_10158_),
    .B(_10163_),
    .X(_10165_));
 sky130_fd_sc_hd__or2_2 _23543_ (.A(_10164_),
    .B(_10165_),
    .X(_10166_));
 sky130_fd_sc_hd__a21oi_2 _23544_ (.A1(_10125_),
    .A2(_10128_),
    .B1(_10166_),
    .Y(_10167_));
 sky130_fd_sc_hd__and3_2 _23545_ (.A(_10125_),
    .B(_10128_),
    .C(_10166_),
    .X(_10168_));
 sky130_fd_sc_hd__or2_2 _23546_ (.A(_10167_),
    .B(_10168_),
    .X(_10169_));
 sky130_fd_sc_hd__nor2_2 _23547_ (.A(_10152_),
    .B(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__xor2_2 _23548_ (.A(_10152_),
    .B(_10169_),
    .X(_10171_));
 sky130_fd_sc_hd__o21a_2 _23549_ (.A1(_10130_),
    .A2(_10132_),
    .B1(_10171_),
    .X(_10172_));
 sky130_fd_sc_hd__o21ai_2 _23550_ (.A1(_10130_),
    .A2(_10132_),
    .B1(_10171_),
    .Y(_10173_));
 sky130_fd_sc_hd__nor3_2 _23551_ (.A(_10130_),
    .B(_10132_),
    .C(_10171_),
    .Y(_10174_));
 sky130_fd_sc_hd__a211oi_2 _23552_ (.A1(_10109_),
    .A2(_10111_),
    .B1(_10172_),
    .C1(_10174_),
    .Y(_10175_));
 sky130_fd_sc_hd__a211o_2 _23553_ (.A1(_10109_),
    .A2(_10111_),
    .B1(_10172_),
    .C1(_10174_),
    .X(_10176_));
 sky130_fd_sc_hd__o211a_2 _23554_ (.A1(_10172_),
    .A2(_10174_),
    .B1(_10109_),
    .C1(_10111_),
    .X(_10177_));
 sky130_fd_sc_hd__a211oi_2 _23555_ (.A1(_10134_),
    .A2(_10136_),
    .B1(_10175_),
    .C1(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__o211a_2 _23556_ (.A1(_10175_),
    .A2(_10177_),
    .B1(_10134_),
    .C1(_10136_),
    .X(_10179_));
 sky130_fd_sc_hd__o31a_2 _23557_ (.A1(_10099_),
    .A2(_10102_),
    .A3(_10138_),
    .B1(_10139_),
    .X(_10180_));
 sky130_fd_sc_hd__o21bai_2 _23558_ (.A1(_10178_),
    .A2(_10179_),
    .B1_N(_10180_),
    .Y(_10181_));
 sky130_fd_sc_hd__nor3b_2 _23559_ (.A(_10178_),
    .B(_10179_),
    .C_N(_10180_),
    .Y(_10182_));
 sky130_fd_sc_hd__nor2_2 _23560_ (.A(_11258_),
    .B(_10182_),
    .Y(_10183_));
 sky130_fd_sc_hd__a22o_2 _23561_ (.A1(_11258_),
    .A2(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[10] ),
    .B1(_10181_),
    .B2(_10183_),
    .X(_01924_));
 sky130_fd_sc_hd__nor2_2 _23562_ (.A(_10178_),
    .B(_10182_),
    .Y(_10184_));
 sky130_fd_sc_hd__a21oi_2 _23563_ (.A1(\systolic_inst.A_outs[0][6] ),
    .A2(_10154_),
    .B1(_10156_),
    .Y(_10185_));
 sky130_fd_sc_hd__and3_2 _23564_ (.A(\systolic_inst.B_outs[0][5] ),
    .B(\systolic_inst.A_outs[0][6] ),
    .C(_10025_),
    .X(_10186_));
 sky130_fd_sc_hd__a21oi_2 _23565_ (.A1(\systolic_inst.B_outs[0][5] ),
    .A2(\systolic_inst.A_outs[0][6] ),
    .B1(_10025_),
    .Y(_10187_));
 sky130_fd_sc_hd__nor2_2 _23566_ (.A(_10186_),
    .B(_10187_),
    .Y(_10188_));
 sky130_fd_sc_hd__and2b_2 _23567_ (.A_N(_10185_),
    .B(_10188_),
    .X(_10189_));
 sky130_fd_sc_hd__xnor2_2 _23568_ (.A(_10185_),
    .B(_10188_),
    .Y(_10190_));
 sky130_fd_sc_hd__xnor2_2 _23569_ (.A(_10145_),
    .B(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__o21ai_2 _23570_ (.A1(\systolic_inst.B_outs[0][3] ),
    .A2(\systolic_inst.B_outs[0][4] ),
    .B1(\systolic_inst.A_outs[0][7] ),
    .Y(_10192_));
 sky130_fd_sc_hd__nor2_2 _23571_ (.A(_10154_),
    .B(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__a21oi_2 _23572_ (.A1(\systolic_inst.A_outs[0][5] ),
    .A2(\systolic_inst.B_outs[0][6] ),
    .B1(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__and2_2 _23573_ (.A(\systolic_inst.B_outs[0][6] ),
    .B(_10193_),
    .X(_10195_));
 sky130_fd_sc_hd__a21o_2 _23574_ (.A1(\systolic_inst.A_outs[0][5] ),
    .A2(_10195_),
    .B1(_10194_),
    .X(_10196_));
 sky130_fd_sc_hd__a21oi_2 _23575_ (.A1(_11267_),
    .A2(\systolic_inst.B_outs[0][7] ),
    .B1(_10120_),
    .Y(_10197_));
 sky130_fd_sc_hd__and3_2 _23576_ (.A(_11267_),
    .B(\systolic_inst.B_outs[0][7] ),
    .C(_10120_),
    .X(_10198_));
 sky130_fd_sc_hd__nor2_2 _23577_ (.A(_10197_),
    .B(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__o21bai_2 _23578_ (.A1(_10119_),
    .A2(_10159_),
    .B1_N(_10080_),
    .Y(_10200_));
 sky130_fd_sc_hd__and2_2 _23579_ (.A(_10199_),
    .B(_10200_),
    .X(_10201_));
 sky130_fd_sc_hd__xnor2_2 _23580_ (.A(_10199_),
    .B(_10200_),
    .Y(_10202_));
 sky130_fd_sc_hd__nor2_2 _23581_ (.A(_10196_),
    .B(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__xor2_2 _23582_ (.A(_10196_),
    .B(_10202_),
    .X(_10204_));
 sky130_fd_sc_hd__o21a_2 _23583_ (.A1(_10161_),
    .A2(_10164_),
    .B1(_10204_),
    .X(_10205_));
 sky130_fd_sc_hd__nor3_2 _23584_ (.A(_10161_),
    .B(_10164_),
    .C(_10204_),
    .Y(_10206_));
 sky130_fd_sc_hd__or2_2 _23585_ (.A(_10205_),
    .B(_10206_),
    .X(_10207_));
 sky130_fd_sc_hd__nor2_2 _23586_ (.A(_10191_),
    .B(_10207_),
    .Y(_10208_));
 sky130_fd_sc_hd__and2_2 _23587_ (.A(_10191_),
    .B(_10207_),
    .X(_10209_));
 sky130_fd_sc_hd__nor2_2 _23588_ (.A(_10208_),
    .B(_10209_),
    .Y(_10210_));
 sky130_fd_sc_hd__o21a_2 _23589_ (.A1(_10167_),
    .A2(_10170_),
    .B1(_10210_),
    .X(_10211_));
 sky130_fd_sc_hd__nor3_2 _23590_ (.A(_10167_),
    .B(_10170_),
    .C(_10210_),
    .Y(_10212_));
 sky130_fd_sc_hd__a211oi_2 _23591_ (.A1(_10148_),
    .A2(_10151_),
    .B1(_10211_),
    .C1(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__o211a_2 _23592_ (.A1(_10211_),
    .A2(_10212_),
    .B1(_10148_),
    .C1(_10151_),
    .X(_10214_));
 sky130_fd_sc_hd__a211oi_2 _23593_ (.A1(_10173_),
    .A2(_10176_),
    .B1(_10213_),
    .C1(_10214_),
    .Y(_10215_));
 sky130_fd_sc_hd__o211a_2 _23594_ (.A1(_10213_),
    .A2(_10214_),
    .B1(_10173_),
    .C1(_10176_),
    .X(_10216_));
 sky130_fd_sc_hd__inv_2 _23595_ (.A(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__nor2_2 _23596_ (.A(_10215_),
    .B(_10216_),
    .Y(_10218_));
 sky130_fd_sc_hd__xnor2_2 _23597_ (.A(_10184_),
    .B(_10218_),
    .Y(_10219_));
 sky130_fd_sc_hd__mux2_1 _23598_ (.A0(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[11] ),
    .A1(_10219_),
    .S(\systolic_inst.ce_local ),
    .X(_01925_));
 sky130_fd_sc_hd__a21o_2 _23599_ (.A1(_10145_),
    .A2(_10190_),
    .B1(_10189_),
    .X(_10220_));
 sky130_fd_sc_hd__a31o_2 _23600_ (.A1(\systolic_inst.A_outs[0][5] ),
    .A2(\systolic_inst.B_outs[0][6] ),
    .A3(_10193_),
    .B1(_10154_),
    .X(_10221_));
 sky130_fd_sc_hd__o21ai_2 _23601_ (.A1(\systolic_inst.B_outs[0][0] ),
    .A2(\systolic_inst.B_outs[0][5] ),
    .B1(\systolic_inst.A_outs[0][7] ),
    .Y(_10222_));
 sky130_fd_sc_hd__a21o_2 _23602_ (.A1(\systolic_inst.B_outs[0][0] ),
    .A2(\systolic_inst.B_outs[0][5] ),
    .B1(_10222_),
    .X(_10223_));
 sky130_fd_sc_hd__nand2b_2 _23603_ (.A_N(_10223_),
    .B(_10221_),
    .Y(_10224_));
 sky130_fd_sc_hd__xnor2_2 _23604_ (.A(_10221_),
    .B(_10223_),
    .Y(_10225_));
 sky130_fd_sc_hd__or2_2 _23605_ (.A(_10186_),
    .B(_10225_),
    .X(_10226_));
 sky130_fd_sc_hd__nand2_2 _23606_ (.A(_10186_),
    .B(_10225_),
    .Y(_10227_));
 sky130_fd_sc_hd__nand2_2 _23607_ (.A(_10226_),
    .B(_10227_),
    .Y(_10228_));
 sky130_fd_sc_hd__a21oi_2 _23608_ (.A1(_11268_),
    .A2(\systolic_inst.B_outs[0][7] ),
    .B1(_10120_),
    .Y(_10229_));
 sky130_fd_sc_hd__and3_2 _23609_ (.A(_11268_),
    .B(\systolic_inst.B_outs[0][7] ),
    .C(_10120_),
    .X(_10230_));
 sky130_fd_sc_hd__nor2_2 _23610_ (.A(_10229_),
    .B(_10230_),
    .Y(_10231_));
 sky130_fd_sc_hd__or2_2 _23611_ (.A(_10080_),
    .B(_10198_),
    .X(_10232_));
 sky130_fd_sc_hd__nand2_2 _23612_ (.A(_10231_),
    .B(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__xnor2_2 _23613_ (.A(_10231_),
    .B(_10232_),
    .Y(_10234_));
 sky130_fd_sc_hd__a21oi_2 _23614_ (.A1(\systolic_inst.B_outs[0][6] ),
    .A2(\systolic_inst.A_outs[0][6] ),
    .B1(_10193_),
    .Y(_10235_));
 sky130_fd_sc_hd__a21o_2 _23615_ (.A1(\systolic_inst.A_outs[0][6] ),
    .A2(_10195_),
    .B1(_10235_),
    .X(_10236_));
 sky130_fd_sc_hd__xor2_2 _23616_ (.A(_10234_),
    .B(_10236_),
    .X(_10237_));
 sky130_fd_sc_hd__o21ai_2 _23617_ (.A1(_10201_),
    .A2(_10203_),
    .B1(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__or3_2 _23618_ (.A(_10201_),
    .B(_10203_),
    .C(_10237_),
    .X(_10239_));
 sky130_fd_sc_hd__nand2_2 _23619_ (.A(_10238_),
    .B(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__or2_2 _23620_ (.A(_10228_),
    .B(_10240_),
    .X(_10241_));
 sky130_fd_sc_hd__nand2_2 _23621_ (.A(_10228_),
    .B(_10240_),
    .Y(_10242_));
 sky130_fd_sc_hd__and2_2 _23622_ (.A(_10241_),
    .B(_10242_),
    .X(_10243_));
 sky130_fd_sc_hd__o21ai_2 _23623_ (.A1(_10205_),
    .A2(_10208_),
    .B1(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__or3_2 _23624_ (.A(_10205_),
    .B(_10208_),
    .C(_10243_),
    .X(_10245_));
 sky130_fd_sc_hd__nand3_2 _23625_ (.A(_10220_),
    .B(_10244_),
    .C(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__a21o_2 _23626_ (.A1(_10244_),
    .A2(_10245_),
    .B1(_10220_),
    .X(_10247_));
 sky130_fd_sc_hd__nand2_2 _23627_ (.A(_10246_),
    .B(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__or2_2 _23628_ (.A(_10211_),
    .B(_10213_),
    .X(_10249_));
 sky130_fd_sc_hd__and3_2 _23629_ (.A(_10246_),
    .B(_10247_),
    .C(_10249_),
    .X(_10250_));
 sky130_fd_sc_hd__xnor2_2 _23630_ (.A(_10248_),
    .B(_10249_),
    .Y(_10251_));
 sky130_fd_sc_hd__o31a_2 _23631_ (.A1(_10178_),
    .A2(_10182_),
    .A3(_10215_),
    .B1(_10217_),
    .X(_10252_));
 sky130_fd_sc_hd__o311a_2 _23632_ (.A1(_10178_),
    .A2(_10182_),
    .A3(_10215_),
    .B1(_10217_),
    .C1(_10251_),
    .X(_10253_));
 sky130_fd_sc_hd__nor2_2 _23633_ (.A(_10251_),
    .B(_10252_),
    .Y(_10254_));
 sky130_fd_sc_hd__nor2_2 _23634_ (.A(_10253_),
    .B(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__mux2_1 _23635_ (.A0(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[12] ),
    .A1(_10255_),
    .S(\systolic_inst.ce_local ),
    .X(_01926_));
 sky130_fd_sc_hd__o21a_2 _23636_ (.A1(_10234_),
    .A2(_10236_),
    .B1(_10233_),
    .X(_10256_));
 sky130_fd_sc_hd__a21oi_2 _23637_ (.A1(_11269_),
    .A2(\systolic_inst.B_outs[0][7] ),
    .B1(_10120_),
    .Y(_10257_));
 sky130_fd_sc_hd__and3_2 _23638_ (.A(_11269_),
    .B(\systolic_inst.B_outs[0][7] ),
    .C(_10120_),
    .X(_10258_));
 sky130_fd_sc_hd__nor2_2 _23639_ (.A(_10257_),
    .B(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__o21a_2 _23640_ (.A1(_10080_),
    .A2(_10230_),
    .B1(_10259_),
    .X(_10260_));
 sky130_fd_sc_hd__or3_2 _23641_ (.A(_10080_),
    .B(_10230_),
    .C(_10259_),
    .X(_10261_));
 sky130_fd_sc_hd__nand2b_2 _23642_ (.A_N(_10260_),
    .B(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__a21oi_2 _23643_ (.A1(\systolic_inst.B_outs[0][6] ),
    .A2(\systolic_inst.A_outs[0][7] ),
    .B1(_10193_),
    .Y(_10263_));
 sky130_fd_sc_hd__or2_2 _23644_ (.A(_10195_),
    .B(_10263_),
    .X(_10264_));
 sky130_fd_sc_hd__xnor2_2 _23645_ (.A(_10262_),
    .B(_10264_),
    .Y(_10265_));
 sky130_fd_sc_hd__nor2_2 _23646_ (.A(_10256_),
    .B(_10265_),
    .Y(_10266_));
 sky130_fd_sc_hd__xnor2_2 _23647_ (.A(_10256_),
    .B(_10265_),
    .Y(_10267_));
 sky130_fd_sc_hd__a21oi_2 _23648_ (.A1(\systolic_inst.A_outs[0][6] ),
    .A2(_10195_),
    .B1(_10154_),
    .Y(_10268_));
 sky130_fd_sc_hd__nor2_2 _23649_ (.A(_10222_),
    .B(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__and2_2 _23650_ (.A(_10222_),
    .B(_10268_),
    .X(_10270_));
 sky130_fd_sc_hd__nor2_2 _23651_ (.A(_10269_),
    .B(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__and2b_2 _23652_ (.A_N(_10267_),
    .B(_10271_),
    .X(_10272_));
 sky130_fd_sc_hd__xor2_2 _23653_ (.A(_10267_),
    .B(_10271_),
    .X(_10273_));
 sky130_fd_sc_hd__a21oi_2 _23654_ (.A1(_10238_),
    .A2(_10241_),
    .B1(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__and3_2 _23655_ (.A(_10238_),
    .B(_10241_),
    .C(_10273_),
    .X(_10275_));
 sky130_fd_sc_hd__a211oi_2 _23656_ (.A1(_10224_),
    .A2(_10227_),
    .B1(_10274_),
    .C1(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__o211a_2 _23657_ (.A1(_10274_),
    .A2(_10275_),
    .B1(_10224_),
    .C1(_10227_),
    .X(_10277_));
 sky130_fd_sc_hd__o211ai_2 _23658_ (.A1(_10276_),
    .A2(_10277_),
    .B1(_10244_),
    .C1(_10246_),
    .Y(_10278_));
 sky130_fd_sc_hd__a211o_2 _23659_ (.A1(_10244_),
    .A2(_10246_),
    .B1(_10276_),
    .C1(_10277_),
    .X(_10279_));
 sky130_fd_sc_hd__and2_2 _23660_ (.A(_10278_),
    .B(_10279_),
    .X(_10280_));
 sky130_fd_sc_hd__nor2_2 _23661_ (.A(_10250_),
    .B(_10253_),
    .Y(_10281_));
 sky130_fd_sc_hd__xnor2_2 _23662_ (.A(_10280_),
    .B(_10281_),
    .Y(_10282_));
 sky130_fd_sc_hd__mux2_1 _23663_ (.A0(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[13] ),
    .A1(_10282_),
    .S(\systolic_inst.ce_local ),
    .X(_01927_));
 sky130_fd_sc_hd__o21bai_2 _23664_ (.A1(_10154_),
    .A2(_10195_),
    .B1_N(_10222_),
    .Y(_10283_));
 sky130_fd_sc_hd__inv_2 _23665_ (.A(_10283_),
    .Y(_10284_));
 sky130_fd_sc_hd__or3b_2 _23666_ (.A(_10154_),
    .B(_10195_),
    .C_N(_10222_),
    .X(_10285_));
 sky130_fd_sc_hd__nand2_2 _23667_ (.A(_10283_),
    .B(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__a21oi_2 _23668_ (.A1(\systolic_inst.B_outs[0][7] ),
    .A2(_11270_),
    .B1(_10120_),
    .Y(_10287_));
 sky130_fd_sc_hd__o21ba_2 _23669_ (.A1(_10258_),
    .A2(_10287_),
    .B1_N(_10080_),
    .X(_10288_));
 sky130_fd_sc_hd__o21a_2 _23670_ (.A1(_10260_),
    .A2(_10288_),
    .B1(_10264_),
    .X(_10289_));
 sky130_fd_sc_hd__a21oi_2 _23671_ (.A1(_10261_),
    .A2(_10288_),
    .B1(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__xnor2_2 _23672_ (.A(_10286_),
    .B(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__o21ai_2 _23673_ (.A1(_10266_),
    .A2(_10272_),
    .B1(_10291_),
    .Y(_10292_));
 sky130_fd_sc_hd__or3_2 _23674_ (.A(_10266_),
    .B(_10272_),
    .C(_10291_),
    .X(_10293_));
 sky130_fd_sc_hd__and2_2 _23675_ (.A(_10292_),
    .B(_10293_),
    .X(_10294_));
 sky130_fd_sc_hd__nand2_2 _23676_ (.A(_10269_),
    .B(_10294_),
    .Y(_10295_));
 sky130_fd_sc_hd__or2_2 _23677_ (.A(_10269_),
    .B(_10294_),
    .X(_10296_));
 sky130_fd_sc_hd__nand2_2 _23678_ (.A(_10295_),
    .B(_10296_),
    .Y(_10297_));
 sky130_fd_sc_hd__nor2_2 _23679_ (.A(_10274_),
    .B(_10276_),
    .Y(_10298_));
 sky130_fd_sc_hd__xnor2_2 _23680_ (.A(_10297_),
    .B(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__a21bo_2 _23681_ (.A1(_10250_),
    .A2(_10278_),
    .B1_N(_10279_),
    .X(_10300_));
 sky130_fd_sc_hd__a21oi_2 _23682_ (.A1(_10253_),
    .A2(_10280_),
    .B1(_10300_),
    .Y(_10301_));
 sky130_fd_sc_hd__nor2_2 _23683_ (.A(_10299_),
    .B(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__xnor2_2 _23684_ (.A(_10299_),
    .B(_10301_),
    .Y(_10303_));
 sky130_fd_sc_hd__nor2_2 _23685_ (.A(\systolic_inst.ce_local ),
    .B(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[14] ),
    .Y(_10304_));
 sky130_fd_sc_hd__a21oi_2 _23686_ (.A1(\systolic_inst.ce_local ),
    .A2(_10303_),
    .B1(_10304_),
    .Y(_01928_));
 sky130_fd_sc_hd__a22o_2 _23687_ (.A1(_10284_),
    .A2(_10290_),
    .B1(_10292_),
    .B2(_10295_),
    .X(_10305_));
 sky130_fd_sc_hd__o221a_2 _23688_ (.A1(_10285_),
    .A2(_10290_),
    .B1(_10297_),
    .B2(_10298_),
    .C1(\systolic_inst.ce_local ),
    .X(_10306_));
 sky130_fd_sc_hd__nand2_2 _23689_ (.A(_10305_),
    .B(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__a2bb2o_2 _23690_ (.A1_N(_10307_),
    .A2_N(_10302_),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B2(_11258_),
    .X(_01929_));
 sky130_fd_sc_hd__a21o_2 _23691_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[0][0] ),
    .B1(\systolic_inst.load_acc ),
    .X(_10308_));
 sky130_fd_sc_hd__a21oi_2 _23692_ (.A1(\systolic_inst.ce_local ),
    .A2(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[0] ),
    .B1(\systolic_inst.acc_wires[0][0] ),
    .Y(_10309_));
 sky130_fd_sc_hd__a21oi_2 _23693_ (.A1(\systolic_inst.ce_local ),
    .A2(_10308_),
    .B1(_10309_),
    .Y(_01930_));
 sky130_fd_sc_hd__and2_2 _23694_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[0][1] ),
    .X(_10310_));
 sky130_fd_sc_hd__nand2_2 _23695_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[0][1] ),
    .Y(_10311_));
 sky130_fd_sc_hd__or2_2 _23696_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[1] ),
    .B(\systolic_inst.acc_wires[0][1] ),
    .X(_10312_));
 sky130_fd_sc_hd__and4_2 _23697_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[0] ),
    .B(\systolic_inst.acc_wires[0][0] ),
    .C(_10311_),
    .D(_10312_),
    .X(_10313_));
 sky130_fd_sc_hd__inv_2 _23698_ (.A(_10313_),
    .Y(_10314_));
 sky130_fd_sc_hd__a22o_2 _23699_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[0][0] ),
    .B1(_10311_),
    .B2(_10312_),
    .X(_10315_));
 sky130_fd_sc_hd__a32o_2 _23700_ (.A1(_11712_),
    .A2(_10314_),
    .A3(_10315_),
    .B1(\systolic_inst.acc_wires[0][1] ),
    .B2(_11258_),
    .X(_01931_));
 sky130_fd_sc_hd__nand2_2 _23701_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[0][2] ),
    .Y(_10316_));
 sky130_fd_sc_hd__or2_2 _23702_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[2] ),
    .B(\systolic_inst.acc_wires[0][2] ),
    .X(_10317_));
 sky130_fd_sc_hd__a31o_2 _23703_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[0] ),
    .A2(\systolic_inst.acc_wires[0][0] ),
    .A3(_10312_),
    .B1(_10310_),
    .X(_10318_));
 sky130_fd_sc_hd__a21o_2 _23704_ (.A1(_10316_),
    .A2(_10317_),
    .B1(_10318_),
    .X(_10319_));
 sky130_fd_sc_hd__and3_2 _23705_ (.A(_10316_),
    .B(_10317_),
    .C(_10318_),
    .X(_10320_));
 sky130_fd_sc_hd__inv_2 _23706_ (.A(_10320_),
    .Y(_10321_));
 sky130_fd_sc_hd__a32o_2 _23707_ (.A1(_11712_),
    .A2(_10319_),
    .A3(_10321_),
    .B1(\systolic_inst.acc_wires[0][2] ),
    .B2(_11258_),
    .X(_01932_));
 sky130_fd_sc_hd__nand2_2 _23708_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[0][3] ),
    .Y(_10322_));
 sky130_fd_sc_hd__or2_2 _23709_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[3] ),
    .B(\systolic_inst.acc_wires[0][3] ),
    .X(_10323_));
 sky130_fd_sc_hd__a21bo_2 _23710_ (.A1(_10317_),
    .A2(_10318_),
    .B1_N(_10316_),
    .X(_10324_));
 sky130_fd_sc_hd__a21o_2 _23711_ (.A1(_10322_),
    .A2(_10323_),
    .B1(_10324_),
    .X(_10325_));
 sky130_fd_sc_hd__and3_2 _23712_ (.A(_10322_),
    .B(_10323_),
    .C(_10324_),
    .X(_10326_));
 sky130_fd_sc_hd__inv_2 _23713_ (.A(_10326_),
    .Y(_10327_));
 sky130_fd_sc_hd__a32o_2 _23714_ (.A1(_11712_),
    .A2(_10325_),
    .A3(_10327_),
    .B1(\systolic_inst.acc_wires[0][3] ),
    .B2(_11258_),
    .X(_01933_));
 sky130_fd_sc_hd__nand2_2 _23715_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[0][4] ),
    .Y(_10328_));
 sky130_fd_sc_hd__or2_2 _23716_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[4] ),
    .B(\systolic_inst.acc_wires[0][4] ),
    .X(_10329_));
 sky130_fd_sc_hd__a21bo_2 _23717_ (.A1(_10323_),
    .A2(_10324_),
    .B1_N(_10322_),
    .X(_10330_));
 sky130_fd_sc_hd__a21o_2 _23718_ (.A1(_10328_),
    .A2(_10329_),
    .B1(_10330_),
    .X(_10331_));
 sky130_fd_sc_hd__and3_2 _23719_ (.A(_10328_),
    .B(_10329_),
    .C(_10330_),
    .X(_10332_));
 sky130_fd_sc_hd__inv_2 _23720_ (.A(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__a32o_2 _23721_ (.A1(_11712_),
    .A2(_10331_),
    .A3(_10333_),
    .B1(\systolic_inst.acc_wires[0][4] ),
    .B2(_11258_),
    .X(_01934_));
 sky130_fd_sc_hd__nand2_2 _23722_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[0][5] ),
    .Y(_10334_));
 sky130_fd_sc_hd__or2_2 _23723_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[5] ),
    .B(\systolic_inst.acc_wires[0][5] ),
    .X(_10335_));
 sky130_fd_sc_hd__a21bo_2 _23724_ (.A1(_10329_),
    .A2(_10330_),
    .B1_N(_10328_),
    .X(_10336_));
 sky130_fd_sc_hd__a21o_2 _23725_ (.A1(_10334_),
    .A2(_10335_),
    .B1(_10336_),
    .X(_10337_));
 sky130_fd_sc_hd__and3_2 _23726_ (.A(_10334_),
    .B(_10335_),
    .C(_10336_),
    .X(_10338_));
 sky130_fd_sc_hd__inv_2 _23727_ (.A(_10338_),
    .Y(_10339_));
 sky130_fd_sc_hd__a32o_2 _23728_ (.A1(_11712_),
    .A2(_10337_),
    .A3(_10339_),
    .B1(\systolic_inst.acc_wires[0][5] ),
    .B2(_11258_),
    .X(_01935_));
 sky130_fd_sc_hd__nand2_2 _23729_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[0][6] ),
    .Y(_10340_));
 sky130_fd_sc_hd__or2_2 _23730_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[6] ),
    .B(\systolic_inst.acc_wires[0][6] ),
    .X(_10341_));
 sky130_fd_sc_hd__a21bo_2 _23731_ (.A1(_10335_),
    .A2(_10336_),
    .B1_N(_10334_),
    .X(_10342_));
 sky130_fd_sc_hd__a21o_2 _23732_ (.A1(_10340_),
    .A2(_10341_),
    .B1(_10342_),
    .X(_10343_));
 sky130_fd_sc_hd__and3_2 _23733_ (.A(_10340_),
    .B(_10341_),
    .C(_10342_),
    .X(_10344_));
 sky130_fd_sc_hd__inv_2 _23734_ (.A(_10344_),
    .Y(_10345_));
 sky130_fd_sc_hd__a32o_2 _23735_ (.A1(_11712_),
    .A2(_10343_),
    .A3(_10345_),
    .B1(\systolic_inst.acc_wires[0][6] ),
    .B2(_11258_),
    .X(_01936_));
 sky130_fd_sc_hd__nand2_2 _23736_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[0][7] ),
    .Y(_10346_));
 sky130_fd_sc_hd__or2_2 _23737_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[7] ),
    .B(\systolic_inst.acc_wires[0][7] ),
    .X(_10347_));
 sky130_fd_sc_hd__a21bo_2 _23738_ (.A1(_10341_),
    .A2(_10342_),
    .B1_N(_10340_),
    .X(_10348_));
 sky130_fd_sc_hd__a21o_2 _23739_ (.A1(_10346_),
    .A2(_10347_),
    .B1(_10348_),
    .X(_10349_));
 sky130_fd_sc_hd__nand3_2 _23740_ (.A(_10346_),
    .B(_10347_),
    .C(_10348_),
    .Y(_10350_));
 sky130_fd_sc_hd__a32o_2 _23741_ (.A1(_11712_),
    .A2(_10349_),
    .A3(_10350_),
    .B1(\systolic_inst.acc_wires[0][7] ),
    .B2(_11258_),
    .X(_01937_));
 sky130_fd_sc_hd__a21bo_2 _23742_ (.A1(_10347_),
    .A2(_10348_),
    .B1_N(_10346_),
    .X(_10351_));
 sky130_fd_sc_hd__xor2_2 _23743_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[0][8] ),
    .X(_10352_));
 sky130_fd_sc_hd__and2_2 _23744_ (.A(_10351_),
    .B(_10352_),
    .X(_10353_));
 sky130_fd_sc_hd__o21ai_2 _23745_ (.A1(_10351_),
    .A2(_10352_),
    .B1(_11712_),
    .Y(_10354_));
 sky130_fd_sc_hd__a2bb2o_2 _23746_ (.A1_N(_10354_),
    .A2_N(_10353_),
    .B1(\systolic_inst.acc_wires[0][8] ),
    .B2(_11258_),
    .X(_01938_));
 sky130_fd_sc_hd__xor2_2 _23747_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[9] ),
    .B(\systolic_inst.acc_wires[0][9] ),
    .X(_10355_));
 sky130_fd_sc_hd__a211o_2 _23748_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[8] ),
    .A2(\systolic_inst.acc_wires[0][8] ),
    .B1(_10353_),
    .C1(_10355_),
    .X(_10356_));
 sky130_fd_sc_hd__nand2_2 _23749_ (.A(_10352_),
    .B(_10355_),
    .Y(_10357_));
 sky130_fd_sc_hd__nand2_2 _23750_ (.A(_10353_),
    .B(_10355_),
    .Y(_10358_));
 sky130_fd_sc_hd__and3_2 _23751_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[8] ),
    .B(\systolic_inst.acc_wires[0][8] ),
    .C(_10355_),
    .X(_10359_));
 sky130_fd_sc_hd__nor2_2 _23752_ (.A(_11713_),
    .B(_10359_),
    .Y(_10360_));
 sky130_fd_sc_hd__a32o_2 _23753_ (.A1(_10356_),
    .A2(_10358_),
    .A3(_10360_),
    .B1(\systolic_inst.acc_wires[0][9] ),
    .B2(_11258_),
    .X(_01939_));
 sky130_fd_sc_hd__nand2_2 _23754_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[0][10] ),
    .Y(_10361_));
 sky130_fd_sc_hd__or2_2 _23755_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[10] ),
    .B(\systolic_inst.acc_wires[0][10] ),
    .X(_10362_));
 sky130_fd_sc_hd__and2_2 _23756_ (.A(_10361_),
    .B(_10362_),
    .X(_10363_));
 sky130_fd_sc_hd__a21oi_2 _23757_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[9] ),
    .A2(\systolic_inst.acc_wires[0][9] ),
    .B1(_10359_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand2_2 _23758_ (.A(_10358_),
    .B(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__xor2_2 _23759_ (.A(_10363_),
    .B(_10365_),
    .X(_10366_));
 sky130_fd_sc_hd__a22o_2 _23760_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][10] ),
    .B1(_11712_),
    .B2(_10366_),
    .X(_01940_));
 sky130_fd_sc_hd__nor2_2 _23761_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[0][11] ),
    .Y(_10367_));
 sky130_fd_sc_hd__or2_2 _23762_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[0][11] ),
    .X(_10368_));
 sky130_fd_sc_hd__nand2_2 _23763_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[11] ),
    .B(\systolic_inst.acc_wires[0][11] ),
    .Y(_10369_));
 sky130_fd_sc_hd__nand2_2 _23764_ (.A(_10368_),
    .B(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__a21bo_2 _23765_ (.A1(_10363_),
    .A2(_10365_),
    .B1_N(_10361_),
    .X(_10371_));
 sky130_fd_sc_hd__xnor2_2 _23766_ (.A(_10370_),
    .B(_10371_),
    .Y(_10372_));
 sky130_fd_sc_hd__a22o_2 _23767_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][11] ),
    .B1(_11712_),
    .B2(_10372_),
    .X(_01941_));
 sky130_fd_sc_hd__nand3_2 _23768_ (.A(_10363_),
    .B(_10368_),
    .C(_10369_),
    .Y(_10373_));
 sky130_fd_sc_hd__nor2_2 _23769_ (.A(_10357_),
    .B(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__o2bb2a_2 _23770_ (.A1_N(_10351_),
    .A2_N(_10374_),
    .B1(_10364_),
    .B2(_10373_),
    .X(_10375_));
 sky130_fd_sc_hd__o21a_2 _23771_ (.A1(_10361_),
    .A2(_10367_),
    .B1(_10369_),
    .X(_10376_));
 sky130_fd_sc_hd__xnor2_2 _23772_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[0][12] ),
    .Y(_10377_));
 sky130_fd_sc_hd__and3_2 _23773_ (.A(_10375_),
    .B(_10376_),
    .C(_10377_),
    .X(_10378_));
 sky130_fd_sc_hd__a21oi_2 _23774_ (.A1(_10375_),
    .A2(_10376_),
    .B1(_10377_),
    .Y(_10379_));
 sky130_fd_sc_hd__nor2_2 _23775_ (.A(_10378_),
    .B(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__a22o_2 _23776_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][12] ),
    .B1(_11712_),
    .B2(_10380_),
    .X(_01942_));
 sky130_fd_sc_hd__xor2_2 _23777_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[13] ),
    .B(\systolic_inst.acc_wires[0][13] ),
    .X(_10381_));
 sky130_fd_sc_hd__a211o_2 _23778_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[12] ),
    .A2(\systolic_inst.acc_wires[0][12] ),
    .B1(_10379_),
    .C1(_10381_),
    .X(_10382_));
 sky130_fd_sc_hd__nand2b_2 _23779_ (.A_N(_10377_),
    .B(_10381_),
    .Y(_10383_));
 sky130_fd_sc_hd__a21o_2 _23780_ (.A1(_10375_),
    .A2(_10376_),
    .B1(_10383_),
    .X(_10384_));
 sky130_fd_sc_hd__and3_2 _23781_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[12] ),
    .B(\systolic_inst.acc_wires[0][12] ),
    .C(_10381_),
    .X(_10385_));
 sky130_fd_sc_hd__nor2_2 _23782_ (.A(_11713_),
    .B(_10385_),
    .Y(_10386_));
 sky130_fd_sc_hd__a32o_2 _23783_ (.A1(_10382_),
    .A2(_10384_),
    .A3(_10386_),
    .B1(\systolic_inst.acc_wires[0][13] ),
    .B2(_11258_),
    .X(_01943_));
 sky130_fd_sc_hd__or2_2 _23784_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[0][14] ),
    .X(_10387_));
 sky130_fd_sc_hd__nand2_2 _23785_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[14] ),
    .B(\systolic_inst.acc_wires[0][14] ),
    .Y(_10388_));
 sky130_fd_sc_hd__and2_2 _23786_ (.A(_10387_),
    .B(_10388_),
    .X(_10389_));
 sky130_fd_sc_hd__a21oi_2 _23787_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[13] ),
    .A2(\systolic_inst.acc_wires[0][13] ),
    .B1(_10385_),
    .Y(_10390_));
 sky130_fd_sc_hd__nand2_2 _23788_ (.A(_10384_),
    .B(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__or2_2 _23789_ (.A(_10389_),
    .B(_10391_),
    .X(_10392_));
 sky130_fd_sc_hd__nand2_2 _23790_ (.A(_10389_),
    .B(_10391_),
    .Y(_10393_));
 sky130_fd_sc_hd__a32o_2 _23791_ (.A1(_11712_),
    .A2(_10392_),
    .A3(_10393_),
    .B1(\systolic_inst.acc_wires[0][14] ),
    .B2(_11258_),
    .X(_01944_));
 sky130_fd_sc_hd__nor2_2 _23792_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][15] ),
    .Y(_10394_));
 sky130_fd_sc_hd__and2_2 _23793_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][15] ),
    .X(_10395_));
 sky130_fd_sc_hd__o211ai_2 _23794_ (.A1(_10394_),
    .A2(_10395_),
    .B1(_10388_),
    .C1(_10393_),
    .Y(_10396_));
 sky130_fd_sc_hd__a211o_2 _23795_ (.A1(_10388_),
    .A2(_10393_),
    .B1(_10394_),
    .C1(_10395_),
    .X(_10397_));
 sky130_fd_sc_hd__a32o_2 _23796_ (.A1(_11712_),
    .A2(_10396_),
    .A3(_10397_),
    .B1(\systolic_inst.acc_wires[0][15] ),
    .B2(_11258_),
    .X(_01945_));
 sky130_fd_sc_hd__or3b_2 _23797_ (.A(_10394_),
    .B(_10395_),
    .C_N(_10389_),
    .X(_10398_));
 sky130_fd_sc_hd__a21o_2 _23798_ (.A1(_10384_),
    .A2(_10390_),
    .B1(_10398_),
    .X(_10399_));
 sky130_fd_sc_hd__o21ba_2 _23799_ (.A1(_10388_),
    .A2(_10394_),
    .B1_N(_10395_),
    .X(_10400_));
 sky130_fd_sc_hd__and2_2 _23800_ (.A(_10399_),
    .B(_10400_),
    .X(_10401_));
 sky130_fd_sc_hd__xnor2_2 _23801_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][16] ),
    .Y(_10402_));
 sky130_fd_sc_hd__nand2_2 _23802_ (.A(_10401_),
    .B(_10402_),
    .Y(_10403_));
 sky130_fd_sc_hd__nor2_2 _23803_ (.A(_10401_),
    .B(_10402_),
    .Y(_10404_));
 sky130_fd_sc_hd__nor2_2 _23804_ (.A(_11713_),
    .B(_10404_),
    .Y(_10405_));
 sky130_fd_sc_hd__a22o_2 _23805_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][16] ),
    .B1(_10403_),
    .B2(_10405_),
    .X(_01946_));
 sky130_fd_sc_hd__xor2_2 _23806_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][17] ),
    .X(_10406_));
 sky130_fd_sc_hd__inv_2 _23807_ (.A(_10406_),
    .Y(_10407_));
 sky130_fd_sc_hd__a21oi_2 _23808_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[0][16] ),
    .B1(_10404_),
    .Y(_10408_));
 sky130_fd_sc_hd__xnor2_2 _23809_ (.A(_10406_),
    .B(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__a22o_2 _23810_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][17] ),
    .B1(_11712_),
    .B2(_10409_),
    .X(_01947_));
 sky130_fd_sc_hd__or2_2 _23811_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][18] ),
    .X(_10410_));
 sky130_fd_sc_hd__nand2_2 _23812_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][18] ),
    .Y(_10411_));
 sky130_fd_sc_hd__nand2_2 _23813_ (.A(_10410_),
    .B(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__o21a_2 _23814_ (.A1(\systolic_inst.acc_wires[0][16] ),
    .A2(\systolic_inst.acc_wires[0][17] ),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .X(_10413_));
 sky130_fd_sc_hd__a21oi_2 _23815_ (.A1(_10404_),
    .A2(_10406_),
    .B1(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__xor2_2 _23816_ (.A(_10412_),
    .B(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__a22o_2 _23817_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][18] ),
    .B1(_11712_),
    .B2(_10415_),
    .X(_01948_));
 sky130_fd_sc_hd__xnor2_2 _23818_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][19] ),
    .Y(_10416_));
 sky130_fd_sc_hd__o21ai_2 _23819_ (.A1(_10412_),
    .A2(_10414_),
    .B1(_10411_),
    .Y(_10417_));
 sky130_fd_sc_hd__xnor2_2 _23820_ (.A(_10416_),
    .B(_10417_),
    .Y(_10418_));
 sky130_fd_sc_hd__a22o_2 _23821_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][19] ),
    .B1(_11712_),
    .B2(_10418_),
    .X(_01949_));
 sky130_fd_sc_hd__xor2_2 _23822_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][20] ),
    .X(_10419_));
 sky130_fd_sc_hd__or4_2 _23823_ (.A(_10402_),
    .B(_10407_),
    .C(_10412_),
    .D(_10416_),
    .X(_10420_));
 sky130_fd_sc_hd__nor2_2 _23824_ (.A(_10401_),
    .B(_10420_),
    .Y(_10421_));
 sky130_fd_sc_hd__o41a_2 _23825_ (.A1(\systolic_inst.acc_wires[0][16] ),
    .A2(\systolic_inst.acc_wires[0][17] ),
    .A3(\systolic_inst.acc_wires[0][18] ),
    .A4(\systolic_inst.acc_wires[0][19] ),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .X(_10422_));
 sky130_fd_sc_hd__or3_2 _23826_ (.A(_10419_),
    .B(_10421_),
    .C(_10422_),
    .X(_10423_));
 sky130_fd_sc_hd__o21ai_2 _23827_ (.A1(_10421_),
    .A2(_10422_),
    .B1(_10419_),
    .Y(_10424_));
 sky130_fd_sc_hd__a32o_2 _23828_ (.A1(_11712_),
    .A2(_10423_),
    .A3(_10424_),
    .B1(\systolic_inst.acc_wires[0][20] ),
    .B2(_11258_),
    .X(_01950_));
 sky130_fd_sc_hd__xor2_2 _23829_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][21] ),
    .X(_10425_));
 sky130_fd_sc_hd__a21bo_2 _23830_ (.A1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .A2(\systolic_inst.acc_wires[0][20] ),
    .B1_N(_10424_),
    .X(_10426_));
 sky130_fd_sc_hd__xor2_2 _23831_ (.A(_10425_),
    .B(_10426_),
    .X(_10427_));
 sky130_fd_sc_hd__a22o_2 _23832_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][21] ),
    .B1(_11712_),
    .B2(_10427_),
    .X(_01951_));
 sky130_fd_sc_hd__or2_2 _23833_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][22] ),
    .X(_10428_));
 sky130_fd_sc_hd__nand2_2 _23834_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][22] ),
    .Y(_10429_));
 sky130_fd_sc_hd__and2_2 _23835_ (.A(_10428_),
    .B(_10429_),
    .X(_10430_));
 sky130_fd_sc_hd__o21a_2 _23836_ (.A1(\systolic_inst.acc_wires[0][20] ),
    .A2(\systolic_inst.acc_wires[0][21] ),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .X(_10431_));
 sky130_fd_sc_hd__and2b_2 _23837_ (.A_N(_10424_),
    .B(_10425_),
    .X(_10432_));
 sky130_fd_sc_hd__o21ai_2 _23838_ (.A1(_10431_),
    .A2(_10432_),
    .B1(_10430_),
    .Y(_10433_));
 sky130_fd_sc_hd__or3_2 _23839_ (.A(_10430_),
    .B(_10431_),
    .C(_10432_),
    .X(_10434_));
 sky130_fd_sc_hd__a32o_2 _23840_ (.A1(_11712_),
    .A2(_10433_),
    .A3(_10434_),
    .B1(\systolic_inst.acc_wires[0][22] ),
    .B2(_11258_),
    .X(_01952_));
 sky130_fd_sc_hd__xnor2_2 _23841_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][23] ),
    .Y(_10435_));
 sky130_fd_sc_hd__inv_2 _23842_ (.A(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__a21oi_2 _23843_ (.A1(_10429_),
    .A2(_10433_),
    .B1(_10435_),
    .Y(_10437_));
 sky130_fd_sc_hd__a31o_2 _23844_ (.A1(_10429_),
    .A2(_10433_),
    .A3(_10435_),
    .B1(_11713_),
    .X(_10438_));
 sky130_fd_sc_hd__a2bb2o_2 _23845_ (.A1_N(_10438_),
    .A2_N(_10437_),
    .B1(\systolic_inst.acc_wires[0][23] ),
    .B2(_11258_),
    .X(_01953_));
 sky130_fd_sc_hd__nand4_2 _23846_ (.A(_10419_),
    .B(_10425_),
    .C(_10430_),
    .D(_10436_),
    .Y(_10439_));
 sky130_fd_sc_hd__a211o_2 _23847_ (.A1(_10399_),
    .A2(_10400_),
    .B1(_10420_),
    .C1(_10439_),
    .X(_10440_));
 sky130_fd_sc_hd__o41a_2 _23848_ (.A1(\systolic_inst.acc_wires[0][20] ),
    .A2(\systolic_inst.acc_wires[0][21] ),
    .A3(\systolic_inst.acc_wires[0][22] ),
    .A4(\systolic_inst.acc_wires[0][23] ),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .X(_10441_));
 sky130_fd_sc_hd__nor2_2 _23849_ (.A(_10422_),
    .B(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__nor2_2 _23850_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][24] ),
    .Y(_10443_));
 sky130_fd_sc_hd__and2_2 _23851_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][24] ),
    .X(_10444_));
 sky130_fd_sc_hd__or2_2 _23852_ (.A(_10443_),
    .B(_10444_),
    .X(_10445_));
 sky130_fd_sc_hd__a21oi_2 _23853_ (.A1(_10440_),
    .A2(_10442_),
    .B1(_10445_),
    .Y(_10446_));
 sky130_fd_sc_hd__a31o_2 _23854_ (.A1(_10440_),
    .A2(_10442_),
    .A3(_10445_),
    .B1(_11713_),
    .X(_10447_));
 sky130_fd_sc_hd__a2bb2o_2 _23855_ (.A1_N(_10447_),
    .A2_N(_10446_),
    .B1(\systolic_inst.acc_wires[0][24] ),
    .B2(_11258_),
    .X(_01954_));
 sky130_fd_sc_hd__xor2_2 _23856_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][25] ),
    .X(_10448_));
 sky130_fd_sc_hd__or3_2 _23857_ (.A(_10444_),
    .B(_10446_),
    .C(_10448_),
    .X(_10449_));
 sky130_fd_sc_hd__o21ai_2 _23858_ (.A1(_10444_),
    .A2(_10446_),
    .B1(_10448_),
    .Y(_10450_));
 sky130_fd_sc_hd__a32o_2 _23859_ (.A1(_11712_),
    .A2(_10449_),
    .A3(_10450_),
    .B1(\systolic_inst.acc_wires[0][25] ),
    .B2(_11258_),
    .X(_01955_));
 sky130_fd_sc_hd__or2_2 _23860_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][26] ),
    .X(_10451_));
 sky130_fd_sc_hd__nand2_2 _23861_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][26] ),
    .Y(_10452_));
 sky130_fd_sc_hd__nand2_2 _23862_ (.A(_10451_),
    .B(_10452_),
    .Y(_10453_));
 sky130_fd_sc_hd__o21a_2 _23863_ (.A1(\systolic_inst.acc_wires[0][24] ),
    .A2(\systolic_inst.acc_wires[0][25] ),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .X(_10454_));
 sky130_fd_sc_hd__a21o_2 _23864_ (.A1(_10446_),
    .A2(_10448_),
    .B1(_10454_),
    .X(_10455_));
 sky130_fd_sc_hd__xnor2_2 _23865_ (.A(_10453_),
    .B(_10455_),
    .Y(_10456_));
 sky130_fd_sc_hd__a22o_2 _23866_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][26] ),
    .B1(_11712_),
    .B2(_10456_),
    .X(_01956_));
 sky130_fd_sc_hd__xnor2_2 _23867_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][27] ),
    .Y(_10457_));
 sky130_fd_sc_hd__a21bo_2 _23868_ (.A1(_10451_),
    .A2(_10455_),
    .B1_N(_10452_),
    .X(_10458_));
 sky130_fd_sc_hd__xnor2_2 _23869_ (.A(_10457_),
    .B(_10458_),
    .Y(_10459_));
 sky130_fd_sc_hd__a22o_2 _23870_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][27] ),
    .B1(_11712_),
    .B2(_10459_),
    .X(_01957_));
 sky130_fd_sc_hd__nor2_2 _23871_ (.A(_10453_),
    .B(_10457_),
    .Y(_10460_));
 sky130_fd_sc_hd__o21a_2 _23872_ (.A1(\systolic_inst.acc_wires[0][26] ),
    .A2(\systolic_inst.acc_wires[0][27] ),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .X(_10461_));
 sky130_fd_sc_hd__a311oi_2 _23873_ (.A1(_10446_),
    .A2(_10448_),
    .A3(_10460_),
    .B1(_10461_),
    .C1(_10454_),
    .Y(_10462_));
 sky130_fd_sc_hd__or2_2 _23874_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][28] ),
    .X(_10463_));
 sky130_fd_sc_hd__nand2_2 _23875_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][28] ),
    .Y(_10464_));
 sky130_fd_sc_hd__nand2_2 _23876_ (.A(_10463_),
    .B(_10464_),
    .Y(_10465_));
 sky130_fd_sc_hd__xor2_2 _23877_ (.A(_10462_),
    .B(_10465_),
    .X(_10466_));
 sky130_fd_sc_hd__a22o_2 _23878_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][28] ),
    .B1(_11712_),
    .B2(_10466_),
    .X(_01958_));
 sky130_fd_sc_hd__xor2_2 _23879_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][29] ),
    .X(_10467_));
 sky130_fd_sc_hd__inv_2 _23880_ (.A(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__o21a_2 _23881_ (.A1(_10462_),
    .A2(_10465_),
    .B1(_10464_),
    .X(_10469_));
 sky130_fd_sc_hd__xnor2_2 _23882_ (.A(_10467_),
    .B(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__a22o_2 _23883_ (.A1(_11258_),
    .A2(\systolic_inst.acc_wires[0][29] ),
    .B1(_11712_),
    .B2(_10470_),
    .X(_01959_));
 sky130_fd_sc_hd__o21ai_2 _23884_ (.A1(\systolic_inst.acc_wires[0][28] ),
    .A2(\systolic_inst.acc_wires[0][29] ),
    .B1(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .Y(_10471_));
 sky130_fd_sc_hd__o31a_2 _23885_ (.A1(_10462_),
    .A2(_10465_),
    .A3(_10468_),
    .B1(_10471_),
    .X(_10472_));
 sky130_fd_sc_hd__nand2_2 _23886_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][30] ),
    .Y(_10473_));
 sky130_fd_sc_hd__or2_2 _23887_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][30] ),
    .X(_10474_));
 sky130_fd_sc_hd__nand2_2 _23888_ (.A(_10473_),
    .B(_10474_),
    .Y(_10475_));
 sky130_fd_sc_hd__nand2_2 _23889_ (.A(_10472_),
    .B(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__or2_2 _23890_ (.A(_10472_),
    .B(_10475_),
    .X(_10477_));
 sky130_fd_sc_hd__a32o_2 _23891_ (.A1(_11712_),
    .A2(_10476_),
    .A3(_10477_),
    .B1(\systolic_inst.acc_wires[0][30] ),
    .B2(_11258_),
    .X(_01960_));
 sky130_fd_sc_hd__xnor2_2 _23892_ (.A(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ),
    .B(\systolic_inst.acc_wires[0][31] ),
    .Y(_10478_));
 sky130_fd_sc_hd__a21oi_2 _23893_ (.A1(_10473_),
    .A2(_10477_),
    .B1(_10478_),
    .Y(_10479_));
 sky130_fd_sc_hd__a31o_2 _23894_ (.A1(_10473_),
    .A2(_10477_),
    .A3(_10478_),
    .B1(_11713_),
    .X(_10480_));
 sky130_fd_sc_hd__a2bb2o_2 _23895_ (.A1_N(_10480_),
    .A2_N(_10479_),
    .B1(\systolic_inst.acc_wires[0][31] ),
    .B2(_11258_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _23896_ (.A0(\systolic_inst.B_shift[17][0] ),
    .A1(\B_in[72] ),
    .S(_00008_),
    .X(_10481_));
 sky130_fd_sc_hd__mux2_1 _23897_ (.A0(_10481_),
    .A1(\systolic_inst.B_shift[13][0] ),
    .S(_11332_),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _23898_ (.A0(\systolic_inst.B_shift[17][1] ),
    .A1(\B_in[73] ),
    .S(_00008_),
    .X(_10482_));
 sky130_fd_sc_hd__mux2_1 _23899_ (.A0(_10482_),
    .A1(\systolic_inst.B_shift[13][1] ),
    .S(_11332_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _23900_ (.A0(\systolic_inst.B_shift[17][2] ),
    .A1(\B_in[74] ),
    .S(_00008_),
    .X(_10483_));
 sky130_fd_sc_hd__mux2_1 _23901_ (.A0(_10483_),
    .A1(\systolic_inst.B_shift[13][2] ),
    .S(_11332_),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _23902_ (.A0(\systolic_inst.B_shift[17][3] ),
    .A1(\B_in[75] ),
    .S(_00008_),
    .X(_10484_));
 sky130_fd_sc_hd__mux2_1 _23903_ (.A0(_10484_),
    .A1(\systolic_inst.B_shift[13][3] ),
    .S(_11332_),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _23904_ (.A0(\systolic_inst.B_shift[17][4] ),
    .A1(\B_in[76] ),
    .S(_00008_),
    .X(_10485_));
 sky130_fd_sc_hd__mux2_1 _23905_ (.A0(_10485_),
    .A1(\systolic_inst.B_shift[13][4] ),
    .S(_11332_),
    .X(_01966_));
 sky130_fd_sc_hd__mux2_1 _23906_ (.A0(\systolic_inst.B_shift[17][5] ),
    .A1(\B_in[77] ),
    .S(_00008_),
    .X(_10486_));
 sky130_fd_sc_hd__mux2_1 _23907_ (.A0(_10486_),
    .A1(\systolic_inst.B_shift[13][5] ),
    .S(_11332_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _23908_ (.A0(\systolic_inst.B_shift[17][6] ),
    .A1(\B_in[78] ),
    .S(_00008_),
    .X(_10487_));
 sky130_fd_sc_hd__mux2_1 _23909_ (.A0(_10487_),
    .A1(\systolic_inst.B_shift[13][6] ),
    .S(_11332_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _23910_ (.A0(\systolic_inst.B_shift[17][7] ),
    .A1(\B_in[79] ),
    .S(_00008_),
    .X(_10488_));
 sky130_fd_sc_hd__mux2_1 _23911_ (.A0(_10488_),
    .A1(\systolic_inst.B_shift[13][7] ),
    .S(_11332_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _23912_ (.A0(\systolic_inst.B_shift[22][0] ),
    .A1(\B_in[80] ),
    .S(_00008_),
    .X(_10489_));
 sky130_fd_sc_hd__mux2_1 _23913_ (.A0(_10489_),
    .A1(\systolic_inst.B_shift[18][0] ),
    .S(_11332_),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _23914_ (.A0(\systolic_inst.B_shift[22][1] ),
    .A1(\B_in[81] ),
    .S(_00008_),
    .X(_10490_));
 sky130_fd_sc_hd__mux2_1 _23915_ (.A0(_10490_),
    .A1(\systolic_inst.B_shift[18][1] ),
    .S(_11332_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _23916_ (.A0(\systolic_inst.B_shift[22][2] ),
    .A1(\B_in[82] ),
    .S(_00008_),
    .X(_10491_));
 sky130_fd_sc_hd__mux2_1 _23917_ (.A0(_10491_),
    .A1(\systolic_inst.B_shift[18][2] ),
    .S(_11332_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _23918_ (.A0(\systolic_inst.B_shift[22][3] ),
    .A1(\B_in[83] ),
    .S(_00008_),
    .X(_10492_));
 sky130_fd_sc_hd__mux2_1 _23919_ (.A0(_10492_),
    .A1(\systolic_inst.B_shift[18][3] ),
    .S(_11332_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _23920_ (.A0(\systolic_inst.B_shift[22][4] ),
    .A1(\B_in[84] ),
    .S(_00008_),
    .X(_10493_));
 sky130_fd_sc_hd__mux2_1 _23921_ (.A0(_10493_),
    .A1(\systolic_inst.B_shift[18][4] ),
    .S(_11332_),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_1 _23922_ (.A0(\systolic_inst.B_shift[22][5] ),
    .A1(\B_in[85] ),
    .S(_00008_),
    .X(_10494_));
 sky130_fd_sc_hd__mux2_1 _23923_ (.A0(_10494_),
    .A1(\systolic_inst.B_shift[18][5] ),
    .S(_11332_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _23924_ (.A0(\systolic_inst.B_shift[22][6] ),
    .A1(\B_in[86] ),
    .S(_00008_),
    .X(_10495_));
 sky130_fd_sc_hd__mux2_1 _23925_ (.A0(_10495_),
    .A1(\systolic_inst.B_shift[18][6] ),
    .S(_11332_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _23926_ (.A0(\systolic_inst.B_shift[22][7] ),
    .A1(\B_in[87] ),
    .S(_00008_),
    .X(_10496_));
 sky130_fd_sc_hd__mux2_1 _23927_ (.A0(_10496_),
    .A1(\systolic_inst.B_shift[18][7] ),
    .S(_11332_),
    .X(_01977_));
 sky130_fd_sc_hd__a22o_2 _23928_ (.A1(\systolic_inst.A_shift[3][0] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[24] ),
    .X(_01978_));
 sky130_fd_sc_hd__a22o_2 _23929_ (.A1(\systolic_inst.A_shift[3][1] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[25] ),
    .X(_01979_));
 sky130_fd_sc_hd__a22o_2 _23930_ (.A1(\systolic_inst.A_shift[3][2] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[26] ),
    .X(_01980_));
 sky130_fd_sc_hd__a22o_2 _23931_ (.A1(\systolic_inst.A_shift[3][3] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[27] ),
    .X(_01981_));
 sky130_fd_sc_hd__a22o_2 _23932_ (.A1(\systolic_inst.A_shift[3][4] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[28] ),
    .X(_01982_));
 sky130_fd_sc_hd__a22o_2 _23933_ (.A1(\systolic_inst.A_shift[3][5] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[29] ),
    .X(_01983_));
 sky130_fd_sc_hd__a22o_2 _23934_ (.A1(\systolic_inst.A_shift[3][6] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[30] ),
    .X(_01984_));
 sky130_fd_sc_hd__a22o_2 _23935_ (.A1(\systolic_inst.A_shift[3][7] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[31] ),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _23936_ (.A0(\systolic_inst.B_shift[14][0] ),
    .A1(\B_in[16] ),
    .S(_00008_),
    .X(_10497_));
 sky130_fd_sc_hd__mux2_1 _23937_ (.A0(_10497_),
    .A1(\systolic_inst.B_shift[10][0] ),
    .S(_11332_),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_1 _23938_ (.A0(\systolic_inst.B_shift[14][1] ),
    .A1(\B_in[17] ),
    .S(_00008_),
    .X(_10498_));
 sky130_fd_sc_hd__mux2_1 _23939_ (.A0(_10498_),
    .A1(\systolic_inst.B_shift[10][1] ),
    .S(_11332_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _23940_ (.A0(\systolic_inst.B_shift[14][2] ),
    .A1(\B_in[18] ),
    .S(_00008_),
    .X(_10499_));
 sky130_fd_sc_hd__mux2_1 _23941_ (.A0(_10499_),
    .A1(\systolic_inst.B_shift[10][2] ),
    .S(_11332_),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _23942_ (.A0(\systolic_inst.B_shift[14][3] ),
    .A1(\B_in[19] ),
    .S(_00008_),
    .X(_10500_));
 sky130_fd_sc_hd__mux2_1 _23943_ (.A0(_10500_),
    .A1(\systolic_inst.B_shift[10][3] ),
    .S(_11332_),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_1 _23944_ (.A0(\systolic_inst.B_shift[14][4] ),
    .A1(\B_in[20] ),
    .S(_00008_),
    .X(_10501_));
 sky130_fd_sc_hd__mux2_1 _23945_ (.A0(_10501_),
    .A1(\systolic_inst.B_shift[10][4] ),
    .S(_11332_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _23946_ (.A0(\systolic_inst.B_shift[14][5] ),
    .A1(\B_in[21] ),
    .S(_00008_),
    .X(_10502_));
 sky130_fd_sc_hd__mux2_1 _23947_ (.A0(_10502_),
    .A1(\systolic_inst.B_shift[10][5] ),
    .S(_11332_),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _23948_ (.A0(\systolic_inst.B_shift[14][6] ),
    .A1(\B_in[22] ),
    .S(_00008_),
    .X(_10503_));
 sky130_fd_sc_hd__mux2_1 _23949_ (.A0(_10503_),
    .A1(\systolic_inst.B_shift[10][6] ),
    .S(_11332_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_1 _23950_ (.A0(\systolic_inst.B_shift[14][7] ),
    .A1(\B_in[23] ),
    .S(_00008_),
    .X(_10504_));
 sky130_fd_sc_hd__mux2_1 _23951_ (.A0(_10504_),
    .A1(\systolic_inst.B_shift[10][7] ),
    .S(_11332_),
    .X(_01993_));
 sky130_fd_sc_hd__and2_2 _23952_ (.A(\systolic_inst.ce_local ),
    .B(rst_n),
    .X(_10505_));
 sky130_fd_sc_hd__a22o_2 _23953_ (.A1(\systolic_inst.B_shift[11][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[15][0] ),
    .X(_01994_));
 sky130_fd_sc_hd__a22o_2 _23954_ (.A1(\systolic_inst.B_shift[11][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[15][1] ),
    .X(_01995_));
 sky130_fd_sc_hd__a22o_2 _23955_ (.A1(\systolic_inst.B_shift[11][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[15][2] ),
    .X(_01996_));
 sky130_fd_sc_hd__a22o_2 _23956_ (.A1(\systolic_inst.B_shift[11][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[15][3] ),
    .X(_01997_));
 sky130_fd_sc_hd__a22o_2 _23957_ (.A1(\systolic_inst.B_shift[11][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[15][4] ),
    .X(_01998_));
 sky130_fd_sc_hd__a22o_2 _23958_ (.A1(\systolic_inst.B_shift[11][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[15][5] ),
    .X(_01999_));
 sky130_fd_sc_hd__a22o_2 _23959_ (.A1(\systolic_inst.B_shift[11][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[15][6] ),
    .X(_02000_));
 sky130_fd_sc_hd__a22o_2 _23960_ (.A1(\systolic_inst.B_shift[11][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[15][7] ),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_1 _23961_ (.A0(\systolic_inst.B_shift[13][0] ),
    .A1(\B_in[40] ),
    .S(_00008_),
    .X(_10506_));
 sky130_fd_sc_hd__mux2_1 _23962_ (.A0(_10506_),
    .A1(\systolic_inst.B_shift[9][0] ),
    .S(_11332_),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_1 _23963_ (.A0(\systolic_inst.B_shift[13][1] ),
    .A1(\B_in[41] ),
    .S(_00008_),
    .X(_10507_));
 sky130_fd_sc_hd__mux2_1 _23964_ (.A0(_10507_),
    .A1(\systolic_inst.B_shift[9][1] ),
    .S(_11332_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _23965_ (.A0(\systolic_inst.B_shift[13][2] ),
    .A1(\B_in[42] ),
    .S(_00008_),
    .X(_10508_));
 sky130_fd_sc_hd__mux2_1 _23966_ (.A0(_10508_),
    .A1(\systolic_inst.B_shift[9][2] ),
    .S(_11332_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _23967_ (.A0(\systolic_inst.B_shift[13][3] ),
    .A1(\B_in[43] ),
    .S(_00008_),
    .X(_10509_));
 sky130_fd_sc_hd__mux2_1 _23968_ (.A0(_10509_),
    .A1(\systolic_inst.B_shift[9][3] ),
    .S(_11332_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _23969_ (.A0(\systolic_inst.B_shift[13][4] ),
    .A1(\B_in[44] ),
    .S(_00008_),
    .X(_10510_));
 sky130_fd_sc_hd__mux2_1 _23970_ (.A0(_10510_),
    .A1(\systolic_inst.B_shift[9][4] ),
    .S(_11332_),
    .X(_02006_));
 sky130_fd_sc_hd__mux2_1 _23971_ (.A0(\systolic_inst.B_shift[13][5] ),
    .A1(\B_in[45] ),
    .S(_00008_),
    .X(_10511_));
 sky130_fd_sc_hd__mux2_1 _23972_ (.A0(_10511_),
    .A1(\systolic_inst.B_shift[9][5] ),
    .S(_11332_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_1 _23973_ (.A0(\systolic_inst.B_shift[13][6] ),
    .A1(\B_in[46] ),
    .S(_00008_),
    .X(_10512_));
 sky130_fd_sc_hd__mux2_1 _23974_ (.A0(_10512_),
    .A1(\systolic_inst.B_shift[9][6] ),
    .S(_11332_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _23975_ (.A0(\systolic_inst.B_shift[13][7] ),
    .A1(\B_in[47] ),
    .S(_00008_),
    .X(_10513_));
 sky130_fd_sc_hd__mux2_1 _23976_ (.A0(_10513_),
    .A1(\systolic_inst.B_shift[9][7] ),
    .S(_11332_),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _23977_ (.A0(\systolic_inst.B_shift[12][0] ),
    .A1(\B_in[64] ),
    .S(_00008_),
    .X(_10514_));
 sky130_fd_sc_hd__mux2_1 _23978_ (.A0(_10514_),
    .A1(\systolic_inst.B_shift[8][0] ),
    .S(_11332_),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_1 _23979_ (.A0(\systolic_inst.B_shift[12][1] ),
    .A1(\B_in[65] ),
    .S(_00008_),
    .X(_10515_));
 sky130_fd_sc_hd__mux2_1 _23980_ (.A0(_10515_),
    .A1(\systolic_inst.B_shift[8][1] ),
    .S(_11332_),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_1 _23981_ (.A0(\systolic_inst.B_shift[12][2] ),
    .A1(\B_in[66] ),
    .S(_00008_),
    .X(_10516_));
 sky130_fd_sc_hd__mux2_1 _23982_ (.A0(_10516_),
    .A1(\systolic_inst.B_shift[8][2] ),
    .S(_11332_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _23983_ (.A0(\systolic_inst.B_shift[12][3] ),
    .A1(\B_in[67] ),
    .S(_00008_),
    .X(_10517_));
 sky130_fd_sc_hd__mux2_1 _23984_ (.A0(_10517_),
    .A1(\systolic_inst.B_shift[8][3] ),
    .S(_11332_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _23985_ (.A0(\systolic_inst.B_shift[12][4] ),
    .A1(\B_in[68] ),
    .S(_00008_),
    .X(_10518_));
 sky130_fd_sc_hd__mux2_1 _23986_ (.A0(_10518_),
    .A1(\systolic_inst.B_shift[8][4] ),
    .S(_11332_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _23987_ (.A0(\systolic_inst.B_shift[12][5] ),
    .A1(\B_in[69] ),
    .S(_00008_),
    .X(_10519_));
 sky130_fd_sc_hd__mux2_1 _23988_ (.A0(_10519_),
    .A1(\systolic_inst.B_shift[8][5] ),
    .S(_11332_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _23989_ (.A0(\systolic_inst.B_shift[12][6] ),
    .A1(\B_in[70] ),
    .S(_00008_),
    .X(_10520_));
 sky130_fd_sc_hd__mux2_1 _23990_ (.A0(_10520_),
    .A1(\systolic_inst.B_shift[8][6] ),
    .S(_11332_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _23991_ (.A0(\systolic_inst.B_shift[12][7] ),
    .A1(\B_in[71] ),
    .S(_00008_),
    .X(_10521_));
 sky130_fd_sc_hd__mux2_1 _23992_ (.A0(_10521_),
    .A1(\systolic_inst.B_shift[8][7] ),
    .S(_11332_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _23993_ (.A0(\systolic_inst.B_shift[9][0] ),
    .A1(\B_in[8] ),
    .S(_00008_),
    .X(_10522_));
 sky130_fd_sc_hd__mux2_1 _23994_ (.A0(_10522_),
    .A1(\systolic_inst.B_shift[5][0] ),
    .S(_11332_),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _23995_ (.A0(\systolic_inst.B_shift[9][1] ),
    .A1(\B_in[9] ),
    .S(_00008_),
    .X(_10523_));
 sky130_fd_sc_hd__mux2_1 _23996_ (.A0(_10523_),
    .A1(\systolic_inst.B_shift[5][1] ),
    .S(_11332_),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _23997_ (.A0(\systolic_inst.B_shift[9][2] ),
    .A1(\B_in[10] ),
    .S(_00008_),
    .X(_10524_));
 sky130_fd_sc_hd__mux2_1 _23998_ (.A0(_10524_),
    .A1(\systolic_inst.B_shift[5][2] ),
    .S(_11332_),
    .X(_02020_));
 sky130_fd_sc_hd__mux2_1 _23999_ (.A0(\systolic_inst.B_shift[9][3] ),
    .A1(\B_in[11] ),
    .S(_00008_),
    .X(_10525_));
 sky130_fd_sc_hd__mux2_1 _24000_ (.A0(_10525_),
    .A1(\systolic_inst.B_shift[5][3] ),
    .S(_11332_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _24001_ (.A0(\systolic_inst.B_shift[9][4] ),
    .A1(\B_in[12] ),
    .S(_00008_),
    .X(_10526_));
 sky130_fd_sc_hd__mux2_1 _24002_ (.A0(_10526_),
    .A1(\systolic_inst.B_shift[5][4] ),
    .S(_11332_),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_1 _24003_ (.A0(\systolic_inst.B_shift[9][5] ),
    .A1(\B_in[13] ),
    .S(_00008_),
    .X(_10527_));
 sky130_fd_sc_hd__mux2_1 _24004_ (.A0(_10527_),
    .A1(\systolic_inst.B_shift[5][5] ),
    .S(_11332_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _24005_ (.A0(\systolic_inst.B_shift[9][6] ),
    .A1(\B_in[14] ),
    .S(_00008_),
    .X(_10528_));
 sky130_fd_sc_hd__mux2_1 _24006_ (.A0(_10528_),
    .A1(\systolic_inst.B_shift[5][6] ),
    .S(_11332_),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _24007_ (.A0(\systolic_inst.B_shift[9][7] ),
    .A1(\B_in[15] ),
    .S(_00008_),
    .X(_10529_));
 sky130_fd_sc_hd__mux2_1 _24008_ (.A0(_10529_),
    .A1(\systolic_inst.B_shift[5][7] ),
    .S(_11332_),
    .X(_02025_));
 sky130_fd_sc_hd__a22o_2 _24009_ (.A1(\systolic_inst.B_shift[7][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[11][0] ),
    .X(_02026_));
 sky130_fd_sc_hd__a22o_2 _24010_ (.A1(\systolic_inst.B_shift[7][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[11][1] ),
    .X(_02027_));
 sky130_fd_sc_hd__a22o_2 _24011_ (.A1(\systolic_inst.B_shift[7][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[11][2] ),
    .X(_02028_));
 sky130_fd_sc_hd__a22o_2 _24012_ (.A1(\systolic_inst.B_shift[7][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[11][3] ),
    .X(_02029_));
 sky130_fd_sc_hd__a22o_2 _24013_ (.A1(\systolic_inst.B_shift[7][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[11][4] ),
    .X(_02030_));
 sky130_fd_sc_hd__a22o_2 _24014_ (.A1(\systolic_inst.B_shift[7][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[11][5] ),
    .X(_02031_));
 sky130_fd_sc_hd__a22o_2 _24015_ (.A1(\systolic_inst.B_shift[7][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[11][6] ),
    .X(_02032_));
 sky130_fd_sc_hd__a22o_2 _24016_ (.A1(\systolic_inst.B_shift[7][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[11][7] ),
    .X(_02033_));
 sky130_fd_sc_hd__a22o_2 _24017_ (.A1(\systolic_inst.B_shift[6][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[10][0] ),
    .X(_02034_));
 sky130_fd_sc_hd__a22o_2 _24018_ (.A1(\systolic_inst.B_shift[6][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[10][1] ),
    .X(_02035_));
 sky130_fd_sc_hd__a22o_2 _24019_ (.A1(\systolic_inst.B_shift[6][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[10][2] ),
    .X(_02036_));
 sky130_fd_sc_hd__a22o_2 _24020_ (.A1(\systolic_inst.B_shift[6][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[10][3] ),
    .X(_02037_));
 sky130_fd_sc_hd__a22o_2 _24021_ (.A1(\systolic_inst.B_shift[6][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[10][4] ),
    .X(_02038_));
 sky130_fd_sc_hd__a22o_2 _24022_ (.A1(\systolic_inst.B_shift[6][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[10][5] ),
    .X(_02039_));
 sky130_fd_sc_hd__a22o_2 _24023_ (.A1(\systolic_inst.B_shift[6][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[10][6] ),
    .X(_02040_));
 sky130_fd_sc_hd__a22o_2 _24024_ (.A1(\systolic_inst.B_shift[6][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[10][7] ),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _24025_ (.A0(\systolic_inst.B_shift[8][0] ),
    .A1(\B_in[32] ),
    .S(_00008_),
    .X(_10530_));
 sky130_fd_sc_hd__mux2_1 _24026_ (.A0(_10530_),
    .A1(\systolic_inst.B_shift[4][0] ),
    .S(_11332_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _24027_ (.A0(\systolic_inst.B_shift[8][1] ),
    .A1(\B_in[33] ),
    .S(_00008_),
    .X(_10531_));
 sky130_fd_sc_hd__mux2_1 _24028_ (.A0(_10531_),
    .A1(\systolic_inst.B_shift[4][1] ),
    .S(_11332_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _24029_ (.A0(\systolic_inst.B_shift[8][2] ),
    .A1(\B_in[34] ),
    .S(_00008_),
    .X(_10532_));
 sky130_fd_sc_hd__mux2_1 _24030_ (.A0(_10532_),
    .A1(\systolic_inst.B_shift[4][2] ),
    .S(_11332_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _24031_ (.A0(\systolic_inst.B_shift[8][3] ),
    .A1(\B_in[35] ),
    .S(_00008_),
    .X(_10533_));
 sky130_fd_sc_hd__mux2_1 _24032_ (.A0(_10533_),
    .A1(\systolic_inst.B_shift[4][3] ),
    .S(_11332_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _24033_ (.A0(\systolic_inst.B_shift[8][4] ),
    .A1(\B_in[36] ),
    .S(_00008_),
    .X(_10534_));
 sky130_fd_sc_hd__mux2_1 _24034_ (.A0(_10534_),
    .A1(\systolic_inst.B_shift[4][4] ),
    .S(_11332_),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _24035_ (.A0(\systolic_inst.B_shift[8][5] ),
    .A1(\B_in[37] ),
    .S(_00008_),
    .X(_10535_));
 sky130_fd_sc_hd__mux2_1 _24036_ (.A0(_10535_),
    .A1(\systolic_inst.B_shift[4][5] ),
    .S(_11332_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _24037_ (.A0(\systolic_inst.B_shift[8][6] ),
    .A1(\B_in[38] ),
    .S(_00008_),
    .X(_10536_));
 sky130_fd_sc_hd__mux2_1 _24038_ (.A0(_10536_),
    .A1(\systolic_inst.B_shift[4][6] ),
    .S(_11332_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _24039_ (.A0(\systolic_inst.B_shift[8][7] ),
    .A1(\B_in[39] ),
    .S(_00008_),
    .X(_10537_));
 sky130_fd_sc_hd__mux2_1 _24040_ (.A0(_10537_),
    .A1(\systolic_inst.B_shift[4][7] ),
    .S(_11332_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _24041_ (.A0(\systolic_inst.B_shift[4][0] ),
    .A1(\B_in[0] ),
    .S(_00008_),
    .X(_10538_));
 sky130_fd_sc_hd__mux2_1 _24042_ (.A0(_10538_),
    .A1(\systolic_inst.B_shift[0][0] ),
    .S(_11332_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _24043_ (.A0(\systolic_inst.B_shift[4][1] ),
    .A1(\B_in[1] ),
    .S(_00008_),
    .X(_10539_));
 sky130_fd_sc_hd__mux2_1 _24044_ (.A0(_10539_),
    .A1(\systolic_inst.B_shift[0][1] ),
    .S(_11332_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _24045_ (.A0(\systolic_inst.B_shift[4][2] ),
    .A1(\B_in[2] ),
    .S(_00008_),
    .X(_10540_));
 sky130_fd_sc_hd__mux2_1 _24046_ (.A0(_10540_),
    .A1(\systolic_inst.B_shift[0][2] ),
    .S(_11332_),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _24047_ (.A0(\systolic_inst.B_shift[4][3] ),
    .A1(\B_in[3] ),
    .S(_00008_),
    .X(_10541_));
 sky130_fd_sc_hd__mux2_1 _24048_ (.A0(_10541_),
    .A1(\systolic_inst.B_shift[0][3] ),
    .S(_11332_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _24049_ (.A0(\systolic_inst.B_shift[4][4] ),
    .A1(\B_in[4] ),
    .S(_00008_),
    .X(_10542_));
 sky130_fd_sc_hd__mux2_1 _24050_ (.A0(_10542_),
    .A1(\systolic_inst.B_shift[0][4] ),
    .S(_11332_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _24051_ (.A0(\systolic_inst.B_shift[4][5] ),
    .A1(\B_in[5] ),
    .S(_00008_),
    .X(_10543_));
 sky130_fd_sc_hd__mux2_1 _24052_ (.A0(_10543_),
    .A1(\systolic_inst.B_shift[0][5] ),
    .S(_11332_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _24053_ (.A0(\systolic_inst.B_shift[4][6] ),
    .A1(\B_in[6] ),
    .S(_00008_),
    .X(_10544_));
 sky130_fd_sc_hd__mux2_1 _24054_ (.A0(_10544_),
    .A1(\systolic_inst.B_shift[0][6] ),
    .S(_11332_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _24055_ (.A0(\systolic_inst.B_shift[4][7] ),
    .A1(\B_in[7] ),
    .S(_00008_),
    .X(_10545_));
 sky130_fd_sc_hd__mux2_1 _24056_ (.A0(_10545_),
    .A1(\systolic_inst.B_shift[0][7] ),
    .S(_11332_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _24057_ (.A0(\systolic_inst.B_shift[19][0] ),
    .A1(\B_in[24] ),
    .S(_00008_),
    .X(_10546_));
 sky130_fd_sc_hd__mux2_1 _24058_ (.A0(_10546_),
    .A1(\systolic_inst.B_shift[15][0] ),
    .S(_11332_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _24059_ (.A0(\systolic_inst.B_shift[19][1] ),
    .A1(\B_in[25] ),
    .S(_00008_),
    .X(_10547_));
 sky130_fd_sc_hd__mux2_1 _24060_ (.A0(_10547_),
    .A1(\systolic_inst.B_shift[15][1] ),
    .S(_11332_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _24061_ (.A0(\systolic_inst.B_shift[19][2] ),
    .A1(\B_in[26] ),
    .S(_00008_),
    .X(_10548_));
 sky130_fd_sc_hd__mux2_1 _24062_ (.A0(_10548_),
    .A1(\systolic_inst.B_shift[15][2] ),
    .S(_11332_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _24063_ (.A0(\systolic_inst.B_shift[19][3] ),
    .A1(\B_in[27] ),
    .S(_00008_),
    .X(_10549_));
 sky130_fd_sc_hd__mux2_1 _24064_ (.A0(_10549_),
    .A1(\systolic_inst.B_shift[15][3] ),
    .S(_11332_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _24065_ (.A0(\systolic_inst.B_shift[19][4] ),
    .A1(\B_in[28] ),
    .S(_00008_),
    .X(_10550_));
 sky130_fd_sc_hd__mux2_1 _24066_ (.A0(_10550_),
    .A1(\systolic_inst.B_shift[15][4] ),
    .S(_11332_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _24067_ (.A0(\systolic_inst.B_shift[19][5] ),
    .A1(\B_in[29] ),
    .S(_00008_),
    .X(_10551_));
 sky130_fd_sc_hd__mux2_1 _24068_ (.A0(_10551_),
    .A1(\systolic_inst.B_shift[15][5] ),
    .S(_11332_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _24069_ (.A0(\systolic_inst.B_shift[19][6] ),
    .A1(\B_in[30] ),
    .S(_00008_),
    .X(_10552_));
 sky130_fd_sc_hd__mux2_1 _24070_ (.A0(_10552_),
    .A1(\systolic_inst.B_shift[15][6] ),
    .S(_11332_),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _24071_ (.A0(\systolic_inst.B_shift[19][7] ),
    .A1(\B_in[31] ),
    .S(_00008_),
    .X(_10553_));
 sky130_fd_sc_hd__mux2_1 _24072_ (.A0(_10553_),
    .A1(\systolic_inst.B_shift[15][7] ),
    .S(_11332_),
    .X(_02065_));
 sky130_fd_sc_hd__a22o_2 _24073_ (.A1(\systolic_inst.B_shift[3][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[7][0] ),
    .X(_02066_));
 sky130_fd_sc_hd__a22o_2 _24074_ (.A1(\systolic_inst.B_shift[3][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[7][1] ),
    .X(_02067_));
 sky130_fd_sc_hd__a22o_2 _24075_ (.A1(\systolic_inst.B_shift[3][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[7][2] ),
    .X(_02068_));
 sky130_fd_sc_hd__a22o_2 _24076_ (.A1(\systolic_inst.B_shift[3][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[7][3] ),
    .X(_02069_));
 sky130_fd_sc_hd__a22o_2 _24077_ (.A1(\systolic_inst.B_shift[3][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[7][4] ),
    .X(_02070_));
 sky130_fd_sc_hd__a22o_2 _24078_ (.A1(\systolic_inst.B_shift[3][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[7][5] ),
    .X(_02071_));
 sky130_fd_sc_hd__a22o_2 _24079_ (.A1(\systolic_inst.B_shift[3][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[7][6] ),
    .X(_02072_));
 sky130_fd_sc_hd__a22o_2 _24080_ (.A1(\systolic_inst.B_shift[3][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[7][7] ),
    .X(_02073_));
 sky130_fd_sc_hd__a22o_2 _24081_ (.A1(\systolic_inst.B_shift[2][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[6][0] ),
    .X(_02074_));
 sky130_fd_sc_hd__a22o_2 _24082_ (.A1(\systolic_inst.B_shift[2][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[6][1] ),
    .X(_02075_));
 sky130_fd_sc_hd__a22o_2 _24083_ (.A1(\systolic_inst.B_shift[2][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[6][2] ),
    .X(_02076_));
 sky130_fd_sc_hd__a22o_2 _24084_ (.A1(\systolic_inst.B_shift[2][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[6][3] ),
    .X(_02077_));
 sky130_fd_sc_hd__a22o_2 _24085_ (.A1(\systolic_inst.B_shift[2][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[6][4] ),
    .X(_02078_));
 sky130_fd_sc_hd__a22o_2 _24086_ (.A1(\systolic_inst.B_shift[2][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[6][5] ),
    .X(_02079_));
 sky130_fd_sc_hd__a22o_2 _24087_ (.A1(\systolic_inst.B_shift[2][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[6][6] ),
    .X(_02080_));
 sky130_fd_sc_hd__a22o_2 _24088_ (.A1(\systolic_inst.B_shift[2][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[6][7] ),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_1 _24089_ (.A0(\systolic_inst.B_shift[23][0] ),
    .A1(\B_in[56] ),
    .S(_00008_),
    .X(_10554_));
 sky130_fd_sc_hd__mux2_1 _24090_ (.A0(_10554_),
    .A1(\systolic_inst.B_shift[19][0] ),
    .S(_11332_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _24091_ (.A0(\systolic_inst.B_shift[23][1] ),
    .A1(\B_in[57] ),
    .S(_00008_),
    .X(_10555_));
 sky130_fd_sc_hd__mux2_1 _24092_ (.A0(_10555_),
    .A1(\systolic_inst.B_shift[19][1] ),
    .S(_11332_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_1 _24093_ (.A0(\systolic_inst.B_shift[23][2] ),
    .A1(\B_in[58] ),
    .S(_00008_),
    .X(_10556_));
 sky130_fd_sc_hd__mux2_1 _24094_ (.A0(_10556_),
    .A1(\systolic_inst.B_shift[19][2] ),
    .S(_11332_),
    .X(_02084_));
 sky130_fd_sc_hd__mux2_1 _24095_ (.A0(\systolic_inst.B_shift[23][3] ),
    .A1(\B_in[59] ),
    .S(_00008_),
    .X(_10557_));
 sky130_fd_sc_hd__mux2_1 _24096_ (.A0(_10557_),
    .A1(\systolic_inst.B_shift[19][3] ),
    .S(_11332_),
    .X(_02085_));
 sky130_fd_sc_hd__mux2_1 _24097_ (.A0(\systolic_inst.B_shift[23][4] ),
    .A1(\B_in[60] ),
    .S(_00008_),
    .X(_10558_));
 sky130_fd_sc_hd__mux2_1 _24098_ (.A0(_10558_),
    .A1(\systolic_inst.B_shift[19][4] ),
    .S(_11332_),
    .X(_02086_));
 sky130_fd_sc_hd__mux2_1 _24099_ (.A0(\systolic_inst.B_shift[23][5] ),
    .A1(\B_in[61] ),
    .S(_00008_),
    .X(_10559_));
 sky130_fd_sc_hd__mux2_1 _24100_ (.A0(_10559_),
    .A1(\systolic_inst.B_shift[19][5] ),
    .S(_11332_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_1 _24101_ (.A0(\systolic_inst.B_shift[23][6] ),
    .A1(\B_in[62] ),
    .S(_00008_),
    .X(_10560_));
 sky130_fd_sc_hd__mux2_1 _24102_ (.A0(_10560_),
    .A1(\systolic_inst.B_shift[19][6] ),
    .S(_11332_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _24103_ (.A0(\systolic_inst.B_shift[23][7] ),
    .A1(\B_in[63] ),
    .S(_00008_),
    .X(_10561_));
 sky130_fd_sc_hd__mux2_1 _24104_ (.A0(_10561_),
    .A1(\systolic_inst.B_shift[19][7] ),
    .S(_11332_),
    .X(_02089_));
 sky130_fd_sc_hd__a22o_2 _24105_ (.A1(\systolic_inst.B_shift[1][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[5][0] ),
    .X(_02090_));
 sky130_fd_sc_hd__a22o_2 _24106_ (.A1(\systolic_inst.B_shift[1][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[5][1] ),
    .X(_02091_));
 sky130_fd_sc_hd__a22o_2 _24107_ (.A1(\systolic_inst.B_shift[1][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[5][2] ),
    .X(_02092_));
 sky130_fd_sc_hd__a22o_2 _24108_ (.A1(\systolic_inst.B_shift[1][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[5][3] ),
    .X(_02093_));
 sky130_fd_sc_hd__a22o_2 _24109_ (.A1(\systolic_inst.B_shift[1][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[5][4] ),
    .X(_02094_));
 sky130_fd_sc_hd__a22o_2 _24110_ (.A1(\systolic_inst.B_shift[1][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[5][5] ),
    .X(_02095_));
 sky130_fd_sc_hd__a22o_2 _24111_ (.A1(\systolic_inst.B_shift[1][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[5][6] ),
    .X(_02096_));
 sky130_fd_sc_hd__a22o_2 _24112_ (.A1(\systolic_inst.B_shift[1][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.B_shift[5][7] ),
    .X(_02097_));
 sky130_fd_sc_hd__a22o_2 _24113_ (.A1(\systolic_inst.B_shift[27][0] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[120] ),
    .X(_02098_));
 sky130_fd_sc_hd__a22o_2 _24114_ (.A1(\systolic_inst.B_shift[27][1] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[121] ),
    .X(_02099_));
 sky130_fd_sc_hd__a22o_2 _24115_ (.A1(\systolic_inst.B_shift[27][2] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[122] ),
    .X(_02100_));
 sky130_fd_sc_hd__a22o_2 _24116_ (.A1(\systolic_inst.B_shift[27][3] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[123] ),
    .X(_02101_));
 sky130_fd_sc_hd__a22o_2 _24117_ (.A1(\systolic_inst.B_shift[27][4] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[124] ),
    .X(_02102_));
 sky130_fd_sc_hd__a22o_2 _24118_ (.A1(\systolic_inst.B_shift[27][5] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[125] ),
    .X(_02103_));
 sky130_fd_sc_hd__a22o_2 _24119_ (.A1(\systolic_inst.B_shift[27][6] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[126] ),
    .X(_02104_));
 sky130_fd_sc_hd__a22o_2 _24120_ (.A1(\systolic_inst.B_shift[27][7] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[127] ),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _24121_ (.A0(\systolic_inst.A_shift[30][0] ),
    .A1(\A_in[112] ),
    .S(_00008_),
    .X(_10562_));
 sky130_fd_sc_hd__mux2_1 _24122_ (.A0(_10562_),
    .A1(\systolic_inst.A_shift[29][0] ),
    .S(_11332_),
    .X(_02106_));
 sky130_fd_sc_hd__mux2_1 _24123_ (.A0(\systolic_inst.A_shift[30][1] ),
    .A1(\A_in[113] ),
    .S(_00008_),
    .X(_10563_));
 sky130_fd_sc_hd__mux2_1 _24124_ (.A0(_10563_),
    .A1(\systolic_inst.A_shift[29][1] ),
    .S(_11332_),
    .X(_02107_));
 sky130_fd_sc_hd__mux2_1 _24125_ (.A0(\systolic_inst.A_shift[30][2] ),
    .A1(\A_in[114] ),
    .S(_00008_),
    .X(_10564_));
 sky130_fd_sc_hd__mux2_1 _24126_ (.A0(_10564_),
    .A1(\systolic_inst.A_shift[29][2] ),
    .S(_11332_),
    .X(_02108_));
 sky130_fd_sc_hd__mux2_1 _24127_ (.A0(\systolic_inst.A_shift[30][3] ),
    .A1(\A_in[115] ),
    .S(_00008_),
    .X(_10565_));
 sky130_fd_sc_hd__mux2_1 _24128_ (.A0(_10565_),
    .A1(\systolic_inst.A_shift[29][3] ),
    .S(_11332_),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _24129_ (.A0(\systolic_inst.A_shift[30][4] ),
    .A1(\A_in[116] ),
    .S(_00008_),
    .X(_10566_));
 sky130_fd_sc_hd__mux2_1 _24130_ (.A0(_10566_),
    .A1(\systolic_inst.A_shift[29][4] ),
    .S(_11332_),
    .X(_02110_));
 sky130_fd_sc_hd__mux2_1 _24131_ (.A0(\systolic_inst.A_shift[30][5] ),
    .A1(\A_in[117] ),
    .S(_00008_),
    .X(_10567_));
 sky130_fd_sc_hd__mux2_1 _24132_ (.A0(_10567_),
    .A1(\systolic_inst.A_shift[29][5] ),
    .S(_11332_),
    .X(_02111_));
 sky130_fd_sc_hd__mux2_1 _24133_ (.A0(\systolic_inst.A_shift[30][6] ),
    .A1(\A_in[118] ),
    .S(_00008_),
    .X(_10568_));
 sky130_fd_sc_hd__mux2_1 _24134_ (.A0(_10568_),
    .A1(\systolic_inst.A_shift[29][6] ),
    .S(_11332_),
    .X(_02112_));
 sky130_fd_sc_hd__mux2_1 _24135_ (.A0(\systolic_inst.A_shift[30][7] ),
    .A1(\A_in[119] ),
    .S(_00008_),
    .X(_10569_));
 sky130_fd_sc_hd__mux2_1 _24136_ (.A0(_10569_),
    .A1(\systolic_inst.A_shift[29][7] ),
    .S(_11332_),
    .X(_02113_));
 sky130_fd_sc_hd__mux2_1 _24137_ (.A0(\systolic_inst.A_shift[29][0] ),
    .A1(\A_in[104] ),
    .S(_00008_),
    .X(_10570_));
 sky130_fd_sc_hd__mux2_1 _24138_ (.A0(_10570_),
    .A1(\systolic_inst.A_shift[28][0] ),
    .S(_11332_),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _24139_ (.A0(\systolic_inst.A_shift[29][1] ),
    .A1(\A_in[105] ),
    .S(_00008_),
    .X(_10571_));
 sky130_fd_sc_hd__mux2_1 _24140_ (.A0(_10571_),
    .A1(\systolic_inst.A_shift[28][1] ),
    .S(_11332_),
    .X(_02115_));
 sky130_fd_sc_hd__mux2_1 _24141_ (.A0(\systolic_inst.A_shift[29][2] ),
    .A1(\A_in[106] ),
    .S(_00008_),
    .X(_10572_));
 sky130_fd_sc_hd__mux2_1 _24142_ (.A0(_10572_),
    .A1(\systolic_inst.A_shift[28][2] ),
    .S(_11332_),
    .X(_02116_));
 sky130_fd_sc_hd__mux2_1 _24143_ (.A0(\systolic_inst.A_shift[29][3] ),
    .A1(\A_in[107] ),
    .S(_00008_),
    .X(_10573_));
 sky130_fd_sc_hd__mux2_1 _24144_ (.A0(_10573_),
    .A1(\systolic_inst.A_shift[28][3] ),
    .S(_11332_),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _24145_ (.A0(\systolic_inst.A_shift[29][4] ),
    .A1(\A_in[108] ),
    .S(_00008_),
    .X(_10574_));
 sky130_fd_sc_hd__mux2_1 _24146_ (.A0(_10574_),
    .A1(\systolic_inst.A_shift[28][4] ),
    .S(_11332_),
    .X(_02118_));
 sky130_fd_sc_hd__mux2_1 _24147_ (.A0(\systolic_inst.A_shift[29][5] ),
    .A1(\A_in[109] ),
    .S(_00008_),
    .X(_10575_));
 sky130_fd_sc_hd__mux2_1 _24148_ (.A0(_10575_),
    .A1(\systolic_inst.A_shift[28][5] ),
    .S(_11332_),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _24149_ (.A0(\systolic_inst.A_shift[29][6] ),
    .A1(\A_in[110] ),
    .S(_00008_),
    .X(_10576_));
 sky130_fd_sc_hd__mux2_1 _24150_ (.A0(_10576_),
    .A1(\systolic_inst.A_shift[28][6] ),
    .S(_11332_),
    .X(_02120_));
 sky130_fd_sc_hd__mux2_1 _24151_ (.A0(\systolic_inst.A_shift[29][7] ),
    .A1(\A_in[111] ),
    .S(_00008_),
    .X(_10577_));
 sky130_fd_sc_hd__mux2_1 _24152_ (.A0(_10577_),
    .A1(\systolic_inst.A_shift[28][7] ),
    .S(_11332_),
    .X(_02121_));
 sky130_fd_sc_hd__mux2_1 _24153_ (.A0(\systolic_inst.A_shift[28][0] ),
    .A1(\A_in[96] ),
    .S(_00008_),
    .X(_10578_));
 sky130_fd_sc_hd__mux2_1 _24154_ (.A0(_10578_),
    .A1(\systolic_inst.A_shift[27][0] ),
    .S(_11332_),
    .X(_02122_));
 sky130_fd_sc_hd__mux2_1 _24155_ (.A0(\systolic_inst.A_shift[28][1] ),
    .A1(\A_in[97] ),
    .S(_00008_),
    .X(_10579_));
 sky130_fd_sc_hd__mux2_1 _24156_ (.A0(_10579_),
    .A1(\systolic_inst.A_shift[27][1] ),
    .S(_11332_),
    .X(_02123_));
 sky130_fd_sc_hd__mux2_1 _24157_ (.A0(\systolic_inst.A_shift[28][2] ),
    .A1(\A_in[98] ),
    .S(_00008_),
    .X(_10580_));
 sky130_fd_sc_hd__mux2_1 _24158_ (.A0(_10580_),
    .A1(\systolic_inst.A_shift[27][2] ),
    .S(_11332_),
    .X(_02124_));
 sky130_fd_sc_hd__mux2_1 _24159_ (.A0(\systolic_inst.A_shift[28][3] ),
    .A1(\A_in[99] ),
    .S(_00008_),
    .X(_10581_));
 sky130_fd_sc_hd__mux2_1 _24160_ (.A0(_10581_),
    .A1(\systolic_inst.A_shift[27][3] ),
    .S(_11332_),
    .X(_02125_));
 sky130_fd_sc_hd__mux2_1 _24161_ (.A0(\systolic_inst.A_shift[28][4] ),
    .A1(\A_in[100] ),
    .S(_00008_),
    .X(_10582_));
 sky130_fd_sc_hd__mux2_1 _24162_ (.A0(_10582_),
    .A1(\systolic_inst.A_shift[27][4] ),
    .S(_11332_),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _24163_ (.A0(\systolic_inst.A_shift[28][5] ),
    .A1(\A_in[101] ),
    .S(_00008_),
    .X(_10583_));
 sky130_fd_sc_hd__mux2_1 _24164_ (.A0(_10583_),
    .A1(\systolic_inst.A_shift[27][5] ),
    .S(_11332_),
    .X(_02127_));
 sky130_fd_sc_hd__mux2_1 _24165_ (.A0(\systolic_inst.A_shift[28][6] ),
    .A1(\A_in[102] ),
    .S(_00008_),
    .X(_10584_));
 sky130_fd_sc_hd__mux2_1 _24166_ (.A0(_10584_),
    .A1(\systolic_inst.A_shift[27][6] ),
    .S(_11332_),
    .X(_02128_));
 sky130_fd_sc_hd__mux2_1 _24167_ (.A0(\systolic_inst.A_shift[28][7] ),
    .A1(\A_in[103] ),
    .S(_00008_),
    .X(_10585_));
 sky130_fd_sc_hd__mux2_1 _24168_ (.A0(_10585_),
    .A1(\systolic_inst.A_shift[27][7] ),
    .S(_11332_),
    .X(_02129_));
 sky130_fd_sc_hd__a22o_2 _24169_ (.A1(\systolic_inst.A_shift[26][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[27][0] ),
    .X(_02130_));
 sky130_fd_sc_hd__a22o_2 _24170_ (.A1(\systolic_inst.A_shift[26][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[27][1] ),
    .X(_02131_));
 sky130_fd_sc_hd__a22o_2 _24171_ (.A1(\systolic_inst.A_shift[26][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[27][2] ),
    .X(_02132_));
 sky130_fd_sc_hd__a22o_2 _24172_ (.A1(\systolic_inst.A_shift[26][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[27][3] ),
    .X(_02133_));
 sky130_fd_sc_hd__a22o_2 _24173_ (.A1(\systolic_inst.A_shift[26][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[27][4] ),
    .X(_02134_));
 sky130_fd_sc_hd__a22o_2 _24174_ (.A1(\systolic_inst.A_shift[26][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[27][5] ),
    .X(_02135_));
 sky130_fd_sc_hd__a22o_2 _24175_ (.A1(\systolic_inst.A_shift[26][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[27][6] ),
    .X(_02136_));
 sky130_fd_sc_hd__a22o_2 _24176_ (.A1(\systolic_inst.A_shift[26][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[27][7] ),
    .X(_02137_));
 sky130_fd_sc_hd__a22o_2 _24177_ (.A1(\systolic_inst.A_shift[25][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[26][0] ),
    .X(_02138_));
 sky130_fd_sc_hd__a22o_2 _24178_ (.A1(\systolic_inst.A_shift[25][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[26][1] ),
    .X(_02139_));
 sky130_fd_sc_hd__a22o_2 _24179_ (.A1(\systolic_inst.A_shift[25][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[26][2] ),
    .X(_02140_));
 sky130_fd_sc_hd__a22o_2 _24180_ (.A1(\systolic_inst.A_shift[25][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[26][3] ),
    .X(_02141_));
 sky130_fd_sc_hd__a22o_2 _24181_ (.A1(\systolic_inst.A_shift[25][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[26][4] ),
    .X(_02142_));
 sky130_fd_sc_hd__a22o_2 _24182_ (.A1(\systolic_inst.A_shift[25][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[26][5] ),
    .X(_02143_));
 sky130_fd_sc_hd__a22o_2 _24183_ (.A1(\systolic_inst.A_shift[25][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[26][6] ),
    .X(_02144_));
 sky130_fd_sc_hd__a22o_2 _24184_ (.A1(\systolic_inst.A_shift[25][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[26][7] ),
    .X(_02145_));
 sky130_fd_sc_hd__a22o_2 _24185_ (.A1(\systolic_inst.A_shift[24][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[25][0] ),
    .X(_02146_));
 sky130_fd_sc_hd__a22o_2 _24186_ (.A1(\systolic_inst.A_shift[24][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[25][1] ),
    .X(_02147_));
 sky130_fd_sc_hd__a22o_2 _24187_ (.A1(\systolic_inst.A_shift[24][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[25][2] ),
    .X(_02148_));
 sky130_fd_sc_hd__a22o_2 _24188_ (.A1(\systolic_inst.A_shift[24][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[25][3] ),
    .X(_02149_));
 sky130_fd_sc_hd__a22o_2 _24189_ (.A1(\systolic_inst.A_shift[24][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[25][4] ),
    .X(_02150_));
 sky130_fd_sc_hd__a22o_2 _24190_ (.A1(\systolic_inst.A_shift[24][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[25][5] ),
    .X(_02151_));
 sky130_fd_sc_hd__a22o_2 _24191_ (.A1(\systolic_inst.A_shift[24][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[25][6] ),
    .X(_02152_));
 sky130_fd_sc_hd__a22o_2 _24192_ (.A1(\systolic_inst.A_shift[24][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[25][7] ),
    .X(_02153_));
 sky130_fd_sc_hd__a22o_2 _24193_ (.A1(\systolic_inst.B_shift[22][0] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[112] ),
    .X(_02154_));
 sky130_fd_sc_hd__a22o_2 _24194_ (.A1(\systolic_inst.B_shift[22][1] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[113] ),
    .X(_02155_));
 sky130_fd_sc_hd__a22o_2 _24195_ (.A1(\systolic_inst.B_shift[22][2] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[114] ),
    .X(_02156_));
 sky130_fd_sc_hd__a22o_2 _24196_ (.A1(\systolic_inst.B_shift[22][3] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[115] ),
    .X(_02157_));
 sky130_fd_sc_hd__a22o_2 _24197_ (.A1(\systolic_inst.B_shift[22][4] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[116] ),
    .X(_02158_));
 sky130_fd_sc_hd__a22o_2 _24198_ (.A1(\systolic_inst.B_shift[22][5] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[117] ),
    .X(_02159_));
 sky130_fd_sc_hd__a22o_2 _24199_ (.A1(\systolic_inst.B_shift[22][6] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[118] ),
    .X(_02160_));
 sky130_fd_sc_hd__a22o_2 _24200_ (.A1(\systolic_inst.B_shift[22][7] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[119] ),
    .X(_02161_));
 sky130_fd_sc_hd__mux2_1 _24201_ (.A0(\systolic_inst.A_shift[21][0] ),
    .A1(\A_in[80] ),
    .S(_00008_),
    .X(_10586_));
 sky130_fd_sc_hd__mux2_1 _24202_ (.A0(_10586_),
    .A1(\systolic_inst.A_shift[20][0] ),
    .S(_11332_),
    .X(_02162_));
 sky130_fd_sc_hd__mux2_1 _24203_ (.A0(\systolic_inst.A_shift[21][1] ),
    .A1(\A_in[81] ),
    .S(_00008_),
    .X(_10587_));
 sky130_fd_sc_hd__mux2_1 _24204_ (.A0(_10587_),
    .A1(\systolic_inst.A_shift[20][1] ),
    .S(_11332_),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_1 _24205_ (.A0(\systolic_inst.A_shift[21][2] ),
    .A1(\A_in[82] ),
    .S(_00008_),
    .X(_10588_));
 sky130_fd_sc_hd__mux2_1 _24206_ (.A0(_10588_),
    .A1(\systolic_inst.A_shift[20][2] ),
    .S(_11332_),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_1 _24207_ (.A0(\systolic_inst.A_shift[21][3] ),
    .A1(\A_in[83] ),
    .S(_00008_),
    .X(_10589_));
 sky130_fd_sc_hd__mux2_1 _24208_ (.A0(_10589_),
    .A1(\systolic_inst.A_shift[20][3] ),
    .S(_11332_),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_1 _24209_ (.A0(\systolic_inst.A_shift[21][4] ),
    .A1(\A_in[84] ),
    .S(_00008_),
    .X(_10590_));
 sky130_fd_sc_hd__mux2_1 _24210_ (.A0(_10590_),
    .A1(\systolic_inst.A_shift[20][4] ),
    .S(_11332_),
    .X(_02166_));
 sky130_fd_sc_hd__mux2_1 _24211_ (.A0(\systolic_inst.A_shift[21][5] ),
    .A1(\A_in[85] ),
    .S(_00008_),
    .X(_10591_));
 sky130_fd_sc_hd__mux2_1 _24212_ (.A0(_10591_),
    .A1(\systolic_inst.A_shift[20][5] ),
    .S(_11332_),
    .X(_02167_));
 sky130_fd_sc_hd__mux2_1 _24213_ (.A0(\systolic_inst.A_shift[21][6] ),
    .A1(\A_in[86] ),
    .S(_00008_),
    .X(_10592_));
 sky130_fd_sc_hd__mux2_1 _24214_ (.A0(_10592_),
    .A1(\systolic_inst.A_shift[20][6] ),
    .S(_11332_),
    .X(_02168_));
 sky130_fd_sc_hd__mux2_1 _24215_ (.A0(\systolic_inst.A_shift[21][7] ),
    .A1(\A_in[87] ),
    .S(_00008_),
    .X(_10593_));
 sky130_fd_sc_hd__mux2_1 _24216_ (.A0(_10593_),
    .A1(\systolic_inst.A_shift[20][7] ),
    .S(_11332_),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_1 _24217_ (.A0(\systolic_inst.A_shift[20][0] ),
    .A1(\A_in[72] ),
    .S(_00008_),
    .X(_10594_));
 sky130_fd_sc_hd__mux2_1 _24218_ (.A0(_10594_),
    .A1(\systolic_inst.A_shift[19][0] ),
    .S(_11332_),
    .X(_02170_));
 sky130_fd_sc_hd__mux2_1 _24219_ (.A0(\systolic_inst.A_shift[20][1] ),
    .A1(\A_in[73] ),
    .S(_00008_),
    .X(_10595_));
 sky130_fd_sc_hd__mux2_1 _24220_ (.A0(_10595_),
    .A1(\systolic_inst.A_shift[19][1] ),
    .S(_11332_),
    .X(_02171_));
 sky130_fd_sc_hd__mux2_1 _24221_ (.A0(\systolic_inst.A_shift[20][2] ),
    .A1(\A_in[74] ),
    .S(_00008_),
    .X(_10596_));
 sky130_fd_sc_hd__mux2_1 _24222_ (.A0(_10596_),
    .A1(\systolic_inst.A_shift[19][2] ),
    .S(_11332_),
    .X(_02172_));
 sky130_fd_sc_hd__mux2_1 _24223_ (.A0(\systolic_inst.A_shift[20][3] ),
    .A1(\A_in[75] ),
    .S(_00008_),
    .X(_10597_));
 sky130_fd_sc_hd__mux2_1 _24224_ (.A0(_10597_),
    .A1(\systolic_inst.A_shift[19][3] ),
    .S(_11332_),
    .X(_02173_));
 sky130_fd_sc_hd__mux2_1 _24225_ (.A0(\systolic_inst.A_shift[20][4] ),
    .A1(\A_in[76] ),
    .S(_00008_),
    .X(_10598_));
 sky130_fd_sc_hd__mux2_1 _24226_ (.A0(_10598_),
    .A1(\systolic_inst.A_shift[19][4] ),
    .S(_11332_),
    .X(_02174_));
 sky130_fd_sc_hd__mux2_1 _24227_ (.A0(\systolic_inst.A_shift[20][5] ),
    .A1(\A_in[77] ),
    .S(_00008_),
    .X(_10599_));
 sky130_fd_sc_hd__mux2_1 _24228_ (.A0(_10599_),
    .A1(\systolic_inst.A_shift[19][5] ),
    .S(_11332_),
    .X(_02175_));
 sky130_fd_sc_hd__mux2_1 _24229_ (.A0(\systolic_inst.A_shift[20][6] ),
    .A1(\A_in[78] ),
    .S(_00008_),
    .X(_10600_));
 sky130_fd_sc_hd__mux2_1 _24230_ (.A0(_10600_),
    .A1(\systolic_inst.A_shift[19][6] ),
    .S(_11332_),
    .X(_02176_));
 sky130_fd_sc_hd__mux2_1 _24231_ (.A0(\systolic_inst.A_shift[20][7] ),
    .A1(\A_in[79] ),
    .S(_00008_),
    .X(_10601_));
 sky130_fd_sc_hd__mux2_1 _24232_ (.A0(_10601_),
    .A1(\systolic_inst.A_shift[19][7] ),
    .S(_11332_),
    .X(_02177_));
 sky130_fd_sc_hd__mux2_1 _24233_ (.A0(\systolic_inst.A_shift[19][0] ),
    .A1(\A_in[64] ),
    .S(_00008_),
    .X(_10602_));
 sky130_fd_sc_hd__mux2_1 _24234_ (.A0(_10602_),
    .A1(\systolic_inst.A_shift[18][0] ),
    .S(_11332_),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _24235_ (.A0(\systolic_inst.A_shift[19][1] ),
    .A1(\A_in[65] ),
    .S(_00008_),
    .X(_10603_));
 sky130_fd_sc_hd__mux2_1 _24236_ (.A0(_10603_),
    .A1(\systolic_inst.A_shift[18][1] ),
    .S(_11332_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _24237_ (.A0(\systolic_inst.A_shift[19][2] ),
    .A1(\A_in[66] ),
    .S(_00008_),
    .X(_10604_));
 sky130_fd_sc_hd__mux2_1 _24238_ (.A0(_10604_),
    .A1(\systolic_inst.A_shift[18][2] ),
    .S(_11332_),
    .X(_02180_));
 sky130_fd_sc_hd__mux2_1 _24239_ (.A0(\systolic_inst.A_shift[19][3] ),
    .A1(\A_in[67] ),
    .S(_00008_),
    .X(_10605_));
 sky130_fd_sc_hd__mux2_1 _24240_ (.A0(_10605_),
    .A1(\systolic_inst.A_shift[18][3] ),
    .S(_11332_),
    .X(_02181_));
 sky130_fd_sc_hd__mux2_1 _24241_ (.A0(\systolic_inst.A_shift[19][4] ),
    .A1(\A_in[68] ),
    .S(_00008_),
    .X(_10606_));
 sky130_fd_sc_hd__mux2_1 _24242_ (.A0(_10606_),
    .A1(\systolic_inst.A_shift[18][4] ),
    .S(_11332_),
    .X(_02182_));
 sky130_fd_sc_hd__mux2_1 _24243_ (.A0(\systolic_inst.A_shift[19][5] ),
    .A1(\A_in[69] ),
    .S(_00008_),
    .X(_10607_));
 sky130_fd_sc_hd__mux2_1 _24244_ (.A0(_10607_),
    .A1(\systolic_inst.A_shift[18][5] ),
    .S(_11332_),
    .X(_02183_));
 sky130_fd_sc_hd__mux2_1 _24245_ (.A0(\systolic_inst.A_shift[19][6] ),
    .A1(\A_in[70] ),
    .S(_00008_),
    .X(_10608_));
 sky130_fd_sc_hd__mux2_1 _24246_ (.A0(_10608_),
    .A1(\systolic_inst.A_shift[18][6] ),
    .S(_11332_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _24247_ (.A0(\systolic_inst.A_shift[19][7] ),
    .A1(\A_in[71] ),
    .S(_00008_),
    .X(_10609_));
 sky130_fd_sc_hd__mux2_1 _24248_ (.A0(_10609_),
    .A1(\systolic_inst.A_shift[18][7] ),
    .S(_11332_),
    .X(_02185_));
 sky130_fd_sc_hd__a22o_2 _24249_ (.A1(\systolic_inst.A_shift[17][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[18][0] ),
    .X(_02186_));
 sky130_fd_sc_hd__a22o_2 _24250_ (.A1(\systolic_inst.A_shift[17][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[18][1] ),
    .X(_02187_));
 sky130_fd_sc_hd__a22o_2 _24251_ (.A1(\systolic_inst.A_shift[17][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[18][2] ),
    .X(_02188_));
 sky130_fd_sc_hd__a22o_2 _24252_ (.A1(\systolic_inst.A_shift[17][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[18][3] ),
    .X(_02189_));
 sky130_fd_sc_hd__a22o_2 _24253_ (.A1(\systolic_inst.A_shift[17][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[18][4] ),
    .X(_02190_));
 sky130_fd_sc_hd__a22o_2 _24254_ (.A1(\systolic_inst.A_shift[17][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[18][5] ),
    .X(_02191_));
 sky130_fd_sc_hd__a22o_2 _24255_ (.A1(\systolic_inst.A_shift[17][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[18][6] ),
    .X(_02192_));
 sky130_fd_sc_hd__a22o_2 _24256_ (.A1(\systolic_inst.A_shift[17][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[18][7] ),
    .X(_02193_));
 sky130_fd_sc_hd__a22o_2 _24257_ (.A1(\systolic_inst.A_shift[16][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[17][0] ),
    .X(_02194_));
 sky130_fd_sc_hd__a22o_2 _24258_ (.A1(\systolic_inst.A_shift[16][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[17][1] ),
    .X(_02195_));
 sky130_fd_sc_hd__a22o_2 _24259_ (.A1(\systolic_inst.A_shift[16][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[17][2] ),
    .X(_02196_));
 sky130_fd_sc_hd__a22o_2 _24260_ (.A1(\systolic_inst.A_shift[16][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[17][3] ),
    .X(_02197_));
 sky130_fd_sc_hd__a22o_2 _24261_ (.A1(\systolic_inst.A_shift[16][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[17][4] ),
    .X(_02198_));
 sky130_fd_sc_hd__a22o_2 _24262_ (.A1(\systolic_inst.A_shift[16][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[17][5] ),
    .X(_02199_));
 sky130_fd_sc_hd__a22o_2 _24263_ (.A1(\systolic_inst.A_shift[16][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[17][6] ),
    .X(_02200_));
 sky130_fd_sc_hd__a22o_2 _24264_ (.A1(\systolic_inst.A_shift[16][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[17][7] ),
    .X(_02201_));
 sky130_fd_sc_hd__a22o_2 _24265_ (.A1(\systolic_inst.B_shift[17][0] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[104] ),
    .X(_02202_));
 sky130_fd_sc_hd__a22o_2 _24266_ (.A1(\systolic_inst.B_shift[17][1] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[105] ),
    .X(_02203_));
 sky130_fd_sc_hd__a22o_2 _24267_ (.A1(\systolic_inst.B_shift[17][2] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[106] ),
    .X(_02204_));
 sky130_fd_sc_hd__a22o_2 _24268_ (.A1(\systolic_inst.B_shift[17][3] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[107] ),
    .X(_02205_));
 sky130_fd_sc_hd__a22o_2 _24269_ (.A1(\systolic_inst.B_shift[17][4] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[108] ),
    .X(_02206_));
 sky130_fd_sc_hd__a22o_2 _24270_ (.A1(\systolic_inst.B_shift[17][5] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[109] ),
    .X(_02207_));
 sky130_fd_sc_hd__a22o_2 _24271_ (.A1(\systolic_inst.B_shift[17][6] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[110] ),
    .X(_02208_));
 sky130_fd_sc_hd__a22o_2 _24272_ (.A1(\systolic_inst.B_shift[17][7] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\B_in[111] ),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _24273_ (.A0(\systolic_inst.B_shift[27][0] ),
    .A1(\B_in[88] ),
    .S(_00008_),
    .X(_10610_));
 sky130_fd_sc_hd__mux2_1 _24274_ (.A0(_10610_),
    .A1(\systolic_inst.B_shift[23][0] ),
    .S(_11332_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _24275_ (.A0(\systolic_inst.B_shift[27][1] ),
    .A1(\B_in[89] ),
    .S(_00008_),
    .X(_10611_));
 sky130_fd_sc_hd__mux2_1 _24276_ (.A0(_10611_),
    .A1(\systolic_inst.B_shift[23][1] ),
    .S(_11332_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _24277_ (.A0(\systolic_inst.B_shift[27][2] ),
    .A1(\B_in[90] ),
    .S(_00008_),
    .X(_10612_));
 sky130_fd_sc_hd__mux2_1 _24278_ (.A0(_10612_),
    .A1(\systolic_inst.B_shift[23][2] ),
    .S(_11332_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _24279_ (.A0(\systolic_inst.B_shift[27][3] ),
    .A1(\B_in[91] ),
    .S(_00008_),
    .X(_10613_));
 sky130_fd_sc_hd__mux2_1 _24280_ (.A0(_10613_),
    .A1(\systolic_inst.B_shift[23][3] ),
    .S(_11332_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _24281_ (.A0(\systolic_inst.B_shift[27][4] ),
    .A1(\B_in[92] ),
    .S(_00008_),
    .X(_10614_));
 sky130_fd_sc_hd__mux2_1 _24282_ (.A0(_10614_),
    .A1(\systolic_inst.B_shift[23][4] ),
    .S(_11332_),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _24283_ (.A0(\systolic_inst.B_shift[27][5] ),
    .A1(\B_in[93] ),
    .S(_00008_),
    .X(_10615_));
 sky130_fd_sc_hd__mux2_1 _24284_ (.A0(_10615_),
    .A1(\systolic_inst.B_shift[23][5] ),
    .S(_11332_),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _24285_ (.A0(\systolic_inst.B_shift[27][6] ),
    .A1(\B_in[94] ),
    .S(_00008_),
    .X(_10616_));
 sky130_fd_sc_hd__mux2_1 _24286_ (.A0(_10616_),
    .A1(\systolic_inst.B_shift[23][6] ),
    .S(_11332_),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _24287_ (.A0(\systolic_inst.B_shift[27][7] ),
    .A1(\B_in[95] ),
    .S(_00008_),
    .X(_10617_));
 sky130_fd_sc_hd__mux2_1 _24288_ (.A0(_10617_),
    .A1(\systolic_inst.B_shift[23][7] ),
    .S(_11332_),
    .X(_02217_));
 sky130_fd_sc_hd__mux2_1 _24289_ (.A0(\systolic_inst.A_shift[12][0] ),
    .A1(\A_in[48] ),
    .S(_00008_),
    .X(_10618_));
 sky130_fd_sc_hd__mux2_1 _24290_ (.A0(_10618_),
    .A1(\systolic_inst.A_shift[11][0] ),
    .S(_11332_),
    .X(_02218_));
 sky130_fd_sc_hd__mux2_1 _24291_ (.A0(\systolic_inst.A_shift[12][1] ),
    .A1(\A_in[49] ),
    .S(_00008_),
    .X(_10619_));
 sky130_fd_sc_hd__mux2_1 _24292_ (.A0(_10619_),
    .A1(\systolic_inst.A_shift[11][1] ),
    .S(_11332_),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _24293_ (.A0(\systolic_inst.A_shift[12][2] ),
    .A1(\A_in[50] ),
    .S(_00008_),
    .X(_10620_));
 sky130_fd_sc_hd__mux2_1 _24294_ (.A0(_10620_),
    .A1(\systolic_inst.A_shift[11][2] ),
    .S(_11332_),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _24295_ (.A0(\systolic_inst.A_shift[12][3] ),
    .A1(\A_in[51] ),
    .S(_00008_),
    .X(_10621_));
 sky130_fd_sc_hd__mux2_1 _24296_ (.A0(_10621_),
    .A1(\systolic_inst.A_shift[11][3] ),
    .S(_11332_),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _24297_ (.A0(\systolic_inst.A_shift[12][4] ),
    .A1(\A_in[52] ),
    .S(_00008_),
    .X(_10622_));
 sky130_fd_sc_hd__mux2_1 _24298_ (.A0(_10622_),
    .A1(\systolic_inst.A_shift[11][4] ),
    .S(_11332_),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _24299_ (.A0(\systolic_inst.A_shift[12][5] ),
    .A1(\A_in[53] ),
    .S(_00008_),
    .X(_10623_));
 sky130_fd_sc_hd__mux2_1 _24300_ (.A0(_10623_),
    .A1(\systolic_inst.A_shift[11][5] ),
    .S(_11332_),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _24301_ (.A0(\systolic_inst.A_shift[12][6] ),
    .A1(\A_in[54] ),
    .S(_00008_),
    .X(_10624_));
 sky130_fd_sc_hd__mux2_1 _24302_ (.A0(_10624_),
    .A1(\systolic_inst.A_shift[11][6] ),
    .S(_11332_),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _24303_ (.A0(\systolic_inst.A_shift[12][7] ),
    .A1(\A_in[55] ),
    .S(_00008_),
    .X(_10625_));
 sky130_fd_sc_hd__mux2_1 _24304_ (.A0(_10625_),
    .A1(\systolic_inst.A_shift[11][7] ),
    .S(_11332_),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_1 _24305_ (.A0(\systolic_inst.A_shift[11][0] ),
    .A1(\A_in[40] ),
    .S(_00008_),
    .X(_10626_));
 sky130_fd_sc_hd__mux2_1 _24306_ (.A0(_10626_),
    .A1(\systolic_inst.A_shift[10][0] ),
    .S(_11332_),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _24307_ (.A0(\systolic_inst.A_shift[11][1] ),
    .A1(\A_in[41] ),
    .S(_00008_),
    .X(_10627_));
 sky130_fd_sc_hd__mux2_1 _24308_ (.A0(_10627_),
    .A1(\systolic_inst.A_shift[10][1] ),
    .S(_11332_),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_1 _24309_ (.A0(\systolic_inst.A_shift[11][2] ),
    .A1(\A_in[42] ),
    .S(_00008_),
    .X(_10628_));
 sky130_fd_sc_hd__mux2_1 _24310_ (.A0(_10628_),
    .A1(\systolic_inst.A_shift[10][2] ),
    .S(_11332_),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_1 _24311_ (.A0(\systolic_inst.A_shift[11][3] ),
    .A1(\A_in[43] ),
    .S(_00008_),
    .X(_10629_));
 sky130_fd_sc_hd__mux2_1 _24312_ (.A0(_10629_),
    .A1(\systolic_inst.A_shift[10][3] ),
    .S(_11332_),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _24313_ (.A0(\systolic_inst.A_shift[11][4] ),
    .A1(\A_in[44] ),
    .S(_00008_),
    .X(_10630_));
 sky130_fd_sc_hd__mux2_1 _24314_ (.A0(_10630_),
    .A1(\systolic_inst.A_shift[10][4] ),
    .S(_11332_),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _24315_ (.A0(\systolic_inst.A_shift[11][5] ),
    .A1(\A_in[45] ),
    .S(_00008_),
    .X(_10631_));
 sky130_fd_sc_hd__mux2_1 _24316_ (.A0(_10631_),
    .A1(\systolic_inst.A_shift[10][5] ),
    .S(_11332_),
    .X(_02231_));
 sky130_fd_sc_hd__mux2_1 _24317_ (.A0(\systolic_inst.A_shift[11][6] ),
    .A1(\A_in[46] ),
    .S(_00008_),
    .X(_10632_));
 sky130_fd_sc_hd__mux2_1 _24318_ (.A0(_10632_),
    .A1(\systolic_inst.A_shift[10][6] ),
    .S(_11332_),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _24319_ (.A0(\systolic_inst.A_shift[11][7] ),
    .A1(\A_in[47] ),
    .S(_00008_),
    .X(_10633_));
 sky130_fd_sc_hd__mux2_1 _24320_ (.A0(_10633_),
    .A1(\systolic_inst.A_shift[10][7] ),
    .S(_11332_),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _24321_ (.A0(\systolic_inst.A_shift[10][0] ),
    .A1(\A_in[32] ),
    .S(_00008_),
    .X(_10634_));
 sky130_fd_sc_hd__mux2_1 _24322_ (.A0(_10634_),
    .A1(\systolic_inst.A_shift[9][0] ),
    .S(_11332_),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_1 _24323_ (.A0(\systolic_inst.A_shift[10][1] ),
    .A1(\A_in[33] ),
    .S(_00008_),
    .X(_10635_));
 sky130_fd_sc_hd__mux2_1 _24324_ (.A0(_10635_),
    .A1(\systolic_inst.A_shift[9][1] ),
    .S(_11332_),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _24325_ (.A0(\systolic_inst.A_shift[10][2] ),
    .A1(\A_in[34] ),
    .S(_00008_),
    .X(_10636_));
 sky130_fd_sc_hd__mux2_1 _24326_ (.A0(_10636_),
    .A1(\systolic_inst.A_shift[9][2] ),
    .S(_11332_),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _24327_ (.A0(\systolic_inst.A_shift[10][3] ),
    .A1(\A_in[35] ),
    .S(_00008_),
    .X(_10637_));
 sky130_fd_sc_hd__mux2_1 _24328_ (.A0(_10637_),
    .A1(\systolic_inst.A_shift[9][3] ),
    .S(_11332_),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _24329_ (.A0(\systolic_inst.A_shift[10][4] ),
    .A1(\A_in[36] ),
    .S(_00008_),
    .X(_10638_));
 sky130_fd_sc_hd__mux2_1 _24330_ (.A0(_10638_),
    .A1(\systolic_inst.A_shift[9][4] ),
    .S(_11332_),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _24331_ (.A0(\systolic_inst.A_shift[10][5] ),
    .A1(\A_in[37] ),
    .S(_00008_),
    .X(_10639_));
 sky130_fd_sc_hd__mux2_1 _24332_ (.A0(_10639_),
    .A1(\systolic_inst.A_shift[9][5] ),
    .S(_11332_),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _24333_ (.A0(\systolic_inst.A_shift[10][6] ),
    .A1(\A_in[38] ),
    .S(_00008_),
    .X(_10640_));
 sky130_fd_sc_hd__mux2_1 _24334_ (.A0(_10640_),
    .A1(\systolic_inst.A_shift[9][6] ),
    .S(_11332_),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _24335_ (.A0(\systolic_inst.A_shift[10][7] ),
    .A1(\A_in[39] ),
    .S(_00008_),
    .X(_10641_));
 sky130_fd_sc_hd__mux2_1 _24336_ (.A0(_10641_),
    .A1(\systolic_inst.A_shift[9][7] ),
    .S(_11332_),
    .X(_02241_));
 sky130_fd_sc_hd__a22o_2 _24337_ (.A1(\systolic_inst.A_shift[8][0] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[9][0] ),
    .X(_02242_));
 sky130_fd_sc_hd__a22o_2 _24338_ (.A1(\systolic_inst.A_shift[8][1] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[9][1] ),
    .X(_02243_));
 sky130_fd_sc_hd__a22o_2 _24339_ (.A1(\systolic_inst.A_shift[8][2] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[9][2] ),
    .X(_02244_));
 sky130_fd_sc_hd__a22o_2 _24340_ (.A1(\systolic_inst.A_shift[8][3] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[9][3] ),
    .X(_02245_));
 sky130_fd_sc_hd__a22o_2 _24341_ (.A1(\systolic_inst.A_shift[8][4] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[9][4] ),
    .X(_02246_));
 sky130_fd_sc_hd__a22o_2 _24342_ (.A1(\systolic_inst.A_shift[8][5] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[9][5] ),
    .X(_02247_));
 sky130_fd_sc_hd__a22o_2 _24343_ (.A1(\systolic_inst.A_shift[8][6] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[9][6] ),
    .X(_02248_));
 sky130_fd_sc_hd__a22o_2 _24344_ (.A1(\systolic_inst.A_shift[8][7] ),
    .A2(_11332_),
    .B1(_10505_),
    .B2(\systolic_inst.A_shift[9][7] ),
    .X(_02249_));
 sky130_fd_sc_hd__and2_2 _24345_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[1] ),
    .X(_10642_));
 sky130_fd_sc_hd__nor2_2 _24346_ (.A(done),
    .B(C_out_frame_sync),
    .Y(_10643_));
 sky130_fd_sc_hd__a221o_2 _24347_ (.A1(\C_out[0] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[0] ),
    .C1(_10642_),
    .X(_02250_));
 sky130_fd_sc_hd__and2_2 _24348_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[2] ),
    .X(_10644_));
 sky130_fd_sc_hd__a221o_2 _24349_ (.A1(\C_out[1] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[1] ),
    .C1(_10644_),
    .X(_02251_));
 sky130_fd_sc_hd__and2_2 _24350_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[3] ),
    .X(_10645_));
 sky130_fd_sc_hd__a221o_2 _24351_ (.A1(\C_out[2] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[2] ),
    .C1(_10645_),
    .X(_02252_));
 sky130_fd_sc_hd__and2_2 _24352_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[4] ),
    .X(_10646_));
 sky130_fd_sc_hd__a221o_2 _24353_ (.A1(\C_out[3] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[3] ),
    .C1(_10646_),
    .X(_02253_));
 sky130_fd_sc_hd__and2_2 _24354_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[5] ),
    .X(_10647_));
 sky130_fd_sc_hd__a221o_2 _24355_ (.A1(\C_out[4] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[4] ),
    .C1(_10647_),
    .X(_02254_));
 sky130_fd_sc_hd__and2_2 _24356_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[6] ),
    .X(_10648_));
 sky130_fd_sc_hd__a221o_2 _24357_ (.A1(\C_out[5] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[5] ),
    .C1(_10648_),
    .X(_02255_));
 sky130_fd_sc_hd__and2_2 _24358_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[7] ),
    .X(_10649_));
 sky130_fd_sc_hd__a221o_2 _24359_ (.A1(\C_out[6] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[6] ),
    .C1(_10649_),
    .X(_02256_));
 sky130_fd_sc_hd__and2_2 _24360_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[8] ),
    .X(_10650_));
 sky130_fd_sc_hd__a221o_2 _24361_ (.A1(\C_out[7] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[7] ),
    .C1(_10650_),
    .X(_02257_));
 sky130_fd_sc_hd__and2_2 _24362_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[9] ),
    .X(_10651_));
 sky130_fd_sc_hd__a221o_2 _24363_ (.A1(\C_out[8] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[8] ),
    .C1(_10651_),
    .X(_02258_));
 sky130_fd_sc_hd__and2_2 _24364_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[10] ),
    .X(_10652_));
 sky130_fd_sc_hd__a221o_2 _24365_ (.A1(\C_out[9] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[9] ),
    .C1(_10652_),
    .X(_02259_));
 sky130_fd_sc_hd__and2_2 _24366_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[11] ),
    .X(_10653_));
 sky130_fd_sc_hd__a221o_2 _24367_ (.A1(\C_out[10] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[10] ),
    .C1(_10653_),
    .X(_02260_));
 sky130_fd_sc_hd__and2_2 _24368_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[12] ),
    .X(_10654_));
 sky130_fd_sc_hd__a221o_2 _24369_ (.A1(\C_out[11] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[11] ),
    .C1(_10654_),
    .X(_02261_));
 sky130_fd_sc_hd__and2_2 _24370_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[13] ),
    .X(_10655_));
 sky130_fd_sc_hd__a221o_2 _24371_ (.A1(\C_out[12] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[12] ),
    .C1(_10655_),
    .X(_02262_));
 sky130_fd_sc_hd__and2_2 _24372_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[14] ),
    .X(_10656_));
 sky130_fd_sc_hd__a221o_2 _24373_ (.A1(\C_out[13] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[13] ),
    .C1(_10656_),
    .X(_02263_));
 sky130_fd_sc_hd__and2_2 _24374_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[15] ),
    .X(_10657_));
 sky130_fd_sc_hd__a221o_2 _24375_ (.A1(\C_out[14] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[14] ),
    .C1(_10657_),
    .X(_02264_));
 sky130_fd_sc_hd__and2_2 _24376_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[16] ),
    .X(_10658_));
 sky130_fd_sc_hd__a221o_2 _24377_ (.A1(\C_out[15] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[15] ),
    .C1(_10658_),
    .X(_02265_));
 sky130_fd_sc_hd__and2_2 _24378_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[17] ),
    .X(_10659_));
 sky130_fd_sc_hd__a221o_2 _24379_ (.A1(\C_out[16] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[16] ),
    .C1(_10659_),
    .X(_02266_));
 sky130_fd_sc_hd__and2_2 _24380_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[18] ),
    .X(_10660_));
 sky130_fd_sc_hd__a221o_2 _24381_ (.A1(\C_out[17] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[17] ),
    .C1(_10660_),
    .X(_02267_));
 sky130_fd_sc_hd__and2_2 _24382_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[19] ),
    .X(_10661_));
 sky130_fd_sc_hd__a221o_2 _24383_ (.A1(\C_out[18] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[18] ),
    .C1(_10661_),
    .X(_02268_));
 sky130_fd_sc_hd__and2_2 _24384_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[20] ),
    .X(_10662_));
 sky130_fd_sc_hd__a221o_2 _24385_ (.A1(\C_out[19] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[19] ),
    .C1(_10662_),
    .X(_02269_));
 sky130_fd_sc_hd__and2_2 _24386_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[21] ),
    .X(_10663_));
 sky130_fd_sc_hd__a221o_2 _24387_ (.A1(\C_out[20] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[20] ),
    .C1(_10663_),
    .X(_02270_));
 sky130_fd_sc_hd__and2_2 _24388_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[22] ),
    .X(_10664_));
 sky130_fd_sc_hd__a221o_2 _24389_ (.A1(\C_out[21] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[21] ),
    .C1(_10664_),
    .X(_02271_));
 sky130_fd_sc_hd__and2_2 _24390_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[23] ),
    .X(_10665_));
 sky130_fd_sc_hd__a221o_2 _24391_ (.A1(\C_out[22] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[22] ),
    .C1(_10665_),
    .X(_02272_));
 sky130_fd_sc_hd__and2_2 _24392_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[24] ),
    .X(_10666_));
 sky130_fd_sc_hd__a221o_2 _24393_ (.A1(\C_out[23] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[23] ),
    .C1(_10666_),
    .X(_02273_));
 sky130_fd_sc_hd__and2_2 _24394_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[25] ),
    .X(_10667_));
 sky130_fd_sc_hd__a221o_2 _24395_ (.A1(\C_out[24] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[24] ),
    .C1(_10667_),
    .X(_02274_));
 sky130_fd_sc_hd__and2_2 _24396_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[26] ),
    .X(_10668_));
 sky130_fd_sc_hd__a221o_2 _24397_ (.A1(\C_out[25] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[25] ),
    .C1(_10668_),
    .X(_02275_));
 sky130_fd_sc_hd__and2_2 _24398_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[27] ),
    .X(_10669_));
 sky130_fd_sc_hd__a221o_2 _24399_ (.A1(\C_out[26] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[26] ),
    .C1(_10669_),
    .X(_02276_));
 sky130_fd_sc_hd__and2_2 _24400_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[28] ),
    .X(_10670_));
 sky130_fd_sc_hd__a221o_2 _24401_ (.A1(\C_out[27] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[27] ),
    .C1(_10670_),
    .X(_02277_));
 sky130_fd_sc_hd__and2_2 _24402_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[29] ),
    .X(_10671_));
 sky130_fd_sc_hd__a221o_2 _24403_ (.A1(\C_out[28] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[28] ),
    .C1(_10671_),
    .X(_02278_));
 sky130_fd_sc_hd__and2_2 _24404_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[30] ),
    .X(_10672_));
 sky130_fd_sc_hd__a221o_2 _24405_ (.A1(\C_out[29] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[29] ),
    .C1(_10672_),
    .X(_02279_));
 sky130_fd_sc_hd__and2_2 _24406_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[31] ),
    .X(_10673_));
 sky130_fd_sc_hd__a221o_2 _24407_ (.A1(\C_out[30] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[30] ),
    .C1(_10673_),
    .X(_02280_));
 sky130_fd_sc_hd__and2_2 _24408_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[32] ),
    .X(_10674_));
 sky130_fd_sc_hd__a221o_2 _24409_ (.A1(\C_out[31] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[31] ),
    .C1(_10674_),
    .X(_02281_));
 sky130_fd_sc_hd__and2_2 _24410_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[33] ),
    .X(_10675_));
 sky130_fd_sc_hd__a221o_2 _24411_ (.A1(\C_out[32] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[32] ),
    .C1(_10675_),
    .X(_02282_));
 sky130_fd_sc_hd__and2_2 _24412_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[34] ),
    .X(_10676_));
 sky130_fd_sc_hd__a221o_2 _24413_ (.A1(\C_out[33] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[33] ),
    .C1(_10676_),
    .X(_02283_));
 sky130_fd_sc_hd__and2_2 _24414_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[35] ),
    .X(_10677_));
 sky130_fd_sc_hd__a221o_2 _24415_ (.A1(\C_out[34] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[34] ),
    .C1(_10677_),
    .X(_02284_));
 sky130_fd_sc_hd__and2_2 _24416_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[36] ),
    .X(_10678_));
 sky130_fd_sc_hd__a221o_2 _24417_ (.A1(\C_out[35] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[35] ),
    .C1(_10678_),
    .X(_02285_));
 sky130_fd_sc_hd__and2_2 _24418_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[37] ),
    .X(_10679_));
 sky130_fd_sc_hd__a221o_2 _24419_ (.A1(\C_out[36] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[36] ),
    .C1(_10679_),
    .X(_02286_));
 sky130_fd_sc_hd__and2_2 _24420_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[38] ),
    .X(_10680_));
 sky130_fd_sc_hd__a221o_2 _24421_ (.A1(\C_out[37] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[37] ),
    .C1(_10680_),
    .X(_02287_));
 sky130_fd_sc_hd__and2_2 _24422_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[39] ),
    .X(_10681_));
 sky130_fd_sc_hd__a221o_2 _24423_ (.A1(\C_out[38] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[38] ),
    .C1(_10681_),
    .X(_02288_));
 sky130_fd_sc_hd__and2_2 _24424_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[40] ),
    .X(_10682_));
 sky130_fd_sc_hd__a221o_2 _24425_ (.A1(\C_out[39] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[39] ),
    .C1(_10682_),
    .X(_02289_));
 sky130_fd_sc_hd__and2_2 _24426_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[41] ),
    .X(_10683_));
 sky130_fd_sc_hd__a221o_2 _24427_ (.A1(\C_out[40] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[40] ),
    .C1(_10683_),
    .X(_02290_));
 sky130_fd_sc_hd__and2_2 _24428_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[42] ),
    .X(_10684_));
 sky130_fd_sc_hd__a221o_2 _24429_ (.A1(\C_out[41] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[41] ),
    .C1(_10684_),
    .X(_02291_));
 sky130_fd_sc_hd__and2_2 _24430_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[43] ),
    .X(_10685_));
 sky130_fd_sc_hd__a221o_2 _24431_ (.A1(\C_out[42] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[42] ),
    .C1(_10685_),
    .X(_02292_));
 sky130_fd_sc_hd__and2_2 _24432_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[44] ),
    .X(_10686_));
 sky130_fd_sc_hd__a221o_2 _24433_ (.A1(\C_out[43] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[43] ),
    .C1(_10686_),
    .X(_02293_));
 sky130_fd_sc_hd__and2_2 _24434_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[45] ),
    .X(_10687_));
 sky130_fd_sc_hd__a221o_2 _24435_ (.A1(\C_out[44] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[44] ),
    .C1(_10687_),
    .X(_02294_));
 sky130_fd_sc_hd__and2_2 _24436_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[46] ),
    .X(_10688_));
 sky130_fd_sc_hd__a221o_2 _24437_ (.A1(\C_out[45] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[45] ),
    .C1(_10688_),
    .X(_02295_));
 sky130_fd_sc_hd__and2_2 _24438_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[47] ),
    .X(_10689_));
 sky130_fd_sc_hd__a221o_2 _24439_ (.A1(\C_out[46] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[46] ),
    .C1(_10689_),
    .X(_02296_));
 sky130_fd_sc_hd__and2_2 _24440_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[48] ),
    .X(_10690_));
 sky130_fd_sc_hd__a221o_2 _24441_ (.A1(\C_out[47] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[47] ),
    .C1(_10690_),
    .X(_02297_));
 sky130_fd_sc_hd__and2_2 _24442_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[49] ),
    .X(_10691_));
 sky130_fd_sc_hd__a221o_2 _24443_ (.A1(\C_out[48] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[48] ),
    .C1(_10691_),
    .X(_02298_));
 sky130_fd_sc_hd__and2_2 _24444_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[50] ),
    .X(_10692_));
 sky130_fd_sc_hd__a221o_2 _24445_ (.A1(\C_out[49] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[49] ),
    .C1(_10692_),
    .X(_02299_));
 sky130_fd_sc_hd__and2_2 _24446_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[51] ),
    .X(_10693_));
 sky130_fd_sc_hd__a221o_2 _24447_ (.A1(\C_out[50] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[50] ),
    .C1(_10693_),
    .X(_02300_));
 sky130_fd_sc_hd__and2_2 _24448_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[52] ),
    .X(_10694_));
 sky130_fd_sc_hd__a221o_2 _24449_ (.A1(\C_out[51] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[51] ),
    .C1(_10694_),
    .X(_02301_));
 sky130_fd_sc_hd__and2_2 _24450_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[53] ),
    .X(_10695_));
 sky130_fd_sc_hd__a221o_2 _24451_ (.A1(\C_out[52] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[52] ),
    .C1(_10695_),
    .X(_02302_));
 sky130_fd_sc_hd__and2_2 _24452_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[54] ),
    .X(_10696_));
 sky130_fd_sc_hd__a221o_2 _24453_ (.A1(\C_out[53] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[53] ),
    .C1(_10696_),
    .X(_02303_));
 sky130_fd_sc_hd__and2_2 _24454_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[55] ),
    .X(_10697_));
 sky130_fd_sc_hd__a221o_2 _24455_ (.A1(\C_out[54] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[54] ),
    .C1(_10697_),
    .X(_02304_));
 sky130_fd_sc_hd__and2_2 _24456_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[56] ),
    .X(_10698_));
 sky130_fd_sc_hd__a221o_2 _24457_ (.A1(\C_out[55] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[55] ),
    .C1(_10698_),
    .X(_02305_));
 sky130_fd_sc_hd__and2_2 _24458_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[57] ),
    .X(_10699_));
 sky130_fd_sc_hd__a221o_2 _24459_ (.A1(\C_out[56] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[56] ),
    .C1(_10699_),
    .X(_02306_));
 sky130_fd_sc_hd__and2_2 _24460_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[58] ),
    .X(_10700_));
 sky130_fd_sc_hd__a221o_2 _24461_ (.A1(\C_out[57] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[57] ),
    .C1(_10700_),
    .X(_02307_));
 sky130_fd_sc_hd__and2_2 _24462_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[59] ),
    .X(_10701_));
 sky130_fd_sc_hd__a221o_2 _24463_ (.A1(\C_out[58] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[58] ),
    .C1(_10701_),
    .X(_02308_));
 sky130_fd_sc_hd__and2_2 _24464_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[60] ),
    .X(_10702_));
 sky130_fd_sc_hd__a221o_2 _24465_ (.A1(\C_out[59] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[59] ),
    .C1(_10702_),
    .X(_02309_));
 sky130_fd_sc_hd__and2_2 _24466_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[61] ),
    .X(_10703_));
 sky130_fd_sc_hd__a221o_2 _24467_ (.A1(\C_out[60] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[60] ),
    .C1(_10703_),
    .X(_02310_));
 sky130_fd_sc_hd__and2_2 _24468_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[62] ),
    .X(_10704_));
 sky130_fd_sc_hd__a221o_2 _24469_ (.A1(\C_out[61] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[61] ),
    .C1(_10704_),
    .X(_02311_));
 sky130_fd_sc_hd__and2_2 _24470_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[63] ),
    .X(_10705_));
 sky130_fd_sc_hd__a221o_2 _24471_ (.A1(\C_out[62] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[62] ),
    .C1(_10705_),
    .X(_02312_));
 sky130_fd_sc_hd__and2_2 _24472_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[64] ),
    .X(_10706_));
 sky130_fd_sc_hd__a221o_2 _24473_ (.A1(\C_out[63] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[63] ),
    .C1(_10706_),
    .X(_02313_));
 sky130_fd_sc_hd__and2_2 _24474_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[65] ),
    .X(_10707_));
 sky130_fd_sc_hd__a221o_2 _24475_ (.A1(\C_out[64] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[64] ),
    .C1(_10707_),
    .X(_02314_));
 sky130_fd_sc_hd__and2_2 _24476_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[66] ),
    .X(_10708_));
 sky130_fd_sc_hd__a221o_2 _24477_ (.A1(\C_out[65] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[65] ),
    .C1(_10708_),
    .X(_02315_));
 sky130_fd_sc_hd__and2_2 _24478_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[67] ),
    .X(_10709_));
 sky130_fd_sc_hd__a221o_2 _24479_ (.A1(\C_out[66] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[66] ),
    .C1(_10709_),
    .X(_02316_));
 sky130_fd_sc_hd__and2_2 _24480_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[68] ),
    .X(_10710_));
 sky130_fd_sc_hd__a221o_2 _24481_ (.A1(\C_out[67] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[67] ),
    .C1(_10710_),
    .X(_02317_));
 sky130_fd_sc_hd__and2_2 _24482_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[69] ),
    .X(_10711_));
 sky130_fd_sc_hd__a221o_2 _24483_ (.A1(\C_out[68] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[68] ),
    .C1(_10711_),
    .X(_02318_));
 sky130_fd_sc_hd__and2_2 _24484_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[70] ),
    .X(_10712_));
 sky130_fd_sc_hd__a221o_2 _24485_ (.A1(\C_out[69] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[69] ),
    .C1(_10712_),
    .X(_02319_));
 sky130_fd_sc_hd__and2_2 _24486_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[71] ),
    .X(_10713_));
 sky130_fd_sc_hd__a221o_2 _24487_ (.A1(\C_out[70] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[70] ),
    .C1(_10713_),
    .X(_02320_));
 sky130_fd_sc_hd__and2_2 _24488_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[72] ),
    .X(_10714_));
 sky130_fd_sc_hd__a221o_2 _24489_ (.A1(\C_out[71] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[71] ),
    .C1(_10714_),
    .X(_02321_));
 sky130_fd_sc_hd__and2_2 _24490_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[73] ),
    .X(_10715_));
 sky130_fd_sc_hd__a221o_2 _24491_ (.A1(\C_out[72] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[72] ),
    .C1(_10715_),
    .X(_02322_));
 sky130_fd_sc_hd__and2_2 _24492_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[74] ),
    .X(_10716_));
 sky130_fd_sc_hd__a221o_2 _24493_ (.A1(\C_out[73] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[73] ),
    .C1(_10716_),
    .X(_02323_));
 sky130_fd_sc_hd__and2_2 _24494_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[75] ),
    .X(_10717_));
 sky130_fd_sc_hd__a221o_2 _24495_ (.A1(\C_out[74] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[74] ),
    .C1(_10717_),
    .X(_02324_));
 sky130_fd_sc_hd__and2_2 _24496_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[76] ),
    .X(_10718_));
 sky130_fd_sc_hd__a221o_2 _24497_ (.A1(\C_out[75] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[75] ),
    .C1(_10718_),
    .X(_02325_));
 sky130_fd_sc_hd__and2_2 _24498_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[77] ),
    .X(_10719_));
 sky130_fd_sc_hd__a221o_2 _24499_ (.A1(\C_out[76] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[76] ),
    .C1(_10719_),
    .X(_02326_));
 sky130_fd_sc_hd__and2_2 _24500_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[78] ),
    .X(_10720_));
 sky130_fd_sc_hd__a221o_2 _24501_ (.A1(\C_out[77] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[77] ),
    .C1(_10720_),
    .X(_02327_));
 sky130_fd_sc_hd__and2_2 _24502_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[79] ),
    .X(_10721_));
 sky130_fd_sc_hd__a221o_2 _24503_ (.A1(\C_out[78] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[78] ),
    .C1(_10721_),
    .X(_02328_));
 sky130_fd_sc_hd__and2_2 _24504_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[80] ),
    .X(_10722_));
 sky130_fd_sc_hd__a221o_2 _24505_ (.A1(\C_out[79] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[79] ),
    .C1(_10722_),
    .X(_02329_));
 sky130_fd_sc_hd__and2_2 _24506_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[81] ),
    .X(_10723_));
 sky130_fd_sc_hd__a221o_2 _24507_ (.A1(\C_out[80] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[80] ),
    .C1(_10723_),
    .X(_02330_));
 sky130_fd_sc_hd__and2_2 _24508_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[82] ),
    .X(_10724_));
 sky130_fd_sc_hd__a221o_2 _24509_ (.A1(\C_out[81] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[81] ),
    .C1(_10724_),
    .X(_02331_));
 sky130_fd_sc_hd__and2_2 _24510_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[83] ),
    .X(_10725_));
 sky130_fd_sc_hd__a221o_2 _24511_ (.A1(\C_out[82] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[82] ),
    .C1(_10725_),
    .X(_02332_));
 sky130_fd_sc_hd__and2_2 _24512_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[84] ),
    .X(_10726_));
 sky130_fd_sc_hd__a221o_2 _24513_ (.A1(\C_out[83] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[83] ),
    .C1(_10726_),
    .X(_02333_));
 sky130_fd_sc_hd__and2_2 _24514_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[85] ),
    .X(_10727_));
 sky130_fd_sc_hd__a221o_2 _24515_ (.A1(\C_out[84] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[84] ),
    .C1(_10727_),
    .X(_02334_));
 sky130_fd_sc_hd__and2_2 _24516_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[86] ),
    .X(_10728_));
 sky130_fd_sc_hd__a221o_2 _24517_ (.A1(\C_out[85] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[85] ),
    .C1(_10728_),
    .X(_02335_));
 sky130_fd_sc_hd__and2_2 _24518_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[87] ),
    .X(_10729_));
 sky130_fd_sc_hd__a221o_2 _24519_ (.A1(\C_out[86] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[86] ),
    .C1(_10729_),
    .X(_02336_));
 sky130_fd_sc_hd__and2_2 _24520_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[88] ),
    .X(_10730_));
 sky130_fd_sc_hd__a221o_2 _24521_ (.A1(\C_out[87] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[87] ),
    .C1(_10730_),
    .X(_02337_));
 sky130_fd_sc_hd__and2_2 _24522_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[89] ),
    .X(_10731_));
 sky130_fd_sc_hd__a221o_2 _24523_ (.A1(\C_out[88] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[88] ),
    .C1(_10731_),
    .X(_02338_));
 sky130_fd_sc_hd__and2_2 _24524_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[90] ),
    .X(_10732_));
 sky130_fd_sc_hd__a221o_2 _24525_ (.A1(\C_out[89] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[89] ),
    .C1(_10732_),
    .X(_02339_));
 sky130_fd_sc_hd__and2_2 _24526_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[91] ),
    .X(_10733_));
 sky130_fd_sc_hd__a221o_2 _24527_ (.A1(\C_out[90] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[90] ),
    .C1(_10733_),
    .X(_02340_));
 sky130_fd_sc_hd__and2_2 _24528_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[92] ),
    .X(_10734_));
 sky130_fd_sc_hd__a221o_2 _24529_ (.A1(\C_out[91] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[91] ),
    .C1(_10734_),
    .X(_02341_));
 sky130_fd_sc_hd__and2_2 _24530_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[93] ),
    .X(_10735_));
 sky130_fd_sc_hd__a221o_2 _24531_ (.A1(\C_out[92] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[92] ),
    .C1(_10735_),
    .X(_02342_));
 sky130_fd_sc_hd__and2_2 _24532_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[94] ),
    .X(_10736_));
 sky130_fd_sc_hd__a221o_2 _24533_ (.A1(\C_out[93] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[93] ),
    .C1(_10736_),
    .X(_02343_));
 sky130_fd_sc_hd__and2_2 _24534_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[95] ),
    .X(_10737_));
 sky130_fd_sc_hd__a221o_2 _24535_ (.A1(\C_out[94] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[94] ),
    .C1(_10737_),
    .X(_02344_));
 sky130_fd_sc_hd__and2_2 _24536_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[96] ),
    .X(_10738_));
 sky130_fd_sc_hd__a221o_2 _24537_ (.A1(\C_out[95] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[95] ),
    .C1(_10738_),
    .X(_02345_));
 sky130_fd_sc_hd__and2_2 _24538_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[97] ),
    .X(_10739_));
 sky130_fd_sc_hd__a221o_2 _24539_ (.A1(\C_out[96] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[96] ),
    .C1(_10739_),
    .X(_02346_));
 sky130_fd_sc_hd__and2_2 _24540_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[98] ),
    .X(_10740_));
 sky130_fd_sc_hd__a221o_2 _24541_ (.A1(\C_out[97] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[97] ),
    .C1(_10740_),
    .X(_02347_));
 sky130_fd_sc_hd__and2_2 _24542_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[99] ),
    .X(_10741_));
 sky130_fd_sc_hd__a221o_2 _24543_ (.A1(\C_out[98] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[98] ),
    .C1(_10741_),
    .X(_02348_));
 sky130_fd_sc_hd__and2_2 _24544_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[100] ),
    .X(_10742_));
 sky130_fd_sc_hd__a221o_2 _24545_ (.A1(\C_out[99] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[99] ),
    .C1(_10742_),
    .X(_02349_));
 sky130_fd_sc_hd__and2_2 _24546_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[101] ),
    .X(_10743_));
 sky130_fd_sc_hd__a221o_2 _24547_ (.A1(\C_out[100] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[100] ),
    .C1(_10743_),
    .X(_02350_));
 sky130_fd_sc_hd__and2_2 _24548_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[102] ),
    .X(_10744_));
 sky130_fd_sc_hd__a221o_2 _24549_ (.A1(\C_out[101] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[101] ),
    .C1(_10744_),
    .X(_02351_));
 sky130_fd_sc_hd__and2_2 _24550_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[103] ),
    .X(_10745_));
 sky130_fd_sc_hd__a221o_2 _24551_ (.A1(\C_out[102] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[102] ),
    .C1(_10745_),
    .X(_02352_));
 sky130_fd_sc_hd__and2_2 _24552_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[104] ),
    .X(_10746_));
 sky130_fd_sc_hd__a221o_2 _24553_ (.A1(\C_out[103] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[103] ),
    .C1(_10746_),
    .X(_02353_));
 sky130_fd_sc_hd__and2_2 _24554_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[105] ),
    .X(_10747_));
 sky130_fd_sc_hd__a221o_2 _24555_ (.A1(\C_out[104] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[104] ),
    .C1(_10747_),
    .X(_02354_));
 sky130_fd_sc_hd__and2_2 _24556_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[106] ),
    .X(_10748_));
 sky130_fd_sc_hd__a221o_2 _24557_ (.A1(\C_out[105] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[105] ),
    .C1(_10748_),
    .X(_02355_));
 sky130_fd_sc_hd__and2_2 _24558_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[107] ),
    .X(_10749_));
 sky130_fd_sc_hd__a221o_2 _24559_ (.A1(\C_out[106] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[106] ),
    .C1(_10749_),
    .X(_02356_));
 sky130_fd_sc_hd__and2_2 _24560_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[108] ),
    .X(_10750_));
 sky130_fd_sc_hd__a221o_2 _24561_ (.A1(\C_out[107] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[107] ),
    .C1(_10750_),
    .X(_02357_));
 sky130_fd_sc_hd__and2_2 _24562_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[109] ),
    .X(_10751_));
 sky130_fd_sc_hd__a221o_2 _24563_ (.A1(\C_out[108] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[108] ),
    .C1(_10751_),
    .X(_02358_));
 sky130_fd_sc_hd__and2_2 _24564_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[110] ),
    .X(_10752_));
 sky130_fd_sc_hd__a221o_2 _24565_ (.A1(\C_out[109] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[109] ),
    .C1(_10752_),
    .X(_02359_));
 sky130_fd_sc_hd__and2_2 _24566_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[111] ),
    .X(_10753_));
 sky130_fd_sc_hd__a221o_2 _24567_ (.A1(\C_out[110] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[110] ),
    .C1(_10753_),
    .X(_02360_));
 sky130_fd_sc_hd__and2_2 _24568_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[112] ),
    .X(_10754_));
 sky130_fd_sc_hd__a221o_2 _24569_ (.A1(\C_out[111] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[111] ),
    .C1(_10754_),
    .X(_02361_));
 sky130_fd_sc_hd__and2_2 _24570_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[113] ),
    .X(_10755_));
 sky130_fd_sc_hd__a221o_2 _24571_ (.A1(\C_out[112] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[112] ),
    .C1(_10755_),
    .X(_02362_));
 sky130_fd_sc_hd__and2_2 _24572_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[114] ),
    .X(_10756_));
 sky130_fd_sc_hd__a221o_2 _24573_ (.A1(\C_out[113] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[113] ),
    .C1(_10756_),
    .X(_02363_));
 sky130_fd_sc_hd__and2_2 _24574_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[115] ),
    .X(_10757_));
 sky130_fd_sc_hd__a221o_2 _24575_ (.A1(\C_out[114] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[114] ),
    .C1(_10757_),
    .X(_02364_));
 sky130_fd_sc_hd__and2_2 _24576_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[116] ),
    .X(_10758_));
 sky130_fd_sc_hd__a221o_2 _24577_ (.A1(\C_out[115] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[115] ),
    .C1(_10758_),
    .X(_02365_));
 sky130_fd_sc_hd__and2_2 _24578_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[117] ),
    .X(_10759_));
 sky130_fd_sc_hd__a221o_2 _24579_ (.A1(\C_out[116] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[116] ),
    .C1(_10759_),
    .X(_02366_));
 sky130_fd_sc_hd__and2_2 _24580_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[118] ),
    .X(_10760_));
 sky130_fd_sc_hd__a221o_2 _24581_ (.A1(\C_out[117] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[117] ),
    .C1(_10760_),
    .X(_02367_));
 sky130_fd_sc_hd__and2_2 _24582_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[119] ),
    .X(_10761_));
 sky130_fd_sc_hd__a221o_2 _24583_ (.A1(\C_out[118] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[118] ),
    .C1(_10761_),
    .X(_02368_));
 sky130_fd_sc_hd__and2_2 _24584_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[120] ),
    .X(_10762_));
 sky130_fd_sc_hd__a221o_2 _24585_ (.A1(\C_out[119] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[119] ),
    .C1(_10762_),
    .X(_02369_));
 sky130_fd_sc_hd__and2_2 _24586_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[121] ),
    .X(_10763_));
 sky130_fd_sc_hd__a221o_2 _24587_ (.A1(\C_out[120] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[120] ),
    .C1(_10763_),
    .X(_02370_));
 sky130_fd_sc_hd__and2_2 _24588_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[122] ),
    .X(_10764_));
 sky130_fd_sc_hd__a221o_2 _24589_ (.A1(\C_out[121] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[121] ),
    .C1(_10764_),
    .X(_02371_));
 sky130_fd_sc_hd__and2_2 _24590_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[123] ),
    .X(_10765_));
 sky130_fd_sc_hd__a221o_2 _24591_ (.A1(\C_out[122] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[122] ),
    .C1(_10765_),
    .X(_02372_));
 sky130_fd_sc_hd__and2_2 _24592_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[124] ),
    .X(_10766_));
 sky130_fd_sc_hd__a221o_2 _24593_ (.A1(\C_out[123] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[123] ),
    .C1(_10766_),
    .X(_02373_));
 sky130_fd_sc_hd__and2_2 _24594_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[125] ),
    .X(_10767_));
 sky130_fd_sc_hd__a221o_2 _24595_ (.A1(\C_out[124] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[124] ),
    .C1(_10767_),
    .X(_02374_));
 sky130_fd_sc_hd__and2_2 _24596_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[126] ),
    .X(_10768_));
 sky130_fd_sc_hd__a221o_2 _24597_ (.A1(\C_out[125] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[125] ),
    .C1(_10768_),
    .X(_02375_));
 sky130_fd_sc_hd__and2_2 _24598_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[127] ),
    .X(_10769_));
 sky130_fd_sc_hd__a221o_2 _24599_ (.A1(\C_out[126] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[126] ),
    .C1(_10769_),
    .X(_02376_));
 sky130_fd_sc_hd__and2_2 _24600_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[128] ),
    .X(_10770_));
 sky130_fd_sc_hd__a221o_2 _24601_ (.A1(\C_out[127] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[127] ),
    .C1(_10770_),
    .X(_02377_));
 sky130_fd_sc_hd__and2_2 _24602_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[129] ),
    .X(_10771_));
 sky130_fd_sc_hd__a221o_2 _24603_ (.A1(\C_out[128] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[128] ),
    .C1(_10771_),
    .X(_02378_));
 sky130_fd_sc_hd__and2_2 _24604_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[130] ),
    .X(_10772_));
 sky130_fd_sc_hd__a221o_2 _24605_ (.A1(\C_out[129] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[129] ),
    .C1(_10772_),
    .X(_02379_));
 sky130_fd_sc_hd__and2_2 _24606_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[131] ),
    .X(_10773_));
 sky130_fd_sc_hd__a221o_2 _24607_ (.A1(\C_out[130] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[130] ),
    .C1(_10773_),
    .X(_02380_));
 sky130_fd_sc_hd__and2_2 _24608_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[132] ),
    .X(_10774_));
 sky130_fd_sc_hd__a221o_2 _24609_ (.A1(\C_out[131] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[131] ),
    .C1(_10774_),
    .X(_02381_));
 sky130_fd_sc_hd__and2_2 _24610_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[133] ),
    .X(_10775_));
 sky130_fd_sc_hd__a221o_2 _24611_ (.A1(\C_out[132] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[132] ),
    .C1(_10775_),
    .X(_02382_));
 sky130_fd_sc_hd__and2_2 _24612_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[134] ),
    .X(_10776_));
 sky130_fd_sc_hd__a221o_2 _24613_ (.A1(\C_out[133] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[133] ),
    .C1(_10776_),
    .X(_02383_));
 sky130_fd_sc_hd__and2_2 _24614_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[135] ),
    .X(_10777_));
 sky130_fd_sc_hd__a221o_2 _24615_ (.A1(\C_out[134] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[134] ),
    .C1(_10777_),
    .X(_02384_));
 sky130_fd_sc_hd__and2_2 _24616_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[136] ),
    .X(_10778_));
 sky130_fd_sc_hd__a221o_2 _24617_ (.A1(\C_out[135] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[135] ),
    .C1(_10778_),
    .X(_02385_));
 sky130_fd_sc_hd__and2_2 _24618_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[137] ),
    .X(_10779_));
 sky130_fd_sc_hd__a221o_2 _24619_ (.A1(\C_out[136] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[136] ),
    .C1(_10779_),
    .X(_02386_));
 sky130_fd_sc_hd__and2_2 _24620_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[138] ),
    .X(_10780_));
 sky130_fd_sc_hd__a221o_2 _24621_ (.A1(\C_out[137] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[137] ),
    .C1(_10780_),
    .X(_02387_));
 sky130_fd_sc_hd__and2_2 _24622_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[139] ),
    .X(_10781_));
 sky130_fd_sc_hd__a221o_2 _24623_ (.A1(\C_out[138] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[138] ),
    .C1(_10781_),
    .X(_02388_));
 sky130_fd_sc_hd__and2_2 _24624_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[140] ),
    .X(_10782_));
 sky130_fd_sc_hd__a221o_2 _24625_ (.A1(\C_out[139] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[139] ),
    .C1(_10782_),
    .X(_02389_));
 sky130_fd_sc_hd__and2_2 _24626_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[141] ),
    .X(_10783_));
 sky130_fd_sc_hd__a221o_2 _24627_ (.A1(\C_out[140] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[140] ),
    .C1(_10783_),
    .X(_02390_));
 sky130_fd_sc_hd__and2_2 _24628_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[142] ),
    .X(_10784_));
 sky130_fd_sc_hd__a221o_2 _24629_ (.A1(\C_out[141] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[141] ),
    .C1(_10784_),
    .X(_02391_));
 sky130_fd_sc_hd__and2_2 _24630_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[143] ),
    .X(_10785_));
 sky130_fd_sc_hd__a221o_2 _24631_ (.A1(\C_out[142] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[142] ),
    .C1(_10785_),
    .X(_02392_));
 sky130_fd_sc_hd__and2_2 _24632_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[144] ),
    .X(_10786_));
 sky130_fd_sc_hd__a221o_2 _24633_ (.A1(\C_out[143] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[143] ),
    .C1(_10786_),
    .X(_02393_));
 sky130_fd_sc_hd__and2_2 _24634_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[145] ),
    .X(_10787_));
 sky130_fd_sc_hd__a221o_2 _24635_ (.A1(\C_out[144] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[144] ),
    .C1(_10787_),
    .X(_02394_));
 sky130_fd_sc_hd__and2_2 _24636_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[146] ),
    .X(_10788_));
 sky130_fd_sc_hd__a221o_2 _24637_ (.A1(\C_out[145] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[145] ),
    .C1(_10788_),
    .X(_02395_));
 sky130_fd_sc_hd__and2_2 _24638_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[147] ),
    .X(_10789_));
 sky130_fd_sc_hd__a221o_2 _24639_ (.A1(\C_out[146] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[146] ),
    .C1(_10789_),
    .X(_02396_));
 sky130_fd_sc_hd__and2_2 _24640_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[148] ),
    .X(_10790_));
 sky130_fd_sc_hd__a221o_2 _24641_ (.A1(\C_out[147] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[147] ),
    .C1(_10790_),
    .X(_02397_));
 sky130_fd_sc_hd__and2_2 _24642_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[149] ),
    .X(_10791_));
 sky130_fd_sc_hd__a221o_2 _24643_ (.A1(\C_out[148] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[148] ),
    .C1(_10791_),
    .X(_02398_));
 sky130_fd_sc_hd__and2_2 _24644_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[150] ),
    .X(_10792_));
 sky130_fd_sc_hd__a221o_2 _24645_ (.A1(\C_out[149] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[149] ),
    .C1(_10792_),
    .X(_02399_));
 sky130_fd_sc_hd__and2_2 _24646_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[151] ),
    .X(_10793_));
 sky130_fd_sc_hd__a221o_2 _24647_ (.A1(\C_out[150] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[150] ),
    .C1(_10793_),
    .X(_02400_));
 sky130_fd_sc_hd__and2_2 _24648_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[152] ),
    .X(_10794_));
 sky130_fd_sc_hd__a221o_2 _24649_ (.A1(\C_out[151] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[151] ),
    .C1(_10794_),
    .X(_02401_));
 sky130_fd_sc_hd__and2_2 _24650_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[153] ),
    .X(_10795_));
 sky130_fd_sc_hd__a221o_2 _24651_ (.A1(\C_out[152] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[152] ),
    .C1(_10795_),
    .X(_02402_));
 sky130_fd_sc_hd__and2_2 _24652_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[154] ),
    .X(_10796_));
 sky130_fd_sc_hd__a221o_2 _24653_ (.A1(\C_out[153] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[153] ),
    .C1(_10796_),
    .X(_02403_));
 sky130_fd_sc_hd__and2_2 _24654_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[155] ),
    .X(_10797_));
 sky130_fd_sc_hd__a221o_2 _24655_ (.A1(\C_out[154] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[154] ),
    .C1(_10797_),
    .X(_02404_));
 sky130_fd_sc_hd__and2_2 _24656_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[156] ),
    .X(_10798_));
 sky130_fd_sc_hd__a221o_2 _24657_ (.A1(\C_out[155] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[155] ),
    .C1(_10798_),
    .X(_02405_));
 sky130_fd_sc_hd__and2_2 _24658_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[157] ),
    .X(_10799_));
 sky130_fd_sc_hd__a221o_2 _24659_ (.A1(\C_out[156] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[156] ),
    .C1(_10799_),
    .X(_02406_));
 sky130_fd_sc_hd__and2_2 _24660_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[158] ),
    .X(_10800_));
 sky130_fd_sc_hd__a221o_2 _24661_ (.A1(\C_out[157] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[157] ),
    .C1(_10800_),
    .X(_02407_));
 sky130_fd_sc_hd__and2_2 _24662_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[159] ),
    .X(_10801_));
 sky130_fd_sc_hd__a221o_2 _24663_ (.A1(\C_out[158] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[158] ),
    .C1(_10801_),
    .X(_02408_));
 sky130_fd_sc_hd__and2_2 _24664_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[160] ),
    .X(_10802_));
 sky130_fd_sc_hd__a221o_2 _24665_ (.A1(\C_out[159] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[159] ),
    .C1(_10802_),
    .X(_02409_));
 sky130_fd_sc_hd__and2_2 _24666_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[161] ),
    .X(_10803_));
 sky130_fd_sc_hd__a221o_2 _24667_ (.A1(\C_out[160] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[160] ),
    .C1(_10803_),
    .X(_02410_));
 sky130_fd_sc_hd__and2_2 _24668_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[162] ),
    .X(_10804_));
 sky130_fd_sc_hd__a221o_2 _24669_ (.A1(\C_out[161] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[161] ),
    .C1(_10804_),
    .X(_02411_));
 sky130_fd_sc_hd__and2_2 _24670_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[163] ),
    .X(_10805_));
 sky130_fd_sc_hd__a221o_2 _24671_ (.A1(\C_out[162] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[162] ),
    .C1(_10805_),
    .X(_02412_));
 sky130_fd_sc_hd__and2_2 _24672_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[164] ),
    .X(_10806_));
 sky130_fd_sc_hd__a221o_2 _24673_ (.A1(\C_out[163] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[163] ),
    .C1(_10806_),
    .X(_02413_));
 sky130_fd_sc_hd__and2_2 _24674_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[165] ),
    .X(_10807_));
 sky130_fd_sc_hd__a221o_2 _24675_ (.A1(\C_out[164] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[164] ),
    .C1(_10807_),
    .X(_02414_));
 sky130_fd_sc_hd__and2_2 _24676_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[166] ),
    .X(_10808_));
 sky130_fd_sc_hd__a221o_2 _24677_ (.A1(\C_out[165] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[165] ),
    .C1(_10808_),
    .X(_02415_));
 sky130_fd_sc_hd__and2_2 _24678_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[167] ),
    .X(_10809_));
 sky130_fd_sc_hd__a221o_2 _24679_ (.A1(\C_out[166] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[166] ),
    .C1(_10809_),
    .X(_02416_));
 sky130_fd_sc_hd__and2_2 _24680_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[168] ),
    .X(_10810_));
 sky130_fd_sc_hd__a221o_2 _24681_ (.A1(\C_out[167] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[167] ),
    .C1(_10810_),
    .X(_02417_));
 sky130_fd_sc_hd__and2_2 _24682_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[169] ),
    .X(_10811_));
 sky130_fd_sc_hd__a221o_2 _24683_ (.A1(\C_out[168] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[168] ),
    .C1(_10811_),
    .X(_02418_));
 sky130_fd_sc_hd__and2_2 _24684_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[170] ),
    .X(_10812_));
 sky130_fd_sc_hd__a221o_2 _24685_ (.A1(\C_out[169] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[169] ),
    .C1(_10812_),
    .X(_02419_));
 sky130_fd_sc_hd__and2_2 _24686_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[171] ),
    .X(_10813_));
 sky130_fd_sc_hd__a221o_2 _24687_ (.A1(\C_out[170] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[170] ),
    .C1(_10813_),
    .X(_02420_));
 sky130_fd_sc_hd__and2_2 _24688_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[172] ),
    .X(_10814_));
 sky130_fd_sc_hd__a221o_2 _24689_ (.A1(\C_out[171] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[171] ),
    .C1(_10814_),
    .X(_02421_));
 sky130_fd_sc_hd__and2_2 _24690_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[173] ),
    .X(_10815_));
 sky130_fd_sc_hd__a221o_2 _24691_ (.A1(\C_out[172] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[172] ),
    .C1(_10815_),
    .X(_02422_));
 sky130_fd_sc_hd__and2_2 _24692_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[174] ),
    .X(_10816_));
 sky130_fd_sc_hd__a221o_2 _24693_ (.A1(\C_out[173] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[173] ),
    .C1(_10816_),
    .X(_02423_));
 sky130_fd_sc_hd__and2_2 _24694_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[175] ),
    .X(_10817_));
 sky130_fd_sc_hd__a221o_2 _24695_ (.A1(\C_out[174] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[174] ),
    .C1(_10817_),
    .X(_02424_));
 sky130_fd_sc_hd__and2_2 _24696_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[176] ),
    .X(_10818_));
 sky130_fd_sc_hd__a221o_2 _24697_ (.A1(\C_out[175] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[175] ),
    .C1(_10818_),
    .X(_02425_));
 sky130_fd_sc_hd__and2_2 _24698_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[177] ),
    .X(_10819_));
 sky130_fd_sc_hd__a221o_2 _24699_ (.A1(\C_out[176] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[176] ),
    .C1(_10819_),
    .X(_02426_));
 sky130_fd_sc_hd__and2_2 _24700_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[178] ),
    .X(_10820_));
 sky130_fd_sc_hd__a221o_2 _24701_ (.A1(\C_out[177] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[177] ),
    .C1(_10820_),
    .X(_02427_));
 sky130_fd_sc_hd__and2_2 _24702_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[179] ),
    .X(_10821_));
 sky130_fd_sc_hd__a221o_2 _24703_ (.A1(\C_out[178] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[178] ),
    .C1(_10821_),
    .X(_02428_));
 sky130_fd_sc_hd__and2_2 _24704_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[180] ),
    .X(_10822_));
 sky130_fd_sc_hd__a221o_2 _24705_ (.A1(\C_out[179] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[179] ),
    .C1(_10822_),
    .X(_02429_));
 sky130_fd_sc_hd__and2_2 _24706_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[181] ),
    .X(_10823_));
 sky130_fd_sc_hd__a221o_2 _24707_ (.A1(\C_out[180] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[180] ),
    .C1(_10823_),
    .X(_02430_));
 sky130_fd_sc_hd__and2_2 _24708_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[182] ),
    .X(_10824_));
 sky130_fd_sc_hd__a221o_2 _24709_ (.A1(\C_out[181] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[181] ),
    .C1(_10824_),
    .X(_02431_));
 sky130_fd_sc_hd__and2_2 _24710_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[183] ),
    .X(_10825_));
 sky130_fd_sc_hd__a221o_2 _24711_ (.A1(\C_out[182] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[182] ),
    .C1(_10825_),
    .X(_02432_));
 sky130_fd_sc_hd__and2_2 _24712_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[184] ),
    .X(_10826_));
 sky130_fd_sc_hd__a221o_2 _24713_ (.A1(\C_out[183] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[183] ),
    .C1(_10826_),
    .X(_02433_));
 sky130_fd_sc_hd__and2_2 _24714_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[185] ),
    .X(_10827_));
 sky130_fd_sc_hd__a221o_2 _24715_ (.A1(\C_out[184] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[184] ),
    .C1(_10827_),
    .X(_02434_));
 sky130_fd_sc_hd__and2_2 _24716_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[186] ),
    .X(_10828_));
 sky130_fd_sc_hd__a221o_2 _24717_ (.A1(\C_out[185] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[185] ),
    .C1(_10828_),
    .X(_02435_));
 sky130_fd_sc_hd__and2_2 _24718_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[187] ),
    .X(_10829_));
 sky130_fd_sc_hd__a221o_2 _24719_ (.A1(\C_out[186] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[186] ),
    .C1(_10829_),
    .X(_02436_));
 sky130_fd_sc_hd__and2_2 _24720_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[188] ),
    .X(_10830_));
 sky130_fd_sc_hd__a221o_2 _24721_ (.A1(\C_out[187] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[187] ),
    .C1(_10830_),
    .X(_02437_));
 sky130_fd_sc_hd__and2_2 _24722_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[189] ),
    .X(_10831_));
 sky130_fd_sc_hd__a221o_2 _24723_ (.A1(\C_out[188] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[188] ),
    .C1(_10831_),
    .X(_02438_));
 sky130_fd_sc_hd__and2_2 _24724_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[190] ),
    .X(_10832_));
 sky130_fd_sc_hd__a221o_2 _24725_ (.A1(\C_out[189] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[189] ),
    .C1(_10832_),
    .X(_02439_));
 sky130_fd_sc_hd__and2_2 _24726_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[191] ),
    .X(_10833_));
 sky130_fd_sc_hd__a221o_2 _24727_ (.A1(\C_out[190] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[190] ),
    .C1(_10833_),
    .X(_02440_));
 sky130_fd_sc_hd__and2_2 _24728_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[192] ),
    .X(_10834_));
 sky130_fd_sc_hd__a221o_2 _24729_ (.A1(\C_out[191] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[191] ),
    .C1(_10834_),
    .X(_02441_));
 sky130_fd_sc_hd__and2_2 _24730_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[193] ),
    .X(_10835_));
 sky130_fd_sc_hd__a221o_2 _24731_ (.A1(\C_out[192] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[192] ),
    .C1(_10835_),
    .X(_02442_));
 sky130_fd_sc_hd__and2_2 _24732_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[194] ),
    .X(_10836_));
 sky130_fd_sc_hd__a221o_2 _24733_ (.A1(\C_out[193] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[193] ),
    .C1(_10836_),
    .X(_02443_));
 sky130_fd_sc_hd__and2_2 _24734_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[195] ),
    .X(_10837_));
 sky130_fd_sc_hd__a221o_2 _24735_ (.A1(\C_out[194] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[194] ),
    .C1(_10837_),
    .X(_02444_));
 sky130_fd_sc_hd__and2_2 _24736_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[196] ),
    .X(_10838_));
 sky130_fd_sc_hd__a221o_2 _24737_ (.A1(\C_out[195] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[195] ),
    .C1(_10838_),
    .X(_02445_));
 sky130_fd_sc_hd__and2_2 _24738_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[197] ),
    .X(_10839_));
 sky130_fd_sc_hd__a221o_2 _24739_ (.A1(\C_out[196] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[196] ),
    .C1(_10839_),
    .X(_02446_));
 sky130_fd_sc_hd__and2_2 _24740_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[198] ),
    .X(_10840_));
 sky130_fd_sc_hd__a221o_2 _24741_ (.A1(\C_out[197] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[197] ),
    .C1(_10840_),
    .X(_02447_));
 sky130_fd_sc_hd__and2_2 _24742_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[199] ),
    .X(_10841_));
 sky130_fd_sc_hd__a221o_2 _24743_ (.A1(\C_out[198] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[198] ),
    .C1(_10841_),
    .X(_02448_));
 sky130_fd_sc_hd__and2_2 _24744_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[200] ),
    .X(_10842_));
 sky130_fd_sc_hd__a221o_2 _24745_ (.A1(\C_out[199] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[199] ),
    .C1(_10842_),
    .X(_02449_));
 sky130_fd_sc_hd__and2_2 _24746_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[201] ),
    .X(_10843_));
 sky130_fd_sc_hd__a221o_2 _24747_ (.A1(\C_out[200] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[200] ),
    .C1(_10843_),
    .X(_02450_));
 sky130_fd_sc_hd__and2_2 _24748_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[202] ),
    .X(_10844_));
 sky130_fd_sc_hd__a221o_2 _24749_ (.A1(\C_out[201] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[201] ),
    .C1(_10844_),
    .X(_02451_));
 sky130_fd_sc_hd__and2_2 _24750_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[203] ),
    .X(_10845_));
 sky130_fd_sc_hd__a221o_2 _24751_ (.A1(\C_out[202] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[202] ),
    .C1(_10845_),
    .X(_02452_));
 sky130_fd_sc_hd__and2_2 _24752_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[204] ),
    .X(_10846_));
 sky130_fd_sc_hd__a221o_2 _24753_ (.A1(\C_out[203] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[203] ),
    .C1(_10846_),
    .X(_02453_));
 sky130_fd_sc_hd__and2_2 _24754_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[205] ),
    .X(_10847_));
 sky130_fd_sc_hd__a221o_2 _24755_ (.A1(\C_out[204] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[204] ),
    .C1(_10847_),
    .X(_02454_));
 sky130_fd_sc_hd__and2_2 _24756_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[206] ),
    .X(_10848_));
 sky130_fd_sc_hd__a221o_2 _24757_ (.A1(\C_out[205] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[205] ),
    .C1(_10848_),
    .X(_02455_));
 sky130_fd_sc_hd__and2_2 _24758_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[207] ),
    .X(_10849_));
 sky130_fd_sc_hd__a221o_2 _24759_ (.A1(\C_out[206] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[206] ),
    .C1(_10849_),
    .X(_02456_));
 sky130_fd_sc_hd__and2_2 _24760_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[208] ),
    .X(_10850_));
 sky130_fd_sc_hd__a221o_2 _24761_ (.A1(\C_out[207] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[207] ),
    .C1(_10850_),
    .X(_02457_));
 sky130_fd_sc_hd__and2_2 _24762_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[209] ),
    .X(_10851_));
 sky130_fd_sc_hd__a221o_2 _24763_ (.A1(\C_out[208] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[208] ),
    .C1(_10851_),
    .X(_02458_));
 sky130_fd_sc_hd__and2_2 _24764_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[210] ),
    .X(_10852_));
 sky130_fd_sc_hd__a221o_2 _24765_ (.A1(\C_out[209] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[209] ),
    .C1(_10852_),
    .X(_02459_));
 sky130_fd_sc_hd__and2_2 _24766_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[211] ),
    .X(_10853_));
 sky130_fd_sc_hd__a221o_2 _24767_ (.A1(\C_out[210] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[210] ),
    .C1(_10853_),
    .X(_02460_));
 sky130_fd_sc_hd__and2_2 _24768_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[212] ),
    .X(_10854_));
 sky130_fd_sc_hd__a221o_2 _24769_ (.A1(\C_out[211] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[211] ),
    .C1(_10854_),
    .X(_02461_));
 sky130_fd_sc_hd__and2_2 _24770_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[213] ),
    .X(_10855_));
 sky130_fd_sc_hd__a221o_2 _24771_ (.A1(\C_out[212] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[212] ),
    .C1(_10855_),
    .X(_02462_));
 sky130_fd_sc_hd__and2_2 _24772_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[214] ),
    .X(_10856_));
 sky130_fd_sc_hd__a221o_2 _24773_ (.A1(\C_out[213] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[213] ),
    .C1(_10856_),
    .X(_02463_));
 sky130_fd_sc_hd__and2_2 _24774_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[215] ),
    .X(_10857_));
 sky130_fd_sc_hd__a221o_2 _24775_ (.A1(\C_out[214] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[214] ),
    .C1(_10857_),
    .X(_02464_));
 sky130_fd_sc_hd__and2_2 _24776_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[216] ),
    .X(_10858_));
 sky130_fd_sc_hd__a221o_2 _24777_ (.A1(\C_out[215] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[215] ),
    .C1(_10858_),
    .X(_02465_));
 sky130_fd_sc_hd__and2_2 _24778_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[217] ),
    .X(_10859_));
 sky130_fd_sc_hd__a221o_2 _24779_ (.A1(\C_out[216] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[216] ),
    .C1(_10859_),
    .X(_02466_));
 sky130_fd_sc_hd__and2_2 _24780_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[218] ),
    .X(_10860_));
 sky130_fd_sc_hd__a221o_2 _24781_ (.A1(\C_out[217] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[217] ),
    .C1(_10860_),
    .X(_02467_));
 sky130_fd_sc_hd__and2_2 _24782_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[219] ),
    .X(_10861_));
 sky130_fd_sc_hd__a221o_2 _24783_ (.A1(\C_out[218] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[218] ),
    .C1(_10861_),
    .X(_02468_));
 sky130_fd_sc_hd__and2_2 _24784_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[220] ),
    .X(_10862_));
 sky130_fd_sc_hd__a221o_2 _24785_ (.A1(\C_out[219] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[219] ),
    .C1(_10862_),
    .X(_02469_));
 sky130_fd_sc_hd__and2_2 _24786_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[221] ),
    .X(_10863_));
 sky130_fd_sc_hd__a221o_2 _24787_ (.A1(\C_out[220] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[220] ),
    .C1(_10863_),
    .X(_02470_));
 sky130_fd_sc_hd__and2_2 _24788_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[222] ),
    .X(_10864_));
 sky130_fd_sc_hd__a221o_2 _24789_ (.A1(\C_out[221] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[221] ),
    .C1(_10864_),
    .X(_02471_));
 sky130_fd_sc_hd__and2_2 _24790_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[223] ),
    .X(_10865_));
 sky130_fd_sc_hd__a221o_2 _24791_ (.A1(\C_out[222] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[222] ),
    .C1(_10865_),
    .X(_02472_));
 sky130_fd_sc_hd__and2_2 _24792_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[224] ),
    .X(_10866_));
 sky130_fd_sc_hd__a221o_2 _24793_ (.A1(\C_out[223] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[223] ),
    .C1(_10866_),
    .X(_02473_));
 sky130_fd_sc_hd__and2_2 _24794_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[225] ),
    .X(_10867_));
 sky130_fd_sc_hd__a221o_2 _24795_ (.A1(\C_out[224] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[224] ),
    .C1(_10867_),
    .X(_02474_));
 sky130_fd_sc_hd__and2_2 _24796_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[226] ),
    .X(_10868_));
 sky130_fd_sc_hd__a221o_2 _24797_ (.A1(\C_out[225] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[225] ),
    .C1(_10868_),
    .X(_02475_));
 sky130_fd_sc_hd__and2_2 _24798_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[227] ),
    .X(_10869_));
 sky130_fd_sc_hd__a221o_2 _24799_ (.A1(\C_out[226] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[226] ),
    .C1(_10869_),
    .X(_02476_));
 sky130_fd_sc_hd__and2_2 _24800_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[228] ),
    .X(_10870_));
 sky130_fd_sc_hd__a221o_2 _24801_ (.A1(\C_out[227] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[227] ),
    .C1(_10870_),
    .X(_02477_));
 sky130_fd_sc_hd__and2_2 _24802_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[229] ),
    .X(_10871_));
 sky130_fd_sc_hd__a221o_2 _24803_ (.A1(\C_out[228] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[228] ),
    .C1(_10871_),
    .X(_02478_));
 sky130_fd_sc_hd__and2_2 _24804_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[230] ),
    .X(_10872_));
 sky130_fd_sc_hd__a221o_2 _24805_ (.A1(\C_out[229] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[229] ),
    .C1(_10872_),
    .X(_02479_));
 sky130_fd_sc_hd__and2_2 _24806_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[231] ),
    .X(_10873_));
 sky130_fd_sc_hd__a221o_2 _24807_ (.A1(\C_out[230] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[230] ),
    .C1(_10873_),
    .X(_02480_));
 sky130_fd_sc_hd__and2_2 _24808_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[232] ),
    .X(_10874_));
 sky130_fd_sc_hd__a221o_2 _24809_ (.A1(\C_out[231] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[231] ),
    .C1(_10874_),
    .X(_02481_));
 sky130_fd_sc_hd__and2_2 _24810_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[233] ),
    .X(_10875_));
 sky130_fd_sc_hd__a221o_2 _24811_ (.A1(\C_out[232] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[232] ),
    .C1(_10875_),
    .X(_02482_));
 sky130_fd_sc_hd__and2_2 _24812_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[234] ),
    .X(_10876_));
 sky130_fd_sc_hd__a221o_2 _24813_ (.A1(\C_out[233] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[233] ),
    .C1(_10876_),
    .X(_02483_));
 sky130_fd_sc_hd__and2_2 _24814_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[235] ),
    .X(_10877_));
 sky130_fd_sc_hd__a221o_2 _24815_ (.A1(\C_out[234] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[234] ),
    .C1(_10877_),
    .X(_02484_));
 sky130_fd_sc_hd__and2_2 _24816_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[236] ),
    .X(_10878_));
 sky130_fd_sc_hd__a221o_2 _24817_ (.A1(\C_out[235] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[235] ),
    .C1(_10878_),
    .X(_02485_));
 sky130_fd_sc_hd__and2_2 _24818_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[237] ),
    .X(_10879_));
 sky130_fd_sc_hd__a221o_2 _24819_ (.A1(\C_out[236] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[236] ),
    .C1(_10879_),
    .X(_02486_));
 sky130_fd_sc_hd__and2_2 _24820_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[238] ),
    .X(_10880_));
 sky130_fd_sc_hd__a221o_2 _24821_ (.A1(\C_out[237] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[237] ),
    .C1(_10880_),
    .X(_02487_));
 sky130_fd_sc_hd__and2_2 _24822_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[239] ),
    .X(_10881_));
 sky130_fd_sc_hd__a221o_2 _24823_ (.A1(\C_out[238] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[238] ),
    .C1(_10881_),
    .X(_02488_));
 sky130_fd_sc_hd__and2_2 _24824_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[240] ),
    .X(_10882_));
 sky130_fd_sc_hd__a221o_2 _24825_ (.A1(\C_out[239] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[239] ),
    .C1(_10882_),
    .X(_02489_));
 sky130_fd_sc_hd__and2_2 _24826_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[241] ),
    .X(_10883_));
 sky130_fd_sc_hd__a221o_2 _24827_ (.A1(\C_out[240] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[240] ),
    .C1(_10883_),
    .X(_02490_));
 sky130_fd_sc_hd__and2_2 _24828_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[242] ),
    .X(_10884_));
 sky130_fd_sc_hd__a221o_2 _24829_ (.A1(\C_out[241] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[241] ),
    .C1(_10884_),
    .X(_02491_));
 sky130_fd_sc_hd__and2_2 _24830_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[243] ),
    .X(_10885_));
 sky130_fd_sc_hd__a221o_2 _24831_ (.A1(\C_out[242] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[242] ),
    .C1(_10885_),
    .X(_02492_));
 sky130_fd_sc_hd__and2_2 _24832_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[244] ),
    .X(_10886_));
 sky130_fd_sc_hd__a221o_2 _24833_ (.A1(\C_out[243] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[243] ),
    .C1(_10886_),
    .X(_02493_));
 sky130_fd_sc_hd__and2_2 _24834_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[245] ),
    .X(_10887_));
 sky130_fd_sc_hd__a221o_2 _24835_ (.A1(\C_out[244] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[244] ),
    .C1(_10887_),
    .X(_02494_));
 sky130_fd_sc_hd__and2_2 _24836_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[246] ),
    .X(_10888_));
 sky130_fd_sc_hd__a221o_2 _24837_ (.A1(\C_out[245] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[245] ),
    .C1(_10888_),
    .X(_02495_));
 sky130_fd_sc_hd__and2_2 _24838_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[247] ),
    .X(_10889_));
 sky130_fd_sc_hd__a221o_2 _24839_ (.A1(\C_out[246] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[246] ),
    .C1(_10889_),
    .X(_02496_));
 sky130_fd_sc_hd__and2_2 _24840_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[248] ),
    .X(_10890_));
 sky130_fd_sc_hd__a221o_2 _24841_ (.A1(\C_out[247] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[247] ),
    .C1(_10890_),
    .X(_02497_));
 sky130_fd_sc_hd__and2_2 _24842_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[249] ),
    .X(_10891_));
 sky130_fd_sc_hd__a221o_2 _24843_ (.A1(\C_out[248] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[248] ),
    .C1(_10891_),
    .X(_02498_));
 sky130_fd_sc_hd__and2_2 _24844_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[250] ),
    .X(_10892_));
 sky130_fd_sc_hd__a221o_2 _24845_ (.A1(\C_out[249] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[249] ),
    .C1(_10892_),
    .X(_02499_));
 sky130_fd_sc_hd__and2_2 _24846_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[251] ),
    .X(_10893_));
 sky130_fd_sc_hd__a221o_2 _24847_ (.A1(\C_out[250] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[250] ),
    .C1(_10893_),
    .X(_02500_));
 sky130_fd_sc_hd__and2_2 _24848_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[252] ),
    .X(_10894_));
 sky130_fd_sc_hd__a221o_2 _24849_ (.A1(\C_out[251] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[251] ),
    .C1(_10894_),
    .X(_02501_));
 sky130_fd_sc_hd__and2_2 _24850_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[253] ),
    .X(_10895_));
 sky130_fd_sc_hd__a221o_2 _24851_ (.A1(\C_out[252] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[252] ),
    .C1(_10895_),
    .X(_02502_));
 sky130_fd_sc_hd__and2_2 _24852_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[254] ),
    .X(_10896_));
 sky130_fd_sc_hd__a221o_2 _24853_ (.A1(\C_out[253] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[253] ),
    .C1(_10896_),
    .X(_02503_));
 sky130_fd_sc_hd__and2_2 _24854_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[255] ),
    .X(_10897_));
 sky130_fd_sc_hd__a221o_2 _24855_ (.A1(\C_out[254] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[254] ),
    .C1(_10897_),
    .X(_02504_));
 sky130_fd_sc_hd__and2_2 _24856_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[256] ),
    .X(_10898_));
 sky130_fd_sc_hd__a221o_2 _24857_ (.A1(\C_out[255] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[255] ),
    .C1(_10898_),
    .X(_02505_));
 sky130_fd_sc_hd__and2_2 _24858_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[257] ),
    .X(_10899_));
 sky130_fd_sc_hd__a221o_2 _24859_ (.A1(\C_out[256] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[256] ),
    .C1(_10899_),
    .X(_02506_));
 sky130_fd_sc_hd__and2_2 _24860_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[258] ),
    .X(_10900_));
 sky130_fd_sc_hd__a221o_2 _24861_ (.A1(\C_out[257] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[257] ),
    .C1(_10900_),
    .X(_02507_));
 sky130_fd_sc_hd__and2_2 _24862_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[259] ),
    .X(_10901_));
 sky130_fd_sc_hd__a221o_2 _24863_ (.A1(\C_out[258] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[258] ),
    .C1(_10901_),
    .X(_02508_));
 sky130_fd_sc_hd__and2_2 _24864_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[260] ),
    .X(_10902_));
 sky130_fd_sc_hd__a221o_2 _24865_ (.A1(\C_out[259] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[259] ),
    .C1(_10902_),
    .X(_02509_));
 sky130_fd_sc_hd__and2_2 _24866_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[261] ),
    .X(_10903_));
 sky130_fd_sc_hd__a221o_2 _24867_ (.A1(\C_out[260] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[260] ),
    .C1(_10903_),
    .X(_02510_));
 sky130_fd_sc_hd__and2_2 _24868_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[262] ),
    .X(_10904_));
 sky130_fd_sc_hd__a221o_2 _24869_ (.A1(\C_out[261] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[261] ),
    .C1(_10904_),
    .X(_02511_));
 sky130_fd_sc_hd__and2_2 _24870_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[263] ),
    .X(_10905_));
 sky130_fd_sc_hd__a221o_2 _24871_ (.A1(\C_out[262] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[262] ),
    .C1(_10905_),
    .X(_02512_));
 sky130_fd_sc_hd__and2_2 _24872_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[264] ),
    .X(_10906_));
 sky130_fd_sc_hd__a221o_2 _24873_ (.A1(\C_out[263] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[263] ),
    .C1(_10906_),
    .X(_02513_));
 sky130_fd_sc_hd__and2_2 _24874_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[265] ),
    .X(_10907_));
 sky130_fd_sc_hd__a221o_2 _24875_ (.A1(\C_out[264] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[264] ),
    .C1(_10907_),
    .X(_02514_));
 sky130_fd_sc_hd__and2_2 _24876_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[266] ),
    .X(_10908_));
 sky130_fd_sc_hd__a221o_2 _24877_ (.A1(\C_out[265] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[265] ),
    .C1(_10908_),
    .X(_02515_));
 sky130_fd_sc_hd__and2_2 _24878_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[267] ),
    .X(_10909_));
 sky130_fd_sc_hd__a221o_2 _24879_ (.A1(\C_out[266] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[266] ),
    .C1(_10909_),
    .X(_02516_));
 sky130_fd_sc_hd__and2_2 _24880_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[268] ),
    .X(_10910_));
 sky130_fd_sc_hd__a221o_2 _24881_ (.A1(\C_out[267] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[267] ),
    .C1(_10910_),
    .X(_02517_));
 sky130_fd_sc_hd__and2_2 _24882_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[269] ),
    .X(_10911_));
 sky130_fd_sc_hd__a221o_2 _24883_ (.A1(\C_out[268] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[268] ),
    .C1(_10911_),
    .X(_02518_));
 sky130_fd_sc_hd__and2_2 _24884_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[270] ),
    .X(_10912_));
 sky130_fd_sc_hd__a221o_2 _24885_ (.A1(\C_out[269] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[269] ),
    .C1(_10912_),
    .X(_02519_));
 sky130_fd_sc_hd__and2_2 _24886_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[271] ),
    .X(_10913_));
 sky130_fd_sc_hd__a221o_2 _24887_ (.A1(\C_out[270] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[270] ),
    .C1(_10913_),
    .X(_02520_));
 sky130_fd_sc_hd__and2_2 _24888_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[272] ),
    .X(_10914_));
 sky130_fd_sc_hd__a221o_2 _24889_ (.A1(\C_out[271] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[271] ),
    .C1(_10914_),
    .X(_02521_));
 sky130_fd_sc_hd__and2_2 _24890_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[273] ),
    .X(_10915_));
 sky130_fd_sc_hd__a221o_2 _24891_ (.A1(\C_out[272] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[272] ),
    .C1(_10915_),
    .X(_02522_));
 sky130_fd_sc_hd__and2_2 _24892_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[274] ),
    .X(_10916_));
 sky130_fd_sc_hd__a221o_2 _24893_ (.A1(\C_out[273] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[273] ),
    .C1(_10916_),
    .X(_02523_));
 sky130_fd_sc_hd__and2_2 _24894_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[275] ),
    .X(_10917_));
 sky130_fd_sc_hd__a221o_2 _24895_ (.A1(\C_out[274] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[274] ),
    .C1(_10917_),
    .X(_02524_));
 sky130_fd_sc_hd__and2_2 _24896_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[276] ),
    .X(_10918_));
 sky130_fd_sc_hd__a221o_2 _24897_ (.A1(\C_out[275] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[275] ),
    .C1(_10918_),
    .X(_02525_));
 sky130_fd_sc_hd__and2_2 _24898_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[277] ),
    .X(_10919_));
 sky130_fd_sc_hd__a221o_2 _24899_ (.A1(\C_out[276] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[276] ),
    .C1(_10919_),
    .X(_02526_));
 sky130_fd_sc_hd__and2_2 _24900_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[278] ),
    .X(_10920_));
 sky130_fd_sc_hd__a221o_2 _24901_ (.A1(\C_out[277] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[277] ),
    .C1(_10920_),
    .X(_02527_));
 sky130_fd_sc_hd__and2_2 _24902_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[279] ),
    .X(_10921_));
 sky130_fd_sc_hd__a221o_2 _24903_ (.A1(\C_out[278] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[278] ),
    .C1(_10921_),
    .X(_02528_));
 sky130_fd_sc_hd__and2_2 _24904_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[280] ),
    .X(_10922_));
 sky130_fd_sc_hd__a221o_2 _24905_ (.A1(\C_out[279] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[279] ),
    .C1(_10922_),
    .X(_02529_));
 sky130_fd_sc_hd__and2_2 _24906_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[281] ),
    .X(_10923_));
 sky130_fd_sc_hd__a221o_2 _24907_ (.A1(\C_out[280] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[280] ),
    .C1(_10923_),
    .X(_02530_));
 sky130_fd_sc_hd__and2_2 _24908_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[282] ),
    .X(_10924_));
 sky130_fd_sc_hd__a221o_2 _24909_ (.A1(\C_out[281] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[281] ),
    .C1(_10924_),
    .X(_02531_));
 sky130_fd_sc_hd__and2_2 _24910_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[283] ),
    .X(_10925_));
 sky130_fd_sc_hd__a221o_2 _24911_ (.A1(\C_out[282] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[282] ),
    .C1(_10925_),
    .X(_02532_));
 sky130_fd_sc_hd__and2_2 _24912_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[284] ),
    .X(_10926_));
 sky130_fd_sc_hd__a221o_2 _24913_ (.A1(\C_out[283] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[283] ),
    .C1(_10926_),
    .X(_02533_));
 sky130_fd_sc_hd__and2_2 _24914_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[285] ),
    .X(_10927_));
 sky130_fd_sc_hd__a221o_2 _24915_ (.A1(\C_out[284] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[284] ),
    .C1(_10927_),
    .X(_02534_));
 sky130_fd_sc_hd__and2_2 _24916_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[286] ),
    .X(_10928_));
 sky130_fd_sc_hd__a221o_2 _24917_ (.A1(\C_out[285] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[285] ),
    .C1(_10928_),
    .X(_02535_));
 sky130_fd_sc_hd__and2_2 _24918_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[287] ),
    .X(_10929_));
 sky130_fd_sc_hd__a221o_2 _24919_ (.A1(\C_out[286] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[286] ),
    .C1(_10929_),
    .X(_02536_));
 sky130_fd_sc_hd__and2_2 _24920_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[288] ),
    .X(_10930_));
 sky130_fd_sc_hd__a221o_2 _24921_ (.A1(\C_out[287] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[287] ),
    .C1(_10930_),
    .X(_02537_));
 sky130_fd_sc_hd__and2_2 _24922_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[289] ),
    .X(_10931_));
 sky130_fd_sc_hd__a221o_2 _24923_ (.A1(\C_out[288] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[288] ),
    .C1(_10931_),
    .X(_02538_));
 sky130_fd_sc_hd__and2_2 _24924_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[290] ),
    .X(_10932_));
 sky130_fd_sc_hd__a221o_2 _24925_ (.A1(\C_out[289] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[289] ),
    .C1(_10932_),
    .X(_02539_));
 sky130_fd_sc_hd__and2_2 _24926_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[291] ),
    .X(_10933_));
 sky130_fd_sc_hd__a221o_2 _24927_ (.A1(\C_out[290] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[290] ),
    .C1(_10933_),
    .X(_02540_));
 sky130_fd_sc_hd__and2_2 _24928_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[292] ),
    .X(_10934_));
 sky130_fd_sc_hd__a221o_2 _24929_ (.A1(\C_out[291] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[291] ),
    .C1(_10934_),
    .X(_02541_));
 sky130_fd_sc_hd__and2_2 _24930_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[293] ),
    .X(_10935_));
 sky130_fd_sc_hd__a221o_2 _24931_ (.A1(\C_out[292] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[292] ),
    .C1(_10935_),
    .X(_02542_));
 sky130_fd_sc_hd__and2_2 _24932_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[294] ),
    .X(_10936_));
 sky130_fd_sc_hd__a221o_2 _24933_ (.A1(\C_out[293] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[293] ),
    .C1(_10936_),
    .X(_02543_));
 sky130_fd_sc_hd__and2_2 _24934_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[295] ),
    .X(_10937_));
 sky130_fd_sc_hd__a221o_2 _24935_ (.A1(\C_out[294] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[294] ),
    .C1(_10937_),
    .X(_02544_));
 sky130_fd_sc_hd__and2_2 _24936_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[296] ),
    .X(_10938_));
 sky130_fd_sc_hd__a221o_2 _24937_ (.A1(\C_out[295] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[295] ),
    .C1(_10938_),
    .X(_02545_));
 sky130_fd_sc_hd__and2_2 _24938_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[297] ),
    .X(_10939_));
 sky130_fd_sc_hd__a221o_2 _24939_ (.A1(\C_out[296] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[296] ),
    .C1(_10939_),
    .X(_02546_));
 sky130_fd_sc_hd__and2_2 _24940_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[298] ),
    .X(_10940_));
 sky130_fd_sc_hd__a221o_2 _24941_ (.A1(\C_out[297] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[297] ),
    .C1(_10940_),
    .X(_02547_));
 sky130_fd_sc_hd__and2_2 _24942_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[299] ),
    .X(_10941_));
 sky130_fd_sc_hd__a221o_2 _24943_ (.A1(\C_out[298] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[298] ),
    .C1(_10941_),
    .X(_02548_));
 sky130_fd_sc_hd__and2_2 _24944_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[300] ),
    .X(_10942_));
 sky130_fd_sc_hd__a221o_2 _24945_ (.A1(\C_out[299] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[299] ),
    .C1(_10942_),
    .X(_02549_));
 sky130_fd_sc_hd__and2_2 _24946_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[301] ),
    .X(_10943_));
 sky130_fd_sc_hd__a221o_2 _24947_ (.A1(\C_out[300] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[300] ),
    .C1(_10943_),
    .X(_02550_));
 sky130_fd_sc_hd__and2_2 _24948_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[302] ),
    .X(_10944_));
 sky130_fd_sc_hd__a221o_2 _24949_ (.A1(\C_out[301] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[301] ),
    .C1(_10944_),
    .X(_02551_));
 sky130_fd_sc_hd__and2_2 _24950_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[303] ),
    .X(_10945_));
 sky130_fd_sc_hd__a221o_2 _24951_ (.A1(\C_out[302] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[302] ),
    .C1(_10945_),
    .X(_02552_));
 sky130_fd_sc_hd__and2_2 _24952_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[304] ),
    .X(_10946_));
 sky130_fd_sc_hd__a221o_2 _24953_ (.A1(\C_out[303] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[303] ),
    .C1(_10946_),
    .X(_02553_));
 sky130_fd_sc_hd__and2_2 _24954_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[305] ),
    .X(_10947_));
 sky130_fd_sc_hd__a221o_2 _24955_ (.A1(\C_out[304] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[304] ),
    .C1(_10947_),
    .X(_02554_));
 sky130_fd_sc_hd__and2_2 _24956_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[306] ),
    .X(_10948_));
 sky130_fd_sc_hd__a221o_2 _24957_ (.A1(\C_out[305] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[305] ),
    .C1(_10948_),
    .X(_02555_));
 sky130_fd_sc_hd__and2_2 _24958_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[307] ),
    .X(_10949_));
 sky130_fd_sc_hd__a221o_2 _24959_ (.A1(\C_out[306] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[306] ),
    .C1(_10949_),
    .X(_02556_));
 sky130_fd_sc_hd__and2_2 _24960_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[308] ),
    .X(_10950_));
 sky130_fd_sc_hd__a221o_2 _24961_ (.A1(\C_out[307] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[307] ),
    .C1(_10950_),
    .X(_02557_));
 sky130_fd_sc_hd__and2_2 _24962_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[309] ),
    .X(_10951_));
 sky130_fd_sc_hd__a221o_2 _24963_ (.A1(\C_out[308] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[308] ),
    .C1(_10951_),
    .X(_02558_));
 sky130_fd_sc_hd__and2_2 _24964_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[310] ),
    .X(_10952_));
 sky130_fd_sc_hd__a221o_2 _24965_ (.A1(\C_out[309] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[309] ),
    .C1(_10952_),
    .X(_02559_));
 sky130_fd_sc_hd__and2_2 _24966_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[311] ),
    .X(_10953_));
 sky130_fd_sc_hd__a221o_2 _24967_ (.A1(\C_out[310] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[310] ),
    .C1(_10953_),
    .X(_02560_));
 sky130_fd_sc_hd__and2_2 _24968_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[312] ),
    .X(_10954_));
 sky130_fd_sc_hd__a221o_2 _24969_ (.A1(\C_out[311] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[311] ),
    .C1(_10954_),
    .X(_02561_));
 sky130_fd_sc_hd__and2_2 _24970_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[313] ),
    .X(_10955_));
 sky130_fd_sc_hd__a221o_2 _24971_ (.A1(\C_out[312] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[312] ),
    .C1(_10955_),
    .X(_02562_));
 sky130_fd_sc_hd__and2_2 _24972_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[314] ),
    .X(_10956_));
 sky130_fd_sc_hd__a221o_2 _24973_ (.A1(\C_out[313] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[313] ),
    .C1(_10956_),
    .X(_02563_));
 sky130_fd_sc_hd__and2_2 _24974_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[315] ),
    .X(_10957_));
 sky130_fd_sc_hd__a221o_2 _24975_ (.A1(\C_out[314] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[314] ),
    .C1(_10957_),
    .X(_02564_));
 sky130_fd_sc_hd__and2_2 _24976_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[316] ),
    .X(_10958_));
 sky130_fd_sc_hd__a221o_2 _24977_ (.A1(\C_out[315] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[315] ),
    .C1(_10958_),
    .X(_02565_));
 sky130_fd_sc_hd__and2_2 _24978_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[317] ),
    .X(_10959_));
 sky130_fd_sc_hd__a221o_2 _24979_ (.A1(\C_out[316] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[316] ),
    .C1(_10959_),
    .X(_02566_));
 sky130_fd_sc_hd__and2_2 _24980_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[318] ),
    .X(_10960_));
 sky130_fd_sc_hd__a221o_2 _24981_ (.A1(\C_out[317] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[317] ),
    .C1(_10960_),
    .X(_02567_));
 sky130_fd_sc_hd__and2_2 _24982_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[319] ),
    .X(_10961_));
 sky130_fd_sc_hd__a221o_2 _24983_ (.A1(\C_out[318] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[318] ),
    .C1(_10961_),
    .X(_02568_));
 sky130_fd_sc_hd__and2_2 _24984_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[320] ),
    .X(_10962_));
 sky130_fd_sc_hd__a221o_2 _24985_ (.A1(\C_out[319] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[319] ),
    .C1(_10962_),
    .X(_02569_));
 sky130_fd_sc_hd__and2_2 _24986_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[321] ),
    .X(_10963_));
 sky130_fd_sc_hd__a221o_2 _24987_ (.A1(\C_out[320] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[320] ),
    .C1(_10963_),
    .X(_02570_));
 sky130_fd_sc_hd__and2_2 _24988_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[322] ),
    .X(_10964_));
 sky130_fd_sc_hd__a221o_2 _24989_ (.A1(\C_out[321] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[321] ),
    .C1(_10964_),
    .X(_02571_));
 sky130_fd_sc_hd__and2_2 _24990_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[323] ),
    .X(_10965_));
 sky130_fd_sc_hd__a221o_2 _24991_ (.A1(\C_out[322] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[322] ),
    .C1(_10965_),
    .X(_02572_));
 sky130_fd_sc_hd__and2_2 _24992_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[324] ),
    .X(_10966_));
 sky130_fd_sc_hd__a221o_2 _24993_ (.A1(\C_out[323] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[323] ),
    .C1(_10966_),
    .X(_02573_));
 sky130_fd_sc_hd__and2_2 _24994_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[325] ),
    .X(_10967_));
 sky130_fd_sc_hd__a221o_2 _24995_ (.A1(\C_out[324] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[324] ),
    .C1(_10967_),
    .X(_02574_));
 sky130_fd_sc_hd__and2_2 _24996_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[326] ),
    .X(_10968_));
 sky130_fd_sc_hd__a221o_2 _24997_ (.A1(\C_out[325] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[325] ),
    .C1(_10968_),
    .X(_02575_));
 sky130_fd_sc_hd__and2_2 _24998_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[327] ),
    .X(_10969_));
 sky130_fd_sc_hd__a221o_2 _24999_ (.A1(\C_out[326] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[326] ),
    .C1(_10969_),
    .X(_02576_));
 sky130_fd_sc_hd__and2_2 _25000_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[328] ),
    .X(_10970_));
 sky130_fd_sc_hd__a221o_2 _25001_ (.A1(\C_out[327] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[327] ),
    .C1(_10970_),
    .X(_02577_));
 sky130_fd_sc_hd__and2_2 _25002_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[329] ),
    .X(_10971_));
 sky130_fd_sc_hd__a221o_2 _25003_ (.A1(\C_out[328] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[328] ),
    .C1(_10971_),
    .X(_02578_));
 sky130_fd_sc_hd__and2_2 _25004_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[330] ),
    .X(_10972_));
 sky130_fd_sc_hd__a221o_2 _25005_ (.A1(\C_out[329] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[329] ),
    .C1(_10972_),
    .X(_02579_));
 sky130_fd_sc_hd__and2_2 _25006_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[331] ),
    .X(_10973_));
 sky130_fd_sc_hd__a221o_2 _25007_ (.A1(\C_out[330] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[330] ),
    .C1(_10973_),
    .X(_02580_));
 sky130_fd_sc_hd__and2_2 _25008_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[332] ),
    .X(_10974_));
 sky130_fd_sc_hd__a221o_2 _25009_ (.A1(\C_out[331] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[331] ),
    .C1(_10974_),
    .X(_02581_));
 sky130_fd_sc_hd__and2_2 _25010_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[333] ),
    .X(_10975_));
 sky130_fd_sc_hd__a221o_2 _25011_ (.A1(\C_out[332] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[332] ),
    .C1(_10975_),
    .X(_02582_));
 sky130_fd_sc_hd__and2_2 _25012_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[334] ),
    .X(_10976_));
 sky130_fd_sc_hd__a221o_2 _25013_ (.A1(\C_out[333] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[333] ),
    .C1(_10976_),
    .X(_02583_));
 sky130_fd_sc_hd__and2_2 _25014_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[335] ),
    .X(_10977_));
 sky130_fd_sc_hd__a221o_2 _25015_ (.A1(\C_out[334] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[334] ),
    .C1(_10977_),
    .X(_02584_));
 sky130_fd_sc_hd__and2_2 _25016_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[336] ),
    .X(_10978_));
 sky130_fd_sc_hd__a221o_2 _25017_ (.A1(\C_out[335] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[335] ),
    .C1(_10978_),
    .X(_02585_));
 sky130_fd_sc_hd__and2_2 _25018_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[337] ),
    .X(_10979_));
 sky130_fd_sc_hd__a221o_2 _25019_ (.A1(\C_out[336] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[336] ),
    .C1(_10979_),
    .X(_02586_));
 sky130_fd_sc_hd__and2_2 _25020_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[338] ),
    .X(_10980_));
 sky130_fd_sc_hd__a221o_2 _25021_ (.A1(\C_out[337] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[337] ),
    .C1(_10980_),
    .X(_02587_));
 sky130_fd_sc_hd__and2_2 _25022_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[339] ),
    .X(_10981_));
 sky130_fd_sc_hd__a221o_2 _25023_ (.A1(\C_out[338] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[338] ),
    .C1(_10981_),
    .X(_02588_));
 sky130_fd_sc_hd__and2_2 _25024_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[340] ),
    .X(_10982_));
 sky130_fd_sc_hd__a221o_2 _25025_ (.A1(\C_out[339] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[339] ),
    .C1(_10982_),
    .X(_02589_));
 sky130_fd_sc_hd__and2_2 _25026_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[341] ),
    .X(_10983_));
 sky130_fd_sc_hd__a221o_2 _25027_ (.A1(\C_out[340] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[340] ),
    .C1(_10983_),
    .X(_02590_));
 sky130_fd_sc_hd__and2_2 _25028_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[342] ),
    .X(_10984_));
 sky130_fd_sc_hd__a221o_2 _25029_ (.A1(\C_out[341] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[341] ),
    .C1(_10984_),
    .X(_02591_));
 sky130_fd_sc_hd__and2_2 _25030_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[343] ),
    .X(_10985_));
 sky130_fd_sc_hd__a221o_2 _25031_ (.A1(\C_out[342] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[342] ),
    .C1(_10985_),
    .X(_02592_));
 sky130_fd_sc_hd__and2_2 _25032_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[344] ),
    .X(_10986_));
 sky130_fd_sc_hd__a221o_2 _25033_ (.A1(\C_out[343] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[343] ),
    .C1(_10986_),
    .X(_02593_));
 sky130_fd_sc_hd__and2_2 _25034_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[345] ),
    .X(_10987_));
 sky130_fd_sc_hd__a221o_2 _25035_ (.A1(\C_out[344] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[344] ),
    .C1(_10987_),
    .X(_02594_));
 sky130_fd_sc_hd__and2_2 _25036_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[346] ),
    .X(_10988_));
 sky130_fd_sc_hd__a221o_2 _25037_ (.A1(\C_out[345] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[345] ),
    .C1(_10988_),
    .X(_02595_));
 sky130_fd_sc_hd__and2_2 _25038_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[347] ),
    .X(_10989_));
 sky130_fd_sc_hd__a221o_2 _25039_ (.A1(\C_out[346] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[346] ),
    .C1(_10989_),
    .X(_02596_));
 sky130_fd_sc_hd__and2_2 _25040_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[348] ),
    .X(_10990_));
 sky130_fd_sc_hd__a221o_2 _25041_ (.A1(\C_out[347] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[347] ),
    .C1(_10990_),
    .X(_02597_));
 sky130_fd_sc_hd__and2_2 _25042_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[349] ),
    .X(_10991_));
 sky130_fd_sc_hd__a221o_2 _25043_ (.A1(\C_out[348] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[348] ),
    .C1(_10991_),
    .X(_02598_));
 sky130_fd_sc_hd__and2_2 _25044_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[350] ),
    .X(_10992_));
 sky130_fd_sc_hd__a221o_2 _25045_ (.A1(\C_out[349] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[349] ),
    .C1(_10992_),
    .X(_02599_));
 sky130_fd_sc_hd__and2_2 _25046_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[351] ),
    .X(_10993_));
 sky130_fd_sc_hd__a221o_2 _25047_ (.A1(\C_out[350] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[350] ),
    .C1(_10993_),
    .X(_02600_));
 sky130_fd_sc_hd__and2_2 _25048_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[352] ),
    .X(_10994_));
 sky130_fd_sc_hd__a221o_2 _25049_ (.A1(\C_out[351] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[351] ),
    .C1(_10994_),
    .X(_02601_));
 sky130_fd_sc_hd__and2_2 _25050_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[353] ),
    .X(_10995_));
 sky130_fd_sc_hd__a221o_2 _25051_ (.A1(\C_out[352] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[352] ),
    .C1(_10995_),
    .X(_02602_));
 sky130_fd_sc_hd__and2_2 _25052_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[354] ),
    .X(_10996_));
 sky130_fd_sc_hd__a221o_2 _25053_ (.A1(\C_out[353] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[353] ),
    .C1(_10996_),
    .X(_02603_));
 sky130_fd_sc_hd__and2_2 _25054_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[355] ),
    .X(_10997_));
 sky130_fd_sc_hd__a221o_2 _25055_ (.A1(\C_out[354] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[354] ),
    .C1(_10997_),
    .X(_02604_));
 sky130_fd_sc_hd__and2_2 _25056_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[356] ),
    .X(_10998_));
 sky130_fd_sc_hd__a221o_2 _25057_ (.A1(\C_out[355] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[355] ),
    .C1(_10998_),
    .X(_02605_));
 sky130_fd_sc_hd__and2_2 _25058_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[357] ),
    .X(_10999_));
 sky130_fd_sc_hd__a221o_2 _25059_ (.A1(\C_out[356] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[356] ),
    .C1(_10999_),
    .X(_02606_));
 sky130_fd_sc_hd__and2_2 _25060_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[358] ),
    .X(_11000_));
 sky130_fd_sc_hd__a221o_2 _25061_ (.A1(\C_out[357] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[357] ),
    .C1(_11000_),
    .X(_02607_));
 sky130_fd_sc_hd__and2_2 _25062_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[359] ),
    .X(_11001_));
 sky130_fd_sc_hd__a221o_2 _25063_ (.A1(\C_out[358] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[358] ),
    .C1(_11001_),
    .X(_02608_));
 sky130_fd_sc_hd__and2_2 _25064_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[360] ),
    .X(_11002_));
 sky130_fd_sc_hd__a221o_2 _25065_ (.A1(\C_out[359] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[359] ),
    .C1(_11002_),
    .X(_02609_));
 sky130_fd_sc_hd__and2_2 _25066_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[361] ),
    .X(_11003_));
 sky130_fd_sc_hd__a221o_2 _25067_ (.A1(\C_out[360] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[360] ),
    .C1(_11003_),
    .X(_02610_));
 sky130_fd_sc_hd__and2_2 _25068_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[362] ),
    .X(_11004_));
 sky130_fd_sc_hd__a221o_2 _25069_ (.A1(\C_out[361] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[361] ),
    .C1(_11004_),
    .X(_02611_));
 sky130_fd_sc_hd__and2_2 _25070_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[363] ),
    .X(_11005_));
 sky130_fd_sc_hd__a221o_2 _25071_ (.A1(\C_out[362] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[362] ),
    .C1(_11005_),
    .X(_02612_));
 sky130_fd_sc_hd__and2_2 _25072_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[364] ),
    .X(_11006_));
 sky130_fd_sc_hd__a221o_2 _25073_ (.A1(\C_out[363] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[363] ),
    .C1(_11006_),
    .X(_02613_));
 sky130_fd_sc_hd__and2_2 _25074_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[365] ),
    .X(_11007_));
 sky130_fd_sc_hd__a221o_2 _25075_ (.A1(\C_out[364] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[364] ),
    .C1(_11007_),
    .X(_02614_));
 sky130_fd_sc_hd__and2_2 _25076_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[366] ),
    .X(_11008_));
 sky130_fd_sc_hd__a221o_2 _25077_ (.A1(\C_out[365] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[365] ),
    .C1(_11008_),
    .X(_02615_));
 sky130_fd_sc_hd__and2_2 _25078_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[367] ),
    .X(_11009_));
 sky130_fd_sc_hd__a221o_2 _25079_ (.A1(\C_out[366] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[366] ),
    .C1(_11009_),
    .X(_02616_));
 sky130_fd_sc_hd__and2_2 _25080_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[368] ),
    .X(_11010_));
 sky130_fd_sc_hd__a221o_2 _25081_ (.A1(\C_out[367] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[367] ),
    .C1(_11010_),
    .X(_02617_));
 sky130_fd_sc_hd__and2_2 _25082_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[369] ),
    .X(_11011_));
 sky130_fd_sc_hd__a221o_2 _25083_ (.A1(\C_out[368] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[368] ),
    .C1(_11011_),
    .X(_02618_));
 sky130_fd_sc_hd__and2_2 _25084_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[370] ),
    .X(_11012_));
 sky130_fd_sc_hd__a221o_2 _25085_ (.A1(\C_out[369] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[369] ),
    .C1(_11012_),
    .X(_02619_));
 sky130_fd_sc_hd__and2_2 _25086_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[371] ),
    .X(_11013_));
 sky130_fd_sc_hd__a221o_2 _25087_ (.A1(\C_out[370] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[370] ),
    .C1(_11013_),
    .X(_02620_));
 sky130_fd_sc_hd__and2_2 _25088_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[372] ),
    .X(_11014_));
 sky130_fd_sc_hd__a221o_2 _25089_ (.A1(\C_out[371] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[371] ),
    .C1(_11014_),
    .X(_02621_));
 sky130_fd_sc_hd__and2_2 _25090_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[373] ),
    .X(_11015_));
 sky130_fd_sc_hd__a221o_2 _25091_ (.A1(\C_out[372] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[372] ),
    .C1(_11015_),
    .X(_02622_));
 sky130_fd_sc_hd__and2_2 _25092_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[374] ),
    .X(_11016_));
 sky130_fd_sc_hd__a221o_2 _25093_ (.A1(\C_out[373] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[373] ),
    .C1(_11016_),
    .X(_02623_));
 sky130_fd_sc_hd__and2_2 _25094_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[375] ),
    .X(_11017_));
 sky130_fd_sc_hd__a221o_2 _25095_ (.A1(\C_out[374] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[374] ),
    .C1(_11017_),
    .X(_02624_));
 sky130_fd_sc_hd__and2_2 _25096_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[376] ),
    .X(_11018_));
 sky130_fd_sc_hd__a221o_2 _25097_ (.A1(\C_out[375] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[375] ),
    .C1(_11018_),
    .X(_02625_));
 sky130_fd_sc_hd__and2_2 _25098_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[377] ),
    .X(_11019_));
 sky130_fd_sc_hd__a221o_2 _25099_ (.A1(\C_out[376] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[376] ),
    .C1(_11019_),
    .X(_02626_));
 sky130_fd_sc_hd__and2_2 _25100_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[378] ),
    .X(_11020_));
 sky130_fd_sc_hd__a221o_2 _25101_ (.A1(\C_out[377] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[377] ),
    .C1(_11020_),
    .X(_02627_));
 sky130_fd_sc_hd__and2_2 _25102_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[379] ),
    .X(_11021_));
 sky130_fd_sc_hd__a221o_2 _25103_ (.A1(\C_out[378] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[378] ),
    .C1(_11021_),
    .X(_02628_));
 sky130_fd_sc_hd__and2_2 _25104_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[380] ),
    .X(_11022_));
 sky130_fd_sc_hd__a221o_2 _25105_ (.A1(\C_out[379] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[379] ),
    .C1(_11022_),
    .X(_02629_));
 sky130_fd_sc_hd__and2_2 _25106_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[381] ),
    .X(_11023_));
 sky130_fd_sc_hd__a221o_2 _25107_ (.A1(\C_out[380] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[380] ),
    .C1(_11023_),
    .X(_02630_));
 sky130_fd_sc_hd__and2_2 _25108_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[382] ),
    .X(_11024_));
 sky130_fd_sc_hd__a221o_2 _25109_ (.A1(\C_out[381] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[381] ),
    .C1(_11024_),
    .X(_02631_));
 sky130_fd_sc_hd__and2_2 _25110_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[383] ),
    .X(_11025_));
 sky130_fd_sc_hd__a221o_2 _25111_ (.A1(\C_out[382] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[382] ),
    .C1(_11025_),
    .X(_02632_));
 sky130_fd_sc_hd__and2_2 _25112_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[384] ),
    .X(_11026_));
 sky130_fd_sc_hd__a221o_2 _25113_ (.A1(\C_out[383] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[383] ),
    .C1(_11026_),
    .X(_02633_));
 sky130_fd_sc_hd__and2_2 _25114_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[385] ),
    .X(_11027_));
 sky130_fd_sc_hd__a221o_2 _25115_ (.A1(\C_out[384] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[384] ),
    .C1(_11027_),
    .X(_02634_));
 sky130_fd_sc_hd__and2_2 _25116_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[386] ),
    .X(_11028_));
 sky130_fd_sc_hd__a221o_2 _25117_ (.A1(\C_out[385] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[385] ),
    .C1(_11028_),
    .X(_02635_));
 sky130_fd_sc_hd__and2_2 _25118_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[387] ),
    .X(_11029_));
 sky130_fd_sc_hd__a221o_2 _25119_ (.A1(\C_out[386] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[386] ),
    .C1(_11029_),
    .X(_02636_));
 sky130_fd_sc_hd__and2_2 _25120_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[388] ),
    .X(_11030_));
 sky130_fd_sc_hd__a221o_2 _25121_ (.A1(\C_out[387] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[387] ),
    .C1(_11030_),
    .X(_02637_));
 sky130_fd_sc_hd__and2_2 _25122_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[389] ),
    .X(_11031_));
 sky130_fd_sc_hd__a221o_2 _25123_ (.A1(\C_out[388] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[388] ),
    .C1(_11031_),
    .X(_02638_));
 sky130_fd_sc_hd__and2_2 _25124_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[390] ),
    .X(_11032_));
 sky130_fd_sc_hd__a221o_2 _25125_ (.A1(\C_out[389] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[389] ),
    .C1(_11032_),
    .X(_02639_));
 sky130_fd_sc_hd__and2_2 _25126_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[391] ),
    .X(_11033_));
 sky130_fd_sc_hd__a221o_2 _25127_ (.A1(\C_out[390] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[390] ),
    .C1(_11033_),
    .X(_02640_));
 sky130_fd_sc_hd__and2_2 _25128_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[392] ),
    .X(_11034_));
 sky130_fd_sc_hd__a221o_2 _25129_ (.A1(\C_out[391] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[391] ),
    .C1(_11034_),
    .X(_02641_));
 sky130_fd_sc_hd__and2_2 _25130_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[393] ),
    .X(_11035_));
 sky130_fd_sc_hd__a221o_2 _25131_ (.A1(\C_out[392] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[392] ),
    .C1(_11035_),
    .X(_02642_));
 sky130_fd_sc_hd__and2_2 _25132_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[394] ),
    .X(_11036_));
 sky130_fd_sc_hd__a221o_2 _25133_ (.A1(\C_out[393] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[393] ),
    .C1(_11036_),
    .X(_02643_));
 sky130_fd_sc_hd__and2_2 _25134_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[395] ),
    .X(_11037_));
 sky130_fd_sc_hd__a221o_2 _25135_ (.A1(\C_out[394] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[394] ),
    .C1(_11037_),
    .X(_02644_));
 sky130_fd_sc_hd__and2_2 _25136_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[396] ),
    .X(_11038_));
 sky130_fd_sc_hd__a221o_2 _25137_ (.A1(\C_out[395] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[395] ),
    .C1(_11038_),
    .X(_02645_));
 sky130_fd_sc_hd__and2_2 _25138_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[397] ),
    .X(_11039_));
 sky130_fd_sc_hd__a221o_2 _25139_ (.A1(\C_out[396] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[396] ),
    .C1(_11039_),
    .X(_02646_));
 sky130_fd_sc_hd__and2_2 _25140_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[398] ),
    .X(_11040_));
 sky130_fd_sc_hd__a221o_2 _25141_ (.A1(\C_out[397] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[397] ),
    .C1(_11040_),
    .X(_02647_));
 sky130_fd_sc_hd__and2_2 _25142_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[399] ),
    .X(_11041_));
 sky130_fd_sc_hd__a221o_2 _25143_ (.A1(\C_out[398] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[398] ),
    .C1(_11041_),
    .X(_02648_));
 sky130_fd_sc_hd__and2_2 _25144_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[400] ),
    .X(_11042_));
 sky130_fd_sc_hd__a221o_2 _25145_ (.A1(\C_out[399] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[399] ),
    .C1(_11042_),
    .X(_02649_));
 sky130_fd_sc_hd__and2_2 _25146_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[401] ),
    .X(_11043_));
 sky130_fd_sc_hd__a221o_2 _25147_ (.A1(\C_out[400] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[400] ),
    .C1(_11043_),
    .X(_02650_));
 sky130_fd_sc_hd__and2_2 _25148_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[402] ),
    .X(_11044_));
 sky130_fd_sc_hd__a221o_2 _25149_ (.A1(\C_out[401] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[401] ),
    .C1(_11044_),
    .X(_02651_));
 sky130_fd_sc_hd__and2_2 _25150_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[403] ),
    .X(_11045_));
 sky130_fd_sc_hd__a221o_2 _25151_ (.A1(\C_out[402] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[402] ),
    .C1(_11045_),
    .X(_02652_));
 sky130_fd_sc_hd__and2_2 _25152_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[404] ),
    .X(_11046_));
 sky130_fd_sc_hd__a221o_2 _25153_ (.A1(\C_out[403] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[403] ),
    .C1(_11046_),
    .X(_02653_));
 sky130_fd_sc_hd__and2_2 _25154_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[405] ),
    .X(_11047_));
 sky130_fd_sc_hd__a221o_2 _25155_ (.A1(\C_out[404] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[404] ),
    .C1(_11047_),
    .X(_02654_));
 sky130_fd_sc_hd__and2_2 _25156_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[406] ),
    .X(_11048_));
 sky130_fd_sc_hd__a221o_2 _25157_ (.A1(\C_out[405] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[405] ),
    .C1(_11048_),
    .X(_02655_));
 sky130_fd_sc_hd__and2_2 _25158_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[407] ),
    .X(_11049_));
 sky130_fd_sc_hd__a221o_2 _25159_ (.A1(\C_out[406] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[406] ),
    .C1(_11049_),
    .X(_02656_));
 sky130_fd_sc_hd__and2_2 _25160_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[408] ),
    .X(_11050_));
 sky130_fd_sc_hd__a221o_2 _25161_ (.A1(\C_out[407] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[407] ),
    .C1(_11050_),
    .X(_02657_));
 sky130_fd_sc_hd__and2_2 _25162_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[409] ),
    .X(_11051_));
 sky130_fd_sc_hd__a221o_2 _25163_ (.A1(\C_out[408] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[408] ),
    .C1(_11051_),
    .X(_02658_));
 sky130_fd_sc_hd__and2_2 _25164_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[410] ),
    .X(_11052_));
 sky130_fd_sc_hd__a221o_2 _25165_ (.A1(\C_out[409] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[409] ),
    .C1(_11052_),
    .X(_02659_));
 sky130_fd_sc_hd__and2_2 _25166_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[411] ),
    .X(_11053_));
 sky130_fd_sc_hd__a221o_2 _25167_ (.A1(\C_out[410] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[410] ),
    .C1(_11053_),
    .X(_02660_));
 sky130_fd_sc_hd__and2_2 _25168_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[412] ),
    .X(_11054_));
 sky130_fd_sc_hd__a221o_2 _25169_ (.A1(\C_out[411] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[411] ),
    .C1(_11054_),
    .X(_02661_));
 sky130_fd_sc_hd__and2_2 _25170_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[413] ),
    .X(_11055_));
 sky130_fd_sc_hd__a221o_2 _25171_ (.A1(\C_out[412] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[412] ),
    .C1(_11055_),
    .X(_02662_));
 sky130_fd_sc_hd__and2_2 _25172_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[414] ),
    .X(_11056_));
 sky130_fd_sc_hd__a221o_2 _25173_ (.A1(\C_out[413] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[413] ),
    .C1(_11056_),
    .X(_02663_));
 sky130_fd_sc_hd__and2_2 _25174_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[415] ),
    .X(_11057_));
 sky130_fd_sc_hd__a221o_2 _25175_ (.A1(\C_out[414] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[414] ),
    .C1(_11057_),
    .X(_02664_));
 sky130_fd_sc_hd__and2_2 _25176_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[416] ),
    .X(_11058_));
 sky130_fd_sc_hd__a221o_2 _25177_ (.A1(\C_out[415] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[415] ),
    .C1(_11058_),
    .X(_02665_));
 sky130_fd_sc_hd__and2_2 _25178_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[417] ),
    .X(_11059_));
 sky130_fd_sc_hd__a221o_2 _25179_ (.A1(\C_out[416] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[416] ),
    .C1(_11059_),
    .X(_02666_));
 sky130_fd_sc_hd__and2_2 _25180_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[418] ),
    .X(_11060_));
 sky130_fd_sc_hd__a221o_2 _25181_ (.A1(\C_out[417] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[417] ),
    .C1(_11060_),
    .X(_02667_));
 sky130_fd_sc_hd__and2_2 _25182_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[419] ),
    .X(_11061_));
 sky130_fd_sc_hd__a221o_2 _25183_ (.A1(\C_out[418] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[418] ),
    .C1(_11061_),
    .X(_02668_));
 sky130_fd_sc_hd__and2_2 _25184_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[420] ),
    .X(_11062_));
 sky130_fd_sc_hd__a221o_2 _25185_ (.A1(\C_out[419] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[419] ),
    .C1(_11062_),
    .X(_02669_));
 sky130_fd_sc_hd__and2_2 _25186_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[421] ),
    .X(_11063_));
 sky130_fd_sc_hd__a221o_2 _25187_ (.A1(\C_out[420] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[420] ),
    .C1(_11063_),
    .X(_02670_));
 sky130_fd_sc_hd__and2_2 _25188_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[422] ),
    .X(_11064_));
 sky130_fd_sc_hd__a221o_2 _25189_ (.A1(\C_out[421] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[421] ),
    .C1(_11064_),
    .X(_02671_));
 sky130_fd_sc_hd__and2_2 _25190_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[423] ),
    .X(_11065_));
 sky130_fd_sc_hd__a221o_2 _25191_ (.A1(\C_out[422] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[422] ),
    .C1(_11065_),
    .X(_02672_));
 sky130_fd_sc_hd__and2_2 _25192_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[424] ),
    .X(_11066_));
 sky130_fd_sc_hd__a221o_2 _25193_ (.A1(\C_out[423] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[423] ),
    .C1(_11066_),
    .X(_02673_));
 sky130_fd_sc_hd__and2_2 _25194_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[425] ),
    .X(_11067_));
 sky130_fd_sc_hd__a221o_2 _25195_ (.A1(\C_out[424] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[424] ),
    .C1(_11067_),
    .X(_02674_));
 sky130_fd_sc_hd__and2_2 _25196_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[426] ),
    .X(_11068_));
 sky130_fd_sc_hd__a221o_2 _25197_ (.A1(\C_out[425] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[425] ),
    .C1(_11068_),
    .X(_02675_));
 sky130_fd_sc_hd__and2_2 _25198_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[427] ),
    .X(_11069_));
 sky130_fd_sc_hd__a221o_2 _25199_ (.A1(\C_out[426] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[426] ),
    .C1(_11069_),
    .X(_02676_));
 sky130_fd_sc_hd__and2_2 _25200_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[428] ),
    .X(_11070_));
 sky130_fd_sc_hd__a221o_2 _25201_ (.A1(\C_out[427] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[427] ),
    .C1(_11070_),
    .X(_02677_));
 sky130_fd_sc_hd__and2_2 _25202_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[429] ),
    .X(_11071_));
 sky130_fd_sc_hd__a221o_2 _25203_ (.A1(\C_out[428] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[428] ),
    .C1(_11071_),
    .X(_02678_));
 sky130_fd_sc_hd__and2_2 _25204_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[430] ),
    .X(_11072_));
 sky130_fd_sc_hd__a221o_2 _25205_ (.A1(\C_out[429] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[429] ),
    .C1(_11072_),
    .X(_02679_));
 sky130_fd_sc_hd__and2_2 _25206_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[431] ),
    .X(_11073_));
 sky130_fd_sc_hd__a221o_2 _25207_ (.A1(\C_out[430] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[430] ),
    .C1(_11073_),
    .X(_02680_));
 sky130_fd_sc_hd__and2_2 _25208_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[432] ),
    .X(_11074_));
 sky130_fd_sc_hd__a221o_2 _25209_ (.A1(\C_out[431] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[431] ),
    .C1(_11074_),
    .X(_02681_));
 sky130_fd_sc_hd__and2_2 _25210_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[433] ),
    .X(_11075_));
 sky130_fd_sc_hd__a221o_2 _25211_ (.A1(\C_out[432] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[432] ),
    .C1(_11075_),
    .X(_02682_));
 sky130_fd_sc_hd__and2_2 _25212_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[434] ),
    .X(_11076_));
 sky130_fd_sc_hd__a221o_2 _25213_ (.A1(\C_out[433] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[433] ),
    .C1(_11076_),
    .X(_02683_));
 sky130_fd_sc_hd__and2_2 _25214_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[435] ),
    .X(_11077_));
 sky130_fd_sc_hd__a221o_2 _25215_ (.A1(\C_out[434] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[434] ),
    .C1(_11077_),
    .X(_02684_));
 sky130_fd_sc_hd__and2_2 _25216_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[436] ),
    .X(_11078_));
 sky130_fd_sc_hd__a221o_2 _25217_ (.A1(\C_out[435] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[435] ),
    .C1(_11078_),
    .X(_02685_));
 sky130_fd_sc_hd__and2_2 _25218_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[437] ),
    .X(_11079_));
 sky130_fd_sc_hd__a221o_2 _25219_ (.A1(\C_out[436] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[436] ),
    .C1(_11079_),
    .X(_02686_));
 sky130_fd_sc_hd__and2_2 _25220_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[438] ),
    .X(_11080_));
 sky130_fd_sc_hd__a221o_2 _25221_ (.A1(\C_out[437] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[437] ),
    .C1(_11080_),
    .X(_02687_));
 sky130_fd_sc_hd__and2_2 _25222_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[439] ),
    .X(_11081_));
 sky130_fd_sc_hd__a221o_2 _25223_ (.A1(\C_out[438] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[438] ),
    .C1(_11081_),
    .X(_02688_));
 sky130_fd_sc_hd__and2_2 _25224_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[440] ),
    .X(_11082_));
 sky130_fd_sc_hd__a221o_2 _25225_ (.A1(\C_out[439] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[439] ),
    .C1(_11082_),
    .X(_02689_));
 sky130_fd_sc_hd__and2_2 _25226_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[441] ),
    .X(_11083_));
 sky130_fd_sc_hd__a221o_2 _25227_ (.A1(\ser_C.parallel_data[440] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[440] ),
    .C1(_11083_),
    .X(_02690_));
 sky130_fd_sc_hd__and2_2 _25228_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[442] ),
    .X(_11084_));
 sky130_fd_sc_hd__a221o_2 _25229_ (.A1(\ser_C.parallel_data[441] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[441] ),
    .C1(_11084_),
    .X(_02691_));
 sky130_fd_sc_hd__and2_2 _25230_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[443] ),
    .X(_11085_));
 sky130_fd_sc_hd__a221o_2 _25231_ (.A1(\ser_C.parallel_data[442] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[442] ),
    .C1(_11085_),
    .X(_02692_));
 sky130_fd_sc_hd__and2_2 _25232_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[444] ),
    .X(_11086_));
 sky130_fd_sc_hd__a221o_2 _25233_ (.A1(\ser_C.parallel_data[443] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[443] ),
    .C1(_11086_),
    .X(_02693_));
 sky130_fd_sc_hd__and2_2 _25234_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[445] ),
    .X(_11087_));
 sky130_fd_sc_hd__a221o_2 _25235_ (.A1(\ser_C.parallel_data[444] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[444] ),
    .C1(_11087_),
    .X(_02694_));
 sky130_fd_sc_hd__and2_2 _25236_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[446] ),
    .X(_11088_));
 sky130_fd_sc_hd__a221o_2 _25237_ (.A1(\ser_C.parallel_data[445] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[445] ),
    .C1(_11088_),
    .X(_02695_));
 sky130_fd_sc_hd__and2_2 _25238_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[447] ),
    .X(_11089_));
 sky130_fd_sc_hd__a221o_2 _25239_ (.A1(\ser_C.parallel_data[446] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[446] ),
    .C1(_11089_),
    .X(_02696_));
 sky130_fd_sc_hd__and2_2 _25240_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[448] ),
    .X(_11090_));
 sky130_fd_sc_hd__a221o_2 _25241_ (.A1(\ser_C.parallel_data[447] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[447] ),
    .C1(_11090_),
    .X(_02697_));
 sky130_fd_sc_hd__and2_2 _25242_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[449] ),
    .X(_11091_));
 sky130_fd_sc_hd__a221o_2 _25243_ (.A1(\ser_C.parallel_data[448] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[448] ),
    .C1(_11091_),
    .X(_02698_));
 sky130_fd_sc_hd__and2_2 _25244_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[450] ),
    .X(_11092_));
 sky130_fd_sc_hd__a221o_2 _25245_ (.A1(\ser_C.parallel_data[449] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[449] ),
    .C1(_11092_),
    .X(_02699_));
 sky130_fd_sc_hd__and2_2 _25246_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[451] ),
    .X(_11093_));
 sky130_fd_sc_hd__a221o_2 _25247_ (.A1(\ser_C.parallel_data[450] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[450] ),
    .C1(_11093_),
    .X(_02700_));
 sky130_fd_sc_hd__and2_2 _25248_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[452] ),
    .X(_11094_));
 sky130_fd_sc_hd__a221o_2 _25249_ (.A1(\ser_C.parallel_data[451] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[451] ),
    .C1(_11094_),
    .X(_02701_));
 sky130_fd_sc_hd__and2_2 _25250_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[453] ),
    .X(_11095_));
 sky130_fd_sc_hd__a221o_2 _25251_ (.A1(\ser_C.parallel_data[452] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[452] ),
    .C1(_11095_),
    .X(_02702_));
 sky130_fd_sc_hd__and2_2 _25252_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[454] ),
    .X(_11096_));
 sky130_fd_sc_hd__a221o_2 _25253_ (.A1(\ser_C.parallel_data[453] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[453] ),
    .C1(_11096_),
    .X(_02703_));
 sky130_fd_sc_hd__and2_2 _25254_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[455] ),
    .X(_11097_));
 sky130_fd_sc_hd__a221o_2 _25255_ (.A1(\ser_C.parallel_data[454] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[454] ),
    .C1(_11097_),
    .X(_02704_));
 sky130_fd_sc_hd__and2_2 _25256_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[456] ),
    .X(_11098_));
 sky130_fd_sc_hd__a221o_2 _25257_ (.A1(\ser_C.parallel_data[455] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[455] ),
    .C1(_11098_),
    .X(_02705_));
 sky130_fd_sc_hd__and2_2 _25258_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[457] ),
    .X(_11099_));
 sky130_fd_sc_hd__a221o_2 _25259_ (.A1(\ser_C.parallel_data[456] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[456] ),
    .C1(_11099_),
    .X(_02706_));
 sky130_fd_sc_hd__and2_2 _25260_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[458] ),
    .X(_11100_));
 sky130_fd_sc_hd__a221o_2 _25261_ (.A1(\ser_C.parallel_data[457] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[457] ),
    .C1(_11100_),
    .X(_02707_));
 sky130_fd_sc_hd__and2_2 _25262_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[459] ),
    .X(_11101_));
 sky130_fd_sc_hd__a221o_2 _25263_ (.A1(\ser_C.parallel_data[458] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[458] ),
    .C1(_11101_),
    .X(_02708_));
 sky130_fd_sc_hd__and2_2 _25264_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[460] ),
    .X(_11102_));
 sky130_fd_sc_hd__a221o_2 _25265_ (.A1(\ser_C.parallel_data[459] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[459] ),
    .C1(_11102_),
    .X(_02709_));
 sky130_fd_sc_hd__and2_2 _25266_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[461] ),
    .X(_11103_));
 sky130_fd_sc_hd__a221o_2 _25267_ (.A1(\ser_C.parallel_data[460] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[460] ),
    .C1(_11103_),
    .X(_02710_));
 sky130_fd_sc_hd__and2_2 _25268_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[462] ),
    .X(_11104_));
 sky130_fd_sc_hd__a221o_2 _25269_ (.A1(\ser_C.parallel_data[461] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[461] ),
    .C1(_11104_),
    .X(_02711_));
 sky130_fd_sc_hd__and2_2 _25270_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[463] ),
    .X(_11105_));
 sky130_fd_sc_hd__a221o_2 _25271_ (.A1(\ser_C.parallel_data[462] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[462] ),
    .C1(_11105_),
    .X(_02712_));
 sky130_fd_sc_hd__and2_2 _25272_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[464] ),
    .X(_11106_));
 sky130_fd_sc_hd__a221o_2 _25273_ (.A1(\ser_C.parallel_data[463] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[463] ),
    .C1(_11106_),
    .X(_02713_));
 sky130_fd_sc_hd__and2_2 _25274_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[465] ),
    .X(_11107_));
 sky130_fd_sc_hd__a221o_2 _25275_ (.A1(\ser_C.parallel_data[464] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[464] ),
    .C1(_11107_),
    .X(_02714_));
 sky130_fd_sc_hd__and2_2 _25276_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[466] ),
    .X(_11108_));
 sky130_fd_sc_hd__a221o_2 _25277_ (.A1(\ser_C.parallel_data[465] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[465] ),
    .C1(_11108_),
    .X(_02715_));
 sky130_fd_sc_hd__and2_2 _25278_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[467] ),
    .X(_11109_));
 sky130_fd_sc_hd__a221o_2 _25279_ (.A1(\ser_C.parallel_data[466] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[466] ),
    .C1(_11109_),
    .X(_02716_));
 sky130_fd_sc_hd__and2_2 _25280_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[468] ),
    .X(_11110_));
 sky130_fd_sc_hd__a221o_2 _25281_ (.A1(\ser_C.parallel_data[467] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[467] ),
    .C1(_11110_),
    .X(_02717_));
 sky130_fd_sc_hd__and2_2 _25282_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[469] ),
    .X(_11111_));
 sky130_fd_sc_hd__a221o_2 _25283_ (.A1(\ser_C.parallel_data[468] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[468] ),
    .C1(_11111_),
    .X(_02718_));
 sky130_fd_sc_hd__and2_2 _25284_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[470] ),
    .X(_11112_));
 sky130_fd_sc_hd__a221o_2 _25285_ (.A1(\ser_C.parallel_data[469] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[469] ),
    .C1(_11112_),
    .X(_02719_));
 sky130_fd_sc_hd__and2_2 _25286_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[471] ),
    .X(_11113_));
 sky130_fd_sc_hd__a221o_2 _25287_ (.A1(\ser_C.parallel_data[470] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[470] ),
    .C1(_11113_),
    .X(_02720_));
 sky130_fd_sc_hd__and2_2 _25288_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[472] ),
    .X(_11114_));
 sky130_fd_sc_hd__a221o_2 _25289_ (.A1(\ser_C.parallel_data[471] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[471] ),
    .C1(_11114_),
    .X(_02721_));
 sky130_fd_sc_hd__and2_2 _25290_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[473] ),
    .X(_11115_));
 sky130_fd_sc_hd__a221o_2 _25291_ (.A1(\ser_C.parallel_data[472] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[472] ),
    .C1(_11115_),
    .X(_02722_));
 sky130_fd_sc_hd__and2_2 _25292_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[474] ),
    .X(_11116_));
 sky130_fd_sc_hd__a221o_2 _25293_ (.A1(\ser_C.parallel_data[473] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[473] ),
    .C1(_11116_),
    .X(_02723_));
 sky130_fd_sc_hd__and2_2 _25294_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[475] ),
    .X(_11117_));
 sky130_fd_sc_hd__a221o_2 _25295_ (.A1(\ser_C.parallel_data[474] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[474] ),
    .C1(_11117_),
    .X(_02724_));
 sky130_fd_sc_hd__and2_2 _25296_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[476] ),
    .X(_11118_));
 sky130_fd_sc_hd__a221o_2 _25297_ (.A1(\ser_C.parallel_data[475] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[475] ),
    .C1(_11118_),
    .X(_02725_));
 sky130_fd_sc_hd__and2_2 _25298_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[477] ),
    .X(_11119_));
 sky130_fd_sc_hd__a221o_2 _25299_ (.A1(\ser_C.parallel_data[476] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[476] ),
    .C1(_11119_),
    .X(_02726_));
 sky130_fd_sc_hd__and2_2 _25300_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[478] ),
    .X(_11120_));
 sky130_fd_sc_hd__a221o_2 _25301_ (.A1(\ser_C.parallel_data[477] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[477] ),
    .C1(_11120_),
    .X(_02727_));
 sky130_fd_sc_hd__and2_2 _25302_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[479] ),
    .X(_11121_));
 sky130_fd_sc_hd__a221o_2 _25303_ (.A1(\ser_C.parallel_data[478] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[478] ),
    .C1(_11121_),
    .X(_02728_));
 sky130_fd_sc_hd__and2_2 _25304_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[480] ),
    .X(_11122_));
 sky130_fd_sc_hd__a221o_2 _25305_ (.A1(\ser_C.parallel_data[479] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[479] ),
    .C1(_11122_),
    .X(_02729_));
 sky130_fd_sc_hd__and2_2 _25306_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[481] ),
    .X(_11123_));
 sky130_fd_sc_hd__a221o_2 _25307_ (.A1(\ser_C.parallel_data[480] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[480] ),
    .C1(_11123_),
    .X(_02730_));
 sky130_fd_sc_hd__and2_2 _25308_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[482] ),
    .X(_11124_));
 sky130_fd_sc_hd__a221o_2 _25309_ (.A1(\ser_C.parallel_data[481] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[481] ),
    .C1(_11124_),
    .X(_02731_));
 sky130_fd_sc_hd__and2_2 _25310_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[483] ),
    .X(_11125_));
 sky130_fd_sc_hd__a221o_2 _25311_ (.A1(\ser_C.parallel_data[482] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[482] ),
    .C1(_11125_),
    .X(_02732_));
 sky130_fd_sc_hd__and2_2 _25312_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[484] ),
    .X(_11126_));
 sky130_fd_sc_hd__a221o_2 _25313_ (.A1(\ser_C.parallel_data[483] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[483] ),
    .C1(_11126_),
    .X(_02733_));
 sky130_fd_sc_hd__and2_2 _25314_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[485] ),
    .X(_11127_));
 sky130_fd_sc_hd__a221o_2 _25315_ (.A1(\ser_C.parallel_data[484] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[484] ),
    .C1(_11127_),
    .X(_02734_));
 sky130_fd_sc_hd__and2_2 _25316_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[486] ),
    .X(_11128_));
 sky130_fd_sc_hd__a221o_2 _25317_ (.A1(\ser_C.parallel_data[485] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[485] ),
    .C1(_11128_),
    .X(_02735_));
 sky130_fd_sc_hd__and2_2 _25318_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[487] ),
    .X(_11129_));
 sky130_fd_sc_hd__a221o_2 _25319_ (.A1(\ser_C.parallel_data[486] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[486] ),
    .C1(_11129_),
    .X(_02736_));
 sky130_fd_sc_hd__and2_2 _25320_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[488] ),
    .X(_11130_));
 sky130_fd_sc_hd__a221o_2 _25321_ (.A1(\ser_C.parallel_data[487] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[487] ),
    .C1(_11130_),
    .X(_02737_));
 sky130_fd_sc_hd__and2_2 _25322_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[489] ),
    .X(_11131_));
 sky130_fd_sc_hd__a221o_2 _25323_ (.A1(\ser_C.parallel_data[488] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[488] ),
    .C1(_11131_),
    .X(_02738_));
 sky130_fd_sc_hd__and2_2 _25324_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[490] ),
    .X(_11132_));
 sky130_fd_sc_hd__a221o_2 _25325_ (.A1(\ser_C.parallel_data[489] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[489] ),
    .C1(_11132_),
    .X(_02739_));
 sky130_fd_sc_hd__and2_2 _25326_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[491] ),
    .X(_11133_));
 sky130_fd_sc_hd__a221o_2 _25327_ (.A1(\ser_C.parallel_data[490] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[490] ),
    .C1(_11133_),
    .X(_02740_));
 sky130_fd_sc_hd__and2_2 _25328_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[492] ),
    .X(_11134_));
 sky130_fd_sc_hd__a221o_2 _25329_ (.A1(\ser_C.parallel_data[491] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[491] ),
    .C1(_11134_),
    .X(_02741_));
 sky130_fd_sc_hd__and2_2 _25330_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[493] ),
    .X(_11135_));
 sky130_fd_sc_hd__a221o_2 _25331_ (.A1(\ser_C.parallel_data[492] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[492] ),
    .C1(_11135_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_2 _25332_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[494] ),
    .X(_11136_));
 sky130_fd_sc_hd__a221o_2 _25333_ (.A1(\ser_C.parallel_data[493] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[493] ),
    .C1(_11136_),
    .X(_02743_));
 sky130_fd_sc_hd__and2_2 _25334_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[495] ),
    .X(_11137_));
 sky130_fd_sc_hd__a221o_2 _25335_ (.A1(\ser_C.parallel_data[494] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[494] ),
    .C1(_11137_),
    .X(_02744_));
 sky130_fd_sc_hd__and2_2 _25336_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[496] ),
    .X(_11138_));
 sky130_fd_sc_hd__a221o_2 _25337_ (.A1(\ser_C.parallel_data[495] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[495] ),
    .C1(_11138_),
    .X(_02745_));
 sky130_fd_sc_hd__and2_2 _25338_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[497] ),
    .X(_11139_));
 sky130_fd_sc_hd__a221o_2 _25339_ (.A1(\ser_C.parallel_data[496] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[496] ),
    .C1(_11139_),
    .X(_02746_));
 sky130_fd_sc_hd__and2_2 _25340_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[498] ),
    .X(_11140_));
 sky130_fd_sc_hd__a221o_2 _25341_ (.A1(\ser_C.parallel_data[497] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[497] ),
    .C1(_11140_),
    .X(_02747_));
 sky130_fd_sc_hd__and2_2 _25342_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[499] ),
    .X(_11141_));
 sky130_fd_sc_hd__a221o_2 _25343_ (.A1(\ser_C.parallel_data[498] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[498] ),
    .C1(_11141_),
    .X(_02748_));
 sky130_fd_sc_hd__and2_2 _25344_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[500] ),
    .X(_11142_));
 sky130_fd_sc_hd__a221o_2 _25345_ (.A1(\ser_C.parallel_data[499] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[499] ),
    .C1(_11142_),
    .X(_02749_));
 sky130_fd_sc_hd__and2_2 _25346_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[501] ),
    .X(_11143_));
 sky130_fd_sc_hd__a221o_2 _25347_ (.A1(\ser_C.parallel_data[500] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[500] ),
    .C1(_11143_),
    .X(_02750_));
 sky130_fd_sc_hd__and2_2 _25348_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[502] ),
    .X(_11144_));
 sky130_fd_sc_hd__a221o_2 _25349_ (.A1(\ser_C.parallel_data[501] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[501] ),
    .C1(_11144_),
    .X(_02751_));
 sky130_fd_sc_hd__and2_2 _25350_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[503] ),
    .X(_11145_));
 sky130_fd_sc_hd__a221o_2 _25351_ (.A1(\ser_C.parallel_data[502] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[502] ),
    .C1(_11145_),
    .X(_02752_));
 sky130_fd_sc_hd__and2_2 _25352_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[504] ),
    .X(_11146_));
 sky130_fd_sc_hd__a221o_2 _25353_ (.A1(\ser_C.parallel_data[503] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[503] ),
    .C1(_11146_),
    .X(_02753_));
 sky130_fd_sc_hd__and2_2 _25354_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[505] ),
    .X(_11147_));
 sky130_fd_sc_hd__a221o_2 _25355_ (.A1(\ser_C.parallel_data[504] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[504] ),
    .C1(_11147_),
    .X(_02754_));
 sky130_fd_sc_hd__and2_2 _25356_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[506] ),
    .X(_11148_));
 sky130_fd_sc_hd__a221o_2 _25357_ (.A1(\ser_C.parallel_data[505] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[505] ),
    .C1(_11148_),
    .X(_02755_));
 sky130_fd_sc_hd__and2_2 _25358_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[507] ),
    .X(_11149_));
 sky130_fd_sc_hd__a221o_2 _25359_ (.A1(\ser_C.parallel_data[506] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[506] ),
    .C1(_11149_),
    .X(_02756_));
 sky130_fd_sc_hd__and2_2 _25360_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[508] ),
    .X(_11150_));
 sky130_fd_sc_hd__a221o_2 _25361_ (.A1(\ser_C.parallel_data[507] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[507] ),
    .C1(_11150_),
    .X(_02757_));
 sky130_fd_sc_hd__and2_2 _25362_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[509] ),
    .X(_11151_));
 sky130_fd_sc_hd__a221o_2 _25363_ (.A1(\ser_C.parallel_data[508] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[508] ),
    .C1(_11151_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_2 _25364_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[510] ),
    .X(_11152_));
 sky130_fd_sc_hd__a221o_2 _25365_ (.A1(\ser_C.parallel_data[509] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[509] ),
    .C1(_11152_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_2 _25366_ (.A(C_out_frame_sync),
    .B(\ser_C.shift_reg[511] ),
    .X(_11153_));
 sky130_fd_sc_hd__a221o_2 _25367_ (.A1(\ser_C.parallel_data[510] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[510] ),
    .C1(_11153_),
    .X(_02760_));
 sky130_fd_sc_hd__a22o_2 _25368_ (.A1(\ser_C.parallel_data[511] ),
    .A2(_11302_),
    .B1(_10643_),
    .B2(\ser_C.shift_reg[511] ),
    .X(_02761_));
 sky130_fd_sc_hd__mux2_1 _25369_ (.A0(\systolic_inst.B_shift[18][0] ),
    .A1(\B_in[48] ),
    .S(_00008_),
    .X(_11154_));
 sky130_fd_sc_hd__mux2_1 _25370_ (.A0(_11154_),
    .A1(\systolic_inst.B_shift[14][0] ),
    .S(_11332_),
    .X(_02762_));
 sky130_fd_sc_hd__mux2_1 _25371_ (.A0(\systolic_inst.B_shift[18][1] ),
    .A1(\B_in[49] ),
    .S(_00008_),
    .X(_11155_));
 sky130_fd_sc_hd__mux2_1 _25372_ (.A0(_11155_),
    .A1(\systolic_inst.B_shift[14][1] ),
    .S(_11332_),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_1 _25373_ (.A0(\systolic_inst.B_shift[18][2] ),
    .A1(\B_in[50] ),
    .S(_00008_),
    .X(_11156_));
 sky130_fd_sc_hd__mux2_1 _25374_ (.A0(_11156_),
    .A1(\systolic_inst.B_shift[14][2] ),
    .S(_11332_),
    .X(_02764_));
 sky130_fd_sc_hd__mux2_1 _25375_ (.A0(\systolic_inst.B_shift[18][3] ),
    .A1(\B_in[51] ),
    .S(_00008_),
    .X(_11157_));
 sky130_fd_sc_hd__mux2_1 _25376_ (.A0(_11157_),
    .A1(\systolic_inst.B_shift[14][3] ),
    .S(_11332_),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _25377_ (.A0(\systolic_inst.B_shift[18][4] ),
    .A1(\B_in[52] ),
    .S(_00008_),
    .X(_11158_));
 sky130_fd_sc_hd__mux2_1 _25378_ (.A0(_11158_),
    .A1(\systolic_inst.B_shift[14][4] ),
    .S(_11332_),
    .X(_02766_));
 sky130_fd_sc_hd__mux2_1 _25379_ (.A0(\systolic_inst.B_shift[18][5] ),
    .A1(\B_in[53] ),
    .S(_00008_),
    .X(_11159_));
 sky130_fd_sc_hd__mux2_1 _25380_ (.A0(_11159_),
    .A1(\systolic_inst.B_shift[14][5] ),
    .S(_11332_),
    .X(_02767_));
 sky130_fd_sc_hd__mux2_1 _25381_ (.A0(\systolic_inst.B_shift[18][6] ),
    .A1(\B_in[54] ),
    .S(_00008_),
    .X(_11160_));
 sky130_fd_sc_hd__mux2_1 _25382_ (.A0(_11160_),
    .A1(\systolic_inst.B_shift[14][6] ),
    .S(_11332_),
    .X(_02768_));
 sky130_fd_sc_hd__mux2_1 _25383_ (.A0(\systolic_inst.B_shift[18][7] ),
    .A1(\B_in[55] ),
    .S(_00008_),
    .X(_11161_));
 sky130_fd_sc_hd__mux2_1 _25384_ (.A0(_11161_),
    .A1(\systolic_inst.B_shift[14][7] ),
    .S(_11332_),
    .X(_02769_));
 sky130_fd_sc_hd__mux2_1 _25385_ (.A0(\systolic_inst.A_shift[3][0] ),
    .A1(\A_in[16] ),
    .S(_00008_),
    .X(_11162_));
 sky130_fd_sc_hd__mux2_1 _25386_ (.A0(_11162_),
    .A1(\systolic_inst.A_shift[2][0] ),
    .S(_11332_),
    .X(_02770_));
 sky130_fd_sc_hd__mux2_1 _25387_ (.A0(\systolic_inst.A_shift[3][1] ),
    .A1(\A_in[17] ),
    .S(_00008_),
    .X(_11163_));
 sky130_fd_sc_hd__mux2_1 _25388_ (.A0(_11163_),
    .A1(\systolic_inst.A_shift[2][1] ),
    .S(_11332_),
    .X(_02771_));
 sky130_fd_sc_hd__mux2_1 _25389_ (.A0(\systolic_inst.A_shift[3][2] ),
    .A1(\A_in[18] ),
    .S(_00008_),
    .X(_11164_));
 sky130_fd_sc_hd__mux2_1 _25390_ (.A0(_11164_),
    .A1(\systolic_inst.A_shift[2][2] ),
    .S(_11332_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _25391_ (.A0(\systolic_inst.A_shift[3][3] ),
    .A1(\A_in[19] ),
    .S(_00008_),
    .X(_11165_));
 sky130_fd_sc_hd__mux2_1 _25392_ (.A0(_11165_),
    .A1(\systolic_inst.A_shift[2][3] ),
    .S(_11332_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _25393_ (.A0(\systolic_inst.A_shift[3][4] ),
    .A1(\A_in[20] ),
    .S(_00008_),
    .X(_11166_));
 sky130_fd_sc_hd__mux2_1 _25394_ (.A0(_11166_),
    .A1(\systolic_inst.A_shift[2][4] ),
    .S(_11332_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _25395_ (.A0(\systolic_inst.A_shift[3][5] ),
    .A1(\A_in[21] ),
    .S(_00008_),
    .X(_11167_));
 sky130_fd_sc_hd__mux2_1 _25396_ (.A0(_11167_),
    .A1(\systolic_inst.A_shift[2][5] ),
    .S(_11332_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _25397_ (.A0(\systolic_inst.A_shift[3][6] ),
    .A1(\A_in[22] ),
    .S(_00008_),
    .X(_11168_));
 sky130_fd_sc_hd__mux2_1 _25398_ (.A0(_11168_),
    .A1(\systolic_inst.A_shift[2][6] ),
    .S(_11332_),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_1 _25399_ (.A0(\systolic_inst.A_shift[3][7] ),
    .A1(\A_in[23] ),
    .S(_00008_),
    .X(_11169_));
 sky130_fd_sc_hd__mux2_1 _25400_ (.A0(_11169_),
    .A1(\systolic_inst.A_shift[2][7] ),
    .S(_11332_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _25401_ (.A0(\systolic_inst.A_shift[2][0] ),
    .A1(\A_in[8] ),
    .S(_00008_),
    .X(_11170_));
 sky130_fd_sc_hd__mux2_1 _25402_ (.A0(_11170_),
    .A1(\systolic_inst.A_shift[1][0] ),
    .S(_11332_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _25403_ (.A0(\systolic_inst.A_shift[2][1] ),
    .A1(\A_in[9] ),
    .S(_00008_),
    .X(_11171_));
 sky130_fd_sc_hd__mux2_1 _25404_ (.A0(_11171_),
    .A1(\systolic_inst.A_shift[1][1] ),
    .S(_11332_),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _25405_ (.A0(\systolic_inst.A_shift[2][2] ),
    .A1(\A_in[10] ),
    .S(_00008_),
    .X(_11172_));
 sky130_fd_sc_hd__mux2_1 _25406_ (.A0(_11172_),
    .A1(\systolic_inst.A_shift[1][2] ),
    .S(_11332_),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_1 _25407_ (.A0(\systolic_inst.A_shift[2][3] ),
    .A1(\A_in[11] ),
    .S(_00008_),
    .X(_11173_));
 sky130_fd_sc_hd__mux2_1 _25408_ (.A0(_11173_),
    .A1(\systolic_inst.A_shift[1][3] ),
    .S(_11332_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _25409_ (.A0(\systolic_inst.A_shift[2][4] ),
    .A1(\A_in[12] ),
    .S(_00008_),
    .X(_11174_));
 sky130_fd_sc_hd__mux2_1 _25410_ (.A0(_11174_),
    .A1(\systolic_inst.A_shift[1][4] ),
    .S(_11332_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _25411_ (.A0(\systolic_inst.A_shift[2][5] ),
    .A1(\A_in[13] ),
    .S(_00008_),
    .X(_11175_));
 sky130_fd_sc_hd__mux2_1 _25412_ (.A0(_11175_),
    .A1(\systolic_inst.A_shift[1][5] ),
    .S(_11332_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _25413_ (.A0(\systolic_inst.A_shift[2][6] ),
    .A1(\A_in[14] ),
    .S(_00008_),
    .X(_11176_));
 sky130_fd_sc_hd__mux2_1 _25414_ (.A0(_11176_),
    .A1(\systolic_inst.A_shift[1][6] ),
    .S(_11332_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _25415_ (.A0(\systolic_inst.A_shift[2][7] ),
    .A1(\A_in[15] ),
    .S(_00008_),
    .X(_11177_));
 sky130_fd_sc_hd__mux2_1 _25416_ (.A0(_11177_),
    .A1(\systolic_inst.A_shift[1][7] ),
    .S(_11332_),
    .X(_02785_));
 sky130_fd_sc_hd__mux2_1 _25417_ (.A0(\systolic_inst.A_shift[1][0] ),
    .A1(\A_in[0] ),
    .S(_00008_),
    .X(_11178_));
 sky130_fd_sc_hd__mux2_1 _25418_ (.A0(_11178_),
    .A1(\systolic_inst.A_shift[0][0] ),
    .S(_11332_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _25419_ (.A0(\systolic_inst.A_shift[1][1] ),
    .A1(\A_in[1] ),
    .S(_00008_),
    .X(_11179_));
 sky130_fd_sc_hd__mux2_1 _25420_ (.A0(_11179_),
    .A1(\systolic_inst.A_shift[0][1] ),
    .S(_11332_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _25421_ (.A0(\systolic_inst.A_shift[1][2] ),
    .A1(\A_in[2] ),
    .S(_00008_),
    .X(_11180_));
 sky130_fd_sc_hd__mux2_1 _25422_ (.A0(_11180_),
    .A1(\systolic_inst.A_shift[0][2] ),
    .S(_11332_),
    .X(_02788_));
 sky130_fd_sc_hd__mux2_1 _25423_ (.A0(\systolic_inst.A_shift[1][3] ),
    .A1(\A_in[3] ),
    .S(_00008_),
    .X(_11181_));
 sky130_fd_sc_hd__mux2_1 _25424_ (.A0(_11181_),
    .A1(\systolic_inst.A_shift[0][3] ),
    .S(_11332_),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_1 _25425_ (.A0(\systolic_inst.A_shift[1][4] ),
    .A1(\A_in[4] ),
    .S(_00008_),
    .X(_11182_));
 sky130_fd_sc_hd__mux2_1 _25426_ (.A0(_11182_),
    .A1(\systolic_inst.A_shift[0][4] ),
    .S(_11332_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _25427_ (.A0(\systolic_inst.A_shift[1][5] ),
    .A1(\A_in[5] ),
    .S(_00008_),
    .X(_11183_));
 sky130_fd_sc_hd__mux2_1 _25428_ (.A0(_11183_),
    .A1(\systolic_inst.A_shift[0][5] ),
    .S(_11332_),
    .X(_02791_));
 sky130_fd_sc_hd__mux2_1 _25429_ (.A0(\systolic_inst.A_shift[1][6] ),
    .A1(\A_in[6] ),
    .S(_00008_),
    .X(_11184_));
 sky130_fd_sc_hd__mux2_1 _25430_ (.A0(_11184_),
    .A1(\systolic_inst.A_shift[0][6] ),
    .S(_11332_),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_1 _25431_ (.A0(\systolic_inst.A_shift[1][7] ),
    .A1(\A_in[7] ),
    .S(_00008_),
    .X(_11185_));
 sky130_fd_sc_hd__mux2_1 _25432_ (.A0(_11185_),
    .A1(\systolic_inst.A_shift[0][7] ),
    .S(_11332_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_1 _25433_ (.A0(\systolic_inst.ce_local ),
    .A1(_11307_),
    .S(\systolic_inst.cycle_cnt[0] ),
    .X(_02794_));
 sky130_fd_sc_hd__nand2_2 _25434_ (.A(\systolic_inst.cycle_cnt[1] ),
    .B(\systolic_inst.cycle_cnt[0] ),
    .Y(_11186_));
 sky130_fd_sc_hd__or2_2 _25435_ (.A(\systolic_inst.cycle_cnt[1] ),
    .B(\systolic_inst.cycle_cnt[0] ),
    .X(_11187_));
 sky130_fd_sc_hd__a32o_2 _25436_ (.A1(\systolic_inst.ce_local ),
    .A2(_11186_),
    .A3(_11187_),
    .B1(_11307_),
    .B2(\systolic_inst.cycle_cnt[1] ),
    .X(_02795_));
 sky130_fd_sc_hd__a31o_2 _25437_ (.A1(\systolic_inst.cycle_cnt[1] ),
    .A2(\systolic_inst.cycle_cnt[0] ),
    .A3(_11306_),
    .B1(\systolic_inst.cycle_cnt[2] ),
    .X(_11188_));
 sky130_fd_sc_hd__or3_2 _25438_ (.A(_11257_),
    .B(_11258_),
    .C(_11186_),
    .X(_11189_));
 sky130_fd_sc_hd__and3_2 _25439_ (.A(_11279_),
    .B(_11188_),
    .C(_11189_),
    .X(_02796_));
 sky130_fd_sc_hd__and4_2 _25440_ (.A(\systolic_inst.cycle_cnt[1] ),
    .B(\systolic_inst.cycle_cnt[0] ),
    .C(\systolic_inst.cycle_cnt[3] ),
    .D(\systolic_inst.cycle_cnt[2] ),
    .X(_11190_));
 sky130_fd_sc_hd__and2_2 _25441_ (.A(\systolic_inst.ce_local ),
    .B(_11190_),
    .X(_11191_));
 sky130_fd_sc_hd__nand2_2 _25442_ (.A(\systolic_inst.cycle_cnt[3] ),
    .B(_11279_),
    .Y(_11192_));
 sky130_fd_sc_hd__a21oi_2 _25443_ (.A1(_11189_),
    .A2(_11192_),
    .B1(_11191_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand2_2 _25444_ (.A(\systolic_inst.cycle_cnt[4] ),
    .B(_11191_),
    .Y(_11193_));
 sky130_fd_sc_hd__a21o_2 _25445_ (.A1(\systolic_inst.cycle_cnt[4] ),
    .A2(_11279_),
    .B1(_11191_),
    .X(_11194_));
 sky130_fd_sc_hd__and2_2 _25446_ (.A(_11193_),
    .B(_11194_),
    .X(_02798_));
 sky130_fd_sc_hd__and3_2 _25447_ (.A(\systolic_inst.cycle_cnt[5] ),
    .B(\systolic_inst.cycle_cnt[4] ),
    .C(_11190_),
    .X(_11195_));
 sky130_fd_sc_hd__and2_2 _25448_ (.A(\systolic_inst.ce_local ),
    .B(_11195_),
    .X(_11196_));
 sky130_fd_sc_hd__nor2_2 _25449_ (.A(_00008_),
    .B(_11196_),
    .Y(_11197_));
 sky130_fd_sc_hd__a2bb2o_2 _25450_ (.A1_N(_11193_),
    .A2_N(_11196_),
    .B1(_11197_),
    .B2(\systolic_inst.cycle_cnt[5] ),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _25451_ (.A0(_11196_),
    .A1(_11197_),
    .S(\systolic_inst.cycle_cnt[6] ),
    .X(_02800_));
 sky130_fd_sc_hd__a31o_2 _25452_ (.A1(\systolic_inst.cycle_cnt[6] ),
    .A2(_11306_),
    .A3(_11195_),
    .B1(\systolic_inst.cycle_cnt[7] ),
    .X(_11198_));
 sky130_fd_sc_hd__and3_2 _25453_ (.A(\systolic_inst.cycle_cnt[7] ),
    .B(\systolic_inst.cycle_cnt[6] ),
    .C(_11195_),
    .X(_11199_));
 sky130_fd_sc_hd__and2_2 _25454_ (.A(\systolic_inst.ce_local ),
    .B(_11199_),
    .X(_11200_));
 sky130_fd_sc_hd__nor2_2 _25455_ (.A(_00008_),
    .B(_11200_),
    .Y(_11201_));
 sky130_fd_sc_hd__and2_2 _25456_ (.A(_11198_),
    .B(_11201_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _25457_ (.A0(_11200_),
    .A1(_11201_),
    .S(\systolic_inst.cycle_cnt[8] ),
    .X(_02802_));
 sky130_fd_sc_hd__and2_2 _25458_ (.A(\systolic_inst.cycle_cnt[9] ),
    .B(\systolic_inst.cycle_cnt[8] ),
    .X(_11202_));
 sky130_fd_sc_hd__and3_2 _25459_ (.A(\systolic_inst.ce_local ),
    .B(_11199_),
    .C(_11202_),
    .X(_11203_));
 sky130_fd_sc_hd__nor2_2 _25460_ (.A(_00008_),
    .B(_11203_),
    .Y(_11204_));
 sky130_fd_sc_hd__a31o_2 _25461_ (.A1(\systolic_inst.cycle_cnt[8] ),
    .A2(_11306_),
    .A3(_11199_),
    .B1(\systolic_inst.cycle_cnt[9] ),
    .X(_11205_));
 sky130_fd_sc_hd__and2_2 _25462_ (.A(_11204_),
    .B(_11205_),
    .X(_02803_));
 sky130_fd_sc_hd__mux2_1 _25463_ (.A0(_11203_),
    .A1(_11204_),
    .S(\systolic_inst.cycle_cnt[10] ),
    .X(_02804_));
 sky130_fd_sc_hd__and4_2 _25464_ (.A(\systolic_inst.cycle_cnt[11] ),
    .B(\systolic_inst.cycle_cnt[10] ),
    .C(_11199_),
    .D(_11202_),
    .X(_11206_));
 sky130_fd_sc_hd__and2_2 _25465_ (.A(\systolic_inst.ce_local ),
    .B(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__nor2_2 _25466_ (.A(_00008_),
    .B(_11207_),
    .Y(_11208_));
 sky130_fd_sc_hd__a41o_2 _25467_ (.A1(\systolic_inst.cycle_cnt[10] ),
    .A2(_11306_),
    .A3(_11199_),
    .A4(_11202_),
    .B1(\systolic_inst.cycle_cnt[11] ),
    .X(_11209_));
 sky130_fd_sc_hd__and2_2 _25468_ (.A(_11208_),
    .B(_11209_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _25469_ (.A0(_11207_),
    .A1(_11208_),
    .S(\systolic_inst.cycle_cnt[12] ),
    .X(_02806_));
 sky130_fd_sc_hd__and3_2 _25470_ (.A(\systolic_inst.cycle_cnt[13] ),
    .B(\systolic_inst.cycle_cnt[12] ),
    .C(_11206_),
    .X(_11210_));
 sky130_fd_sc_hd__and2_2 _25471_ (.A(\systolic_inst.ce_local ),
    .B(_11210_),
    .X(_11211_));
 sky130_fd_sc_hd__nor2_2 _25472_ (.A(_00008_),
    .B(_11211_),
    .Y(_11212_));
 sky130_fd_sc_hd__a31o_2 _25473_ (.A1(\systolic_inst.cycle_cnt[12] ),
    .A2(_11306_),
    .A3(_11206_),
    .B1(\systolic_inst.cycle_cnt[13] ),
    .X(_11213_));
 sky130_fd_sc_hd__and2_2 _25474_ (.A(_11212_),
    .B(_11213_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _25475_ (.A0(_11211_),
    .A1(_11212_),
    .S(\systolic_inst.cycle_cnt[14] ),
    .X(_02808_));
 sky130_fd_sc_hd__a31o_2 _25476_ (.A1(\systolic_inst.cycle_cnt[14] ),
    .A2(_11306_),
    .A3(_11210_),
    .B1(\systolic_inst.cycle_cnt[15] ),
    .X(_11214_));
 sky130_fd_sc_hd__and3_2 _25477_ (.A(\systolic_inst.cycle_cnt[15] ),
    .B(\systolic_inst.cycle_cnt[14] ),
    .C(_11210_),
    .X(_11215_));
 sky130_fd_sc_hd__and2_2 _25478_ (.A(\systolic_inst.ce_local ),
    .B(_11215_),
    .X(_11216_));
 sky130_fd_sc_hd__nand2_2 _25479_ (.A(\systolic_inst.ce_local ),
    .B(_11215_),
    .Y(_11217_));
 sky130_fd_sc_hd__and3_2 _25480_ (.A(_11279_),
    .B(_11214_),
    .C(_11217_),
    .X(_02809_));
 sky130_fd_sc_hd__or3b_2 _25481_ (.A(_00008_),
    .B(_11216_),
    .C_N(\systolic_inst.cycle_cnt[16] ),
    .X(_11218_));
 sky130_fd_sc_hd__o21ai_2 _25482_ (.A1(\systolic_inst.cycle_cnt[16] ),
    .A2(_11217_),
    .B1(_11218_),
    .Y(_02810_));
 sky130_fd_sc_hd__a31o_2 _25483_ (.A1(\systolic_inst.cycle_cnt[16] ),
    .A2(_11306_),
    .A3(_11215_),
    .B1(\systolic_inst.cycle_cnt[17] ),
    .X(_11219_));
 sky130_fd_sc_hd__and3_2 _25484_ (.A(\systolic_inst.cycle_cnt[17] ),
    .B(\systolic_inst.cycle_cnt[16] ),
    .C(_11216_),
    .X(_11220_));
 sky130_fd_sc_hd__inv_2 _25485_ (.A(_11220_),
    .Y(_11221_));
 sky130_fd_sc_hd__and3_2 _25486_ (.A(_11279_),
    .B(_11219_),
    .C(_11221_),
    .X(_02811_));
 sky130_fd_sc_hd__a41o_2 _25487_ (.A1(\systolic_inst.cycle_cnt[17] ),
    .A2(\systolic_inst.cycle_cnt[16] ),
    .A3(_11306_),
    .A4(_11215_),
    .B1(\systolic_inst.cycle_cnt[18] ),
    .X(_11222_));
 sky130_fd_sc_hd__and2_2 _25488_ (.A(\systolic_inst.cycle_cnt[18] ),
    .B(_11220_),
    .X(_11223_));
 sky130_fd_sc_hd__nor2_2 _25489_ (.A(_00008_),
    .B(_11223_),
    .Y(_11224_));
 sky130_fd_sc_hd__and2_2 _25490_ (.A(_11222_),
    .B(_11224_),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _25491_ (.A0(_11223_),
    .A1(_11224_),
    .S(\systolic_inst.cycle_cnt[19] ),
    .X(_02813_));
 sky130_fd_sc_hd__and3_2 _25492_ (.A(\systolic_inst.cycle_cnt[20] ),
    .B(\systolic_inst.cycle_cnt[19] ),
    .C(_11223_),
    .X(_11225_));
 sky130_fd_sc_hd__a22oi_2 _25493_ (.A1(\systolic_inst.cycle_cnt[20] ),
    .A2(_11279_),
    .B1(_11223_),
    .B2(\systolic_inst.cycle_cnt[19] ),
    .Y(_11226_));
 sky130_fd_sc_hd__nor2_2 _25494_ (.A(_11225_),
    .B(_11226_),
    .Y(_02814_));
 sky130_fd_sc_hd__nor2_2 _25495_ (.A(_00008_),
    .B(_11225_),
    .Y(_11227_));
 sky130_fd_sc_hd__mux2_1 _25496_ (.A0(_11225_),
    .A1(_11227_),
    .S(\systolic_inst.cycle_cnt[21] ),
    .X(_02815_));
 sky130_fd_sc_hd__and3_2 _25497_ (.A(\systolic_inst.cycle_cnt[22] ),
    .B(\systolic_inst.cycle_cnt[21] ),
    .C(_11225_),
    .X(_11228_));
 sky130_fd_sc_hd__a22oi_2 _25498_ (.A1(\systolic_inst.cycle_cnt[22] ),
    .A2(_11279_),
    .B1(_11225_),
    .B2(\systolic_inst.cycle_cnt[21] ),
    .Y(_11229_));
 sky130_fd_sc_hd__nor2_2 _25499_ (.A(_11228_),
    .B(_11229_),
    .Y(_02816_));
 sky130_fd_sc_hd__nor2_2 _25500_ (.A(_00008_),
    .B(_11228_),
    .Y(_11230_));
 sky130_fd_sc_hd__mux2_1 _25501_ (.A0(_11228_),
    .A1(_11230_),
    .S(\systolic_inst.cycle_cnt[23] ),
    .X(_02817_));
 sky130_fd_sc_hd__and3_2 _25502_ (.A(\systolic_inst.cycle_cnt[24] ),
    .B(\systolic_inst.cycle_cnt[23] ),
    .C(_11228_),
    .X(_11231_));
 sky130_fd_sc_hd__a22oi_2 _25503_ (.A1(\systolic_inst.cycle_cnt[24] ),
    .A2(_11279_),
    .B1(_11228_),
    .B2(\systolic_inst.cycle_cnt[23] ),
    .Y(_11232_));
 sky130_fd_sc_hd__nor2_2 _25504_ (.A(_11231_),
    .B(_11232_),
    .Y(_02818_));
 sky130_fd_sc_hd__and2_2 _25505_ (.A(\systolic_inst.cycle_cnt[25] ),
    .B(_11231_),
    .X(_11233_));
 sky130_fd_sc_hd__a21oi_2 _25506_ (.A1(\systolic_inst.cycle_cnt[25] ),
    .A2(_11279_),
    .B1(_11231_),
    .Y(_11234_));
 sky130_fd_sc_hd__nor2_2 _25507_ (.A(_11233_),
    .B(_11234_),
    .Y(_02819_));
 sky130_fd_sc_hd__nor2_2 _25508_ (.A(_00008_),
    .B(_11233_),
    .Y(_11235_));
 sky130_fd_sc_hd__mux2_1 _25509_ (.A0(_11233_),
    .A1(_11235_),
    .S(\systolic_inst.cycle_cnt[26] ),
    .X(_02820_));
 sky130_fd_sc_hd__a22oi_2 _25510_ (.A1(\systolic_inst.cycle_cnt[27] ),
    .A2(_11279_),
    .B1(_11233_),
    .B2(\systolic_inst.cycle_cnt[26] ),
    .Y(_11236_));
 sky130_fd_sc_hd__a31oi_2 _25511_ (.A1(\systolic_inst.cycle_cnt[27] ),
    .A2(\systolic_inst.cycle_cnt[26] ),
    .A3(_11233_),
    .B1(_11236_),
    .Y(_02821_));
 sky130_fd_sc_hd__and4_2 _25512_ (.A(\systolic_inst.cycle_cnt[28] ),
    .B(\systolic_inst.cycle_cnt[27] ),
    .C(\systolic_inst.cycle_cnt[26] ),
    .D(_11233_),
    .X(_11237_));
 sky130_fd_sc_hd__a32o_2 _25513_ (.A1(\systolic_inst.cycle_cnt[27] ),
    .A2(\systolic_inst.cycle_cnt[26] ),
    .A3(_11233_),
    .B1(_11279_),
    .B2(\systolic_inst.cycle_cnt[28] ),
    .X(_11238_));
 sky130_fd_sc_hd__and2b_2 _25514_ (.A_N(_11237_),
    .B(_11238_),
    .X(_02822_));
 sky130_fd_sc_hd__and2_2 _25515_ (.A(\systolic_inst.cycle_cnt[29] ),
    .B(_11237_),
    .X(_11239_));
 sky130_fd_sc_hd__a21oi_2 _25516_ (.A1(\systolic_inst.cycle_cnt[29] ),
    .A2(_11279_),
    .B1(_11237_),
    .Y(_11240_));
 sky130_fd_sc_hd__nor2_2 _25517_ (.A(_11239_),
    .B(_11240_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_2 _25518_ (.A(\systolic_inst.cycle_cnt[30] ),
    .B(_11239_),
    .Y(_11241_));
 sky130_fd_sc_hd__a21o_2 _25519_ (.A1(\systolic_inst.cycle_cnt[30] ),
    .A2(_11279_),
    .B1(_11239_),
    .X(_11242_));
 sky130_fd_sc_hd__and2_2 _25520_ (.A(_11241_),
    .B(_11242_),
    .X(_02824_));
 sky130_fd_sc_hd__nand2_2 _25521_ (.A(\systolic_inst.cycle_cnt[31] ),
    .B(_11279_),
    .Y(_11243_));
 sky130_fd_sc_hd__mux2_1 _25522_ (.A0(\systolic_inst.cycle_cnt[31] ),
    .A1(_11243_),
    .S(_11241_),
    .X(_11244_));
 sky130_fd_sc_hd__inv_2 _25523_ (.A(_11244_),
    .Y(_02825_));
 sky130_fd_sc_hd__mux2_1 _25524_ (.A0(\systolic_inst.acc_wires[0][0] ),
    .A1(\C_out[0] ),
    .S(_11297_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _25525_ (.A0(\systolic_inst.acc_wires[0][1] ),
    .A1(\C_out[1] ),
    .S(_11297_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _25526_ (.A0(\systolic_inst.acc_wires[0][2] ),
    .A1(\C_out[2] ),
    .S(_11297_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _25527_ (.A0(\systolic_inst.acc_wires[0][3] ),
    .A1(\C_out[3] ),
    .S(_11297_),
    .X(_02829_));
 sky130_fd_sc_hd__mux2_1 _25528_ (.A0(\systolic_inst.acc_wires[0][4] ),
    .A1(\C_out[4] ),
    .S(_11297_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _25529_ (.A0(\systolic_inst.acc_wires[0][5] ),
    .A1(\C_out[5] ),
    .S(_11297_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _25530_ (.A0(\systolic_inst.acc_wires[0][6] ),
    .A1(\C_out[6] ),
    .S(_11297_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _25531_ (.A0(\systolic_inst.acc_wires[0][7] ),
    .A1(\C_out[7] ),
    .S(_11297_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _25532_ (.A0(\systolic_inst.acc_wires[0][8] ),
    .A1(\C_out[8] ),
    .S(_11297_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _25533_ (.A0(\systolic_inst.acc_wires[0][9] ),
    .A1(\C_out[9] ),
    .S(_11297_),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _25534_ (.A0(\systolic_inst.acc_wires[0][10] ),
    .A1(\C_out[10] ),
    .S(_11297_),
    .X(_02836_));
 sky130_fd_sc_hd__mux2_1 _25535_ (.A0(\systolic_inst.acc_wires[0][11] ),
    .A1(\C_out[11] ),
    .S(_11297_),
    .X(_02837_));
 sky130_fd_sc_hd__mux2_1 _25536_ (.A0(\systolic_inst.acc_wires[0][12] ),
    .A1(\C_out[12] ),
    .S(_11297_),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_1 _25537_ (.A0(\systolic_inst.acc_wires[0][13] ),
    .A1(\C_out[13] ),
    .S(_11297_),
    .X(_02839_));
 sky130_fd_sc_hd__mux2_1 _25538_ (.A0(\systolic_inst.acc_wires[0][14] ),
    .A1(\C_out[14] ),
    .S(_11297_),
    .X(_02840_));
 sky130_fd_sc_hd__mux2_1 _25539_ (.A0(\systolic_inst.acc_wires[0][15] ),
    .A1(\C_out[15] ),
    .S(_11297_),
    .X(_02841_));
 sky130_fd_sc_hd__mux2_1 _25540_ (.A0(\systolic_inst.acc_wires[0][16] ),
    .A1(\C_out[16] ),
    .S(_11297_),
    .X(_02842_));
 sky130_fd_sc_hd__mux2_1 _25541_ (.A0(\systolic_inst.acc_wires[0][17] ),
    .A1(\C_out[17] ),
    .S(_11297_),
    .X(_02843_));
 sky130_fd_sc_hd__mux2_1 _25542_ (.A0(\systolic_inst.acc_wires[0][18] ),
    .A1(\C_out[18] ),
    .S(_11297_),
    .X(_02844_));
 sky130_fd_sc_hd__mux2_1 _25543_ (.A0(\systolic_inst.acc_wires[0][19] ),
    .A1(\C_out[19] ),
    .S(_11297_),
    .X(_02845_));
 sky130_fd_sc_hd__mux2_1 _25544_ (.A0(\systolic_inst.acc_wires[0][20] ),
    .A1(\C_out[20] ),
    .S(_11297_),
    .X(_02846_));
 sky130_fd_sc_hd__mux2_1 _25545_ (.A0(\systolic_inst.acc_wires[0][21] ),
    .A1(\C_out[21] ),
    .S(_11297_),
    .X(_02847_));
 sky130_fd_sc_hd__mux2_1 _25546_ (.A0(\systolic_inst.acc_wires[0][22] ),
    .A1(\C_out[22] ),
    .S(_11297_),
    .X(_02848_));
 sky130_fd_sc_hd__mux2_1 _25547_ (.A0(\systolic_inst.acc_wires[0][23] ),
    .A1(\C_out[23] ),
    .S(_11297_),
    .X(_02849_));
 sky130_fd_sc_hd__mux2_1 _25548_ (.A0(\systolic_inst.acc_wires[0][24] ),
    .A1(\C_out[24] ),
    .S(_11297_),
    .X(_02850_));
 sky130_fd_sc_hd__mux2_1 _25549_ (.A0(\systolic_inst.acc_wires[0][25] ),
    .A1(\C_out[25] ),
    .S(_11297_),
    .X(_02851_));
 sky130_fd_sc_hd__mux2_1 _25550_ (.A0(\systolic_inst.acc_wires[0][26] ),
    .A1(\C_out[26] ),
    .S(_11297_),
    .X(_02852_));
 sky130_fd_sc_hd__mux2_1 _25551_ (.A0(\systolic_inst.acc_wires[0][27] ),
    .A1(\C_out[27] ),
    .S(_11297_),
    .X(_02853_));
 sky130_fd_sc_hd__mux2_1 _25552_ (.A0(\systolic_inst.acc_wires[0][28] ),
    .A1(\C_out[28] ),
    .S(_11297_),
    .X(_02854_));
 sky130_fd_sc_hd__mux2_1 _25553_ (.A0(\systolic_inst.acc_wires[0][29] ),
    .A1(\C_out[29] ),
    .S(_11297_),
    .X(_02855_));
 sky130_fd_sc_hd__mux2_1 _25554_ (.A0(\systolic_inst.acc_wires[0][30] ),
    .A1(\C_out[30] ),
    .S(_11297_),
    .X(_02856_));
 sky130_fd_sc_hd__mux2_1 _25555_ (.A0(\systolic_inst.acc_wires[0][31] ),
    .A1(\C_out[31] ),
    .S(_11297_),
    .X(_02857_));
 sky130_fd_sc_hd__mux2_1 _25556_ (.A0(\systolic_inst.acc_wires[1][0] ),
    .A1(\C_out[32] ),
    .S(_11297_),
    .X(_02858_));
 sky130_fd_sc_hd__mux2_1 _25557_ (.A0(\systolic_inst.acc_wires[1][1] ),
    .A1(\C_out[33] ),
    .S(_11297_),
    .X(_02859_));
 sky130_fd_sc_hd__mux2_1 _25558_ (.A0(\systolic_inst.acc_wires[1][2] ),
    .A1(\C_out[34] ),
    .S(_11297_),
    .X(_02860_));
 sky130_fd_sc_hd__mux2_1 _25559_ (.A0(\systolic_inst.acc_wires[1][3] ),
    .A1(\C_out[35] ),
    .S(_11297_),
    .X(_02861_));
 sky130_fd_sc_hd__mux2_1 _25560_ (.A0(\systolic_inst.acc_wires[1][4] ),
    .A1(\C_out[36] ),
    .S(_11297_),
    .X(_02862_));
 sky130_fd_sc_hd__mux2_1 _25561_ (.A0(\systolic_inst.acc_wires[1][5] ),
    .A1(\C_out[37] ),
    .S(_11297_),
    .X(_02863_));
 sky130_fd_sc_hd__mux2_1 _25562_ (.A0(\systolic_inst.acc_wires[1][6] ),
    .A1(\C_out[38] ),
    .S(_11297_),
    .X(_02864_));
 sky130_fd_sc_hd__mux2_1 _25563_ (.A0(\systolic_inst.acc_wires[1][7] ),
    .A1(\C_out[39] ),
    .S(_11297_),
    .X(_02865_));
 sky130_fd_sc_hd__mux2_1 _25564_ (.A0(\systolic_inst.acc_wires[1][8] ),
    .A1(\C_out[40] ),
    .S(_11297_),
    .X(_02866_));
 sky130_fd_sc_hd__mux2_1 _25565_ (.A0(\systolic_inst.acc_wires[1][9] ),
    .A1(\C_out[41] ),
    .S(_11297_),
    .X(_02867_));
 sky130_fd_sc_hd__mux2_1 _25566_ (.A0(\systolic_inst.acc_wires[1][10] ),
    .A1(\C_out[42] ),
    .S(_11297_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _25567_ (.A0(\systolic_inst.acc_wires[1][11] ),
    .A1(\C_out[43] ),
    .S(_11297_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_1 _25568_ (.A0(\systolic_inst.acc_wires[1][12] ),
    .A1(\C_out[44] ),
    .S(_11297_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _25569_ (.A0(\systolic_inst.acc_wires[1][13] ),
    .A1(\C_out[45] ),
    .S(_11297_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _25570_ (.A0(\systolic_inst.acc_wires[1][14] ),
    .A1(\C_out[46] ),
    .S(_11297_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _25571_ (.A0(\systolic_inst.acc_wires[1][15] ),
    .A1(\C_out[47] ),
    .S(_11297_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _25572_ (.A0(\systolic_inst.acc_wires[1][16] ),
    .A1(\C_out[48] ),
    .S(_11297_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _25573_ (.A0(\systolic_inst.acc_wires[1][17] ),
    .A1(\C_out[49] ),
    .S(_11297_),
    .X(_02875_));
 sky130_fd_sc_hd__mux2_1 _25574_ (.A0(\systolic_inst.acc_wires[1][18] ),
    .A1(\C_out[50] ),
    .S(_11297_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _25575_ (.A0(\systolic_inst.acc_wires[1][19] ),
    .A1(\C_out[51] ),
    .S(_11297_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _25576_ (.A0(\systolic_inst.acc_wires[1][20] ),
    .A1(\C_out[52] ),
    .S(_11297_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _25577_ (.A0(\systolic_inst.acc_wires[1][21] ),
    .A1(\C_out[53] ),
    .S(_11297_),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _25578_ (.A0(\systolic_inst.acc_wires[1][22] ),
    .A1(\C_out[54] ),
    .S(_11297_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _25579_ (.A0(\systolic_inst.acc_wires[1][23] ),
    .A1(\C_out[55] ),
    .S(_11297_),
    .X(_02881_));
 sky130_fd_sc_hd__mux2_1 _25580_ (.A0(\systolic_inst.acc_wires[1][24] ),
    .A1(\C_out[56] ),
    .S(_11297_),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _25581_ (.A0(\systolic_inst.acc_wires[1][25] ),
    .A1(\C_out[57] ),
    .S(_11297_),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _25582_ (.A0(\systolic_inst.acc_wires[1][26] ),
    .A1(\C_out[58] ),
    .S(_11297_),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_1 _25583_ (.A0(\systolic_inst.acc_wires[1][27] ),
    .A1(\C_out[59] ),
    .S(_11297_),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_1 _25584_ (.A0(\systolic_inst.acc_wires[1][28] ),
    .A1(\C_out[60] ),
    .S(_11297_),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_1 _25585_ (.A0(\systolic_inst.acc_wires[1][29] ),
    .A1(\C_out[61] ),
    .S(_11297_),
    .X(_02887_));
 sky130_fd_sc_hd__mux2_1 _25586_ (.A0(\systolic_inst.acc_wires[1][30] ),
    .A1(\C_out[62] ),
    .S(_11297_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _25587_ (.A0(\systolic_inst.acc_wires[1][31] ),
    .A1(\C_out[63] ),
    .S(_11297_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_1 _25588_ (.A0(\systolic_inst.acc_wires[2][0] ),
    .A1(\C_out[64] ),
    .S(_11297_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_1 _25589_ (.A0(\systolic_inst.acc_wires[2][1] ),
    .A1(\C_out[65] ),
    .S(_11297_),
    .X(_02891_));
 sky130_fd_sc_hd__mux2_1 _25590_ (.A0(\systolic_inst.acc_wires[2][2] ),
    .A1(\C_out[66] ),
    .S(_11297_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _25591_ (.A0(\systolic_inst.acc_wires[2][3] ),
    .A1(\C_out[67] ),
    .S(_11297_),
    .X(_02893_));
 sky130_fd_sc_hd__mux2_1 _25592_ (.A0(\systolic_inst.acc_wires[2][4] ),
    .A1(\C_out[68] ),
    .S(_11297_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _25593_ (.A0(\systolic_inst.acc_wires[2][5] ),
    .A1(\C_out[69] ),
    .S(_11297_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _25594_ (.A0(\systolic_inst.acc_wires[2][6] ),
    .A1(\C_out[70] ),
    .S(_11297_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _25595_ (.A0(\systolic_inst.acc_wires[2][7] ),
    .A1(\C_out[71] ),
    .S(_11297_),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_1 _25596_ (.A0(\systolic_inst.acc_wires[2][8] ),
    .A1(\C_out[72] ),
    .S(_11297_),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_1 _25597_ (.A0(\systolic_inst.acc_wires[2][9] ),
    .A1(\C_out[73] ),
    .S(_11297_),
    .X(_02899_));
 sky130_fd_sc_hd__mux2_1 _25598_ (.A0(\systolic_inst.acc_wires[2][10] ),
    .A1(\C_out[74] ),
    .S(_11297_),
    .X(_02900_));
 sky130_fd_sc_hd__mux2_1 _25599_ (.A0(\systolic_inst.acc_wires[2][11] ),
    .A1(\C_out[75] ),
    .S(_11297_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _25600_ (.A0(\systolic_inst.acc_wires[2][12] ),
    .A1(\C_out[76] ),
    .S(_11297_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_1 _25601_ (.A0(\systolic_inst.acc_wires[2][13] ),
    .A1(\C_out[77] ),
    .S(_11297_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _25602_ (.A0(\systolic_inst.acc_wires[2][14] ),
    .A1(\C_out[78] ),
    .S(_11297_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _25603_ (.A0(\systolic_inst.acc_wires[2][15] ),
    .A1(\C_out[79] ),
    .S(_11297_),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_1 _25604_ (.A0(\systolic_inst.acc_wires[2][16] ),
    .A1(\C_out[80] ),
    .S(_11297_),
    .X(_02906_));
 sky130_fd_sc_hd__mux2_1 _25605_ (.A0(\systolic_inst.acc_wires[2][17] ),
    .A1(\C_out[81] ),
    .S(_11297_),
    .X(_02907_));
 sky130_fd_sc_hd__mux2_1 _25606_ (.A0(\systolic_inst.acc_wires[2][18] ),
    .A1(\C_out[82] ),
    .S(_11297_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _25607_ (.A0(\systolic_inst.acc_wires[2][19] ),
    .A1(\C_out[83] ),
    .S(_11297_),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_1 _25608_ (.A0(\systolic_inst.acc_wires[2][20] ),
    .A1(\C_out[84] ),
    .S(_11297_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _25609_ (.A0(\systolic_inst.acc_wires[2][21] ),
    .A1(\C_out[85] ),
    .S(_11297_),
    .X(_02911_));
 sky130_fd_sc_hd__mux2_1 _25610_ (.A0(\systolic_inst.acc_wires[2][22] ),
    .A1(\C_out[86] ),
    .S(_11297_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _25611_ (.A0(\systolic_inst.acc_wires[2][23] ),
    .A1(\C_out[87] ),
    .S(_11297_),
    .X(_02913_));
 sky130_fd_sc_hd__mux2_1 _25612_ (.A0(\systolic_inst.acc_wires[2][24] ),
    .A1(\C_out[88] ),
    .S(_11297_),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _25613_ (.A0(\systolic_inst.acc_wires[2][25] ),
    .A1(\C_out[89] ),
    .S(_11297_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _25614_ (.A0(\systolic_inst.acc_wires[2][26] ),
    .A1(\C_out[90] ),
    .S(_11297_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _25615_ (.A0(\systolic_inst.acc_wires[2][27] ),
    .A1(\C_out[91] ),
    .S(_11297_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _25616_ (.A0(\systolic_inst.acc_wires[2][28] ),
    .A1(\C_out[92] ),
    .S(_11297_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _25617_ (.A0(\systolic_inst.acc_wires[2][29] ),
    .A1(\C_out[93] ),
    .S(_11297_),
    .X(_02919_));
 sky130_fd_sc_hd__mux2_1 _25618_ (.A0(\systolic_inst.acc_wires[2][30] ),
    .A1(\C_out[94] ),
    .S(_11297_),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_1 _25619_ (.A0(\systolic_inst.acc_wires[2][31] ),
    .A1(\C_out[95] ),
    .S(_11297_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _25620_ (.A0(\systolic_inst.acc_wires[3][0] ),
    .A1(\C_out[96] ),
    .S(_11297_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _25621_ (.A0(\systolic_inst.acc_wires[3][1] ),
    .A1(\C_out[97] ),
    .S(_11297_),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _25622_ (.A0(\systolic_inst.acc_wires[3][2] ),
    .A1(\C_out[98] ),
    .S(_11297_),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_1 _25623_ (.A0(\systolic_inst.acc_wires[3][3] ),
    .A1(\C_out[99] ),
    .S(_11297_),
    .X(_02925_));
 sky130_fd_sc_hd__mux2_1 _25624_ (.A0(\systolic_inst.acc_wires[3][4] ),
    .A1(\C_out[100] ),
    .S(_11297_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _25625_ (.A0(\systolic_inst.acc_wires[3][5] ),
    .A1(\C_out[101] ),
    .S(_11297_),
    .X(_02927_));
 sky130_fd_sc_hd__mux2_1 _25626_ (.A0(\systolic_inst.acc_wires[3][6] ),
    .A1(\C_out[102] ),
    .S(_11297_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_1 _25627_ (.A0(\systolic_inst.acc_wires[3][7] ),
    .A1(\C_out[103] ),
    .S(_11297_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_1 _25628_ (.A0(\systolic_inst.acc_wires[3][8] ),
    .A1(\C_out[104] ),
    .S(_11297_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _25629_ (.A0(\systolic_inst.acc_wires[3][9] ),
    .A1(\C_out[105] ),
    .S(_11297_),
    .X(_02931_));
 sky130_fd_sc_hd__mux2_1 _25630_ (.A0(\systolic_inst.acc_wires[3][10] ),
    .A1(\C_out[106] ),
    .S(_11297_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _25631_ (.A0(\systolic_inst.acc_wires[3][11] ),
    .A1(\C_out[107] ),
    .S(_11297_),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_1 _25632_ (.A0(\systolic_inst.acc_wires[3][12] ),
    .A1(\C_out[108] ),
    .S(_11297_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_1 _25633_ (.A0(\systolic_inst.acc_wires[3][13] ),
    .A1(\C_out[109] ),
    .S(_11297_),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_1 _25634_ (.A0(\systolic_inst.acc_wires[3][14] ),
    .A1(\C_out[110] ),
    .S(_11297_),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_1 _25635_ (.A0(\systolic_inst.acc_wires[3][15] ),
    .A1(\C_out[111] ),
    .S(_11297_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _25636_ (.A0(\systolic_inst.acc_wires[3][16] ),
    .A1(\C_out[112] ),
    .S(_11297_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _25637_ (.A0(\systolic_inst.acc_wires[3][17] ),
    .A1(\C_out[113] ),
    .S(_11297_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _25638_ (.A0(\systolic_inst.acc_wires[3][18] ),
    .A1(\C_out[114] ),
    .S(_11297_),
    .X(_02940_));
 sky130_fd_sc_hd__mux2_1 _25639_ (.A0(\systolic_inst.acc_wires[3][19] ),
    .A1(\C_out[115] ),
    .S(_11297_),
    .X(_02941_));
 sky130_fd_sc_hd__mux2_1 _25640_ (.A0(\systolic_inst.acc_wires[3][20] ),
    .A1(\C_out[116] ),
    .S(_11297_),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_1 _25641_ (.A0(\systolic_inst.acc_wires[3][21] ),
    .A1(\C_out[117] ),
    .S(_11297_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _25642_ (.A0(\systolic_inst.acc_wires[3][22] ),
    .A1(\C_out[118] ),
    .S(_11297_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _25643_ (.A0(\systolic_inst.acc_wires[3][23] ),
    .A1(\C_out[119] ),
    .S(_11297_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_1 _25644_ (.A0(\systolic_inst.acc_wires[3][24] ),
    .A1(\C_out[120] ),
    .S(_11297_),
    .X(_02946_));
 sky130_fd_sc_hd__mux2_1 _25645_ (.A0(\systolic_inst.acc_wires[3][25] ),
    .A1(\C_out[121] ),
    .S(_11297_),
    .X(_02947_));
 sky130_fd_sc_hd__mux2_1 _25646_ (.A0(\systolic_inst.acc_wires[3][26] ),
    .A1(\C_out[122] ),
    .S(_11297_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _25647_ (.A0(\systolic_inst.acc_wires[3][27] ),
    .A1(\C_out[123] ),
    .S(_11297_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _25648_ (.A0(\systolic_inst.acc_wires[3][28] ),
    .A1(\C_out[124] ),
    .S(_11297_),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_1 _25649_ (.A0(\systolic_inst.acc_wires[3][29] ),
    .A1(\C_out[125] ),
    .S(_11297_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _25650_ (.A0(\systolic_inst.acc_wires[3][30] ),
    .A1(\C_out[126] ),
    .S(_11297_),
    .X(_02952_));
 sky130_fd_sc_hd__mux2_1 _25651_ (.A0(\systolic_inst.acc_wires[3][31] ),
    .A1(\C_out[127] ),
    .S(_11297_),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_1 _25652_ (.A0(\systolic_inst.acc_wires[4][0] ),
    .A1(\C_out[128] ),
    .S(_11297_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _25653_ (.A0(\systolic_inst.acc_wires[4][1] ),
    .A1(\C_out[129] ),
    .S(_11297_),
    .X(_02955_));
 sky130_fd_sc_hd__mux2_1 _25654_ (.A0(\systolic_inst.acc_wires[4][2] ),
    .A1(\C_out[130] ),
    .S(_11297_),
    .X(_02956_));
 sky130_fd_sc_hd__mux2_1 _25655_ (.A0(\systolic_inst.acc_wires[4][3] ),
    .A1(\C_out[131] ),
    .S(_11297_),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_1 _25656_ (.A0(\systolic_inst.acc_wires[4][4] ),
    .A1(\C_out[132] ),
    .S(_11297_),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _25657_ (.A0(\systolic_inst.acc_wires[4][5] ),
    .A1(\C_out[133] ),
    .S(_11297_),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_1 _25658_ (.A0(\systolic_inst.acc_wires[4][6] ),
    .A1(\C_out[134] ),
    .S(_11297_),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _25659_ (.A0(\systolic_inst.acc_wires[4][7] ),
    .A1(\C_out[135] ),
    .S(_11297_),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _25660_ (.A0(\systolic_inst.acc_wires[4][8] ),
    .A1(\C_out[136] ),
    .S(_11297_),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _25661_ (.A0(\systolic_inst.acc_wires[4][9] ),
    .A1(\C_out[137] ),
    .S(_11297_),
    .X(_02963_));
 sky130_fd_sc_hd__mux2_1 _25662_ (.A0(\systolic_inst.acc_wires[4][10] ),
    .A1(\C_out[138] ),
    .S(_11297_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _25663_ (.A0(\systolic_inst.acc_wires[4][11] ),
    .A1(\C_out[139] ),
    .S(_11297_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _25664_ (.A0(\systolic_inst.acc_wires[4][12] ),
    .A1(\C_out[140] ),
    .S(_11297_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_1 _25665_ (.A0(\systolic_inst.acc_wires[4][13] ),
    .A1(\C_out[141] ),
    .S(_11297_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _25666_ (.A0(\systolic_inst.acc_wires[4][14] ),
    .A1(\C_out[142] ),
    .S(_11297_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _25667_ (.A0(\systolic_inst.acc_wires[4][15] ),
    .A1(\C_out[143] ),
    .S(_11297_),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _25668_ (.A0(\systolic_inst.acc_wires[4][16] ),
    .A1(\C_out[144] ),
    .S(_11297_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _25669_ (.A0(\systolic_inst.acc_wires[4][17] ),
    .A1(\C_out[145] ),
    .S(_11297_),
    .X(_02971_));
 sky130_fd_sc_hd__mux2_1 _25670_ (.A0(\systolic_inst.acc_wires[4][18] ),
    .A1(\C_out[146] ),
    .S(_11297_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _25671_ (.A0(\systolic_inst.acc_wires[4][19] ),
    .A1(\C_out[147] ),
    .S(_11297_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _25672_ (.A0(\systolic_inst.acc_wires[4][20] ),
    .A1(\C_out[148] ),
    .S(_11297_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_1 _25673_ (.A0(\systolic_inst.acc_wires[4][21] ),
    .A1(\C_out[149] ),
    .S(_11297_),
    .X(_02975_));
 sky130_fd_sc_hd__mux2_1 _25674_ (.A0(\systolic_inst.acc_wires[4][22] ),
    .A1(\C_out[150] ),
    .S(_11297_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _25675_ (.A0(\systolic_inst.acc_wires[4][23] ),
    .A1(\C_out[151] ),
    .S(_11297_),
    .X(_02977_));
 sky130_fd_sc_hd__mux2_1 _25676_ (.A0(\systolic_inst.acc_wires[4][24] ),
    .A1(\C_out[152] ),
    .S(_11297_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_1 _25677_ (.A0(\systolic_inst.acc_wires[4][25] ),
    .A1(\C_out[153] ),
    .S(_11297_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _25678_ (.A0(\systolic_inst.acc_wires[4][26] ),
    .A1(\C_out[154] ),
    .S(_11297_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _25679_ (.A0(\systolic_inst.acc_wires[4][27] ),
    .A1(\C_out[155] ),
    .S(_11297_),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_1 _25680_ (.A0(\systolic_inst.acc_wires[4][28] ),
    .A1(\C_out[156] ),
    .S(_11297_),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_1 _25681_ (.A0(\systolic_inst.acc_wires[4][29] ),
    .A1(\C_out[157] ),
    .S(_11297_),
    .X(_02983_));
 sky130_fd_sc_hd__mux2_1 _25682_ (.A0(\systolic_inst.acc_wires[4][30] ),
    .A1(\C_out[158] ),
    .S(_11297_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _25683_ (.A0(\systolic_inst.acc_wires[4][31] ),
    .A1(\C_out[159] ),
    .S(_11297_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_1 _25684_ (.A0(\systolic_inst.acc_wires[5][0] ),
    .A1(\C_out[160] ),
    .S(_11297_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _25685_ (.A0(\systolic_inst.acc_wires[5][1] ),
    .A1(\C_out[161] ),
    .S(_11297_),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_1 _25686_ (.A0(\systolic_inst.acc_wires[5][2] ),
    .A1(\C_out[162] ),
    .S(_11297_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _25687_ (.A0(\systolic_inst.acc_wires[5][3] ),
    .A1(\C_out[163] ),
    .S(_11297_),
    .X(_02989_));
 sky130_fd_sc_hd__mux2_1 _25688_ (.A0(\systolic_inst.acc_wires[5][4] ),
    .A1(\C_out[164] ),
    .S(_11297_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _25689_ (.A0(\systolic_inst.acc_wires[5][5] ),
    .A1(\C_out[165] ),
    .S(_11297_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _25690_ (.A0(\systolic_inst.acc_wires[5][6] ),
    .A1(\C_out[166] ),
    .S(_11297_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_1 _25691_ (.A0(\systolic_inst.acc_wires[5][7] ),
    .A1(\C_out[167] ),
    .S(_11297_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_1 _25692_ (.A0(\systolic_inst.acc_wires[5][8] ),
    .A1(\C_out[168] ),
    .S(_11297_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _25693_ (.A0(\systolic_inst.acc_wires[5][9] ),
    .A1(\C_out[169] ),
    .S(_11297_),
    .X(_02995_));
 sky130_fd_sc_hd__mux2_1 _25694_ (.A0(\systolic_inst.acc_wires[5][10] ),
    .A1(\C_out[170] ),
    .S(_11297_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_1 _25695_ (.A0(\systolic_inst.acc_wires[5][11] ),
    .A1(\C_out[171] ),
    .S(_11297_),
    .X(_02997_));
 sky130_fd_sc_hd__mux2_1 _25696_ (.A0(\systolic_inst.acc_wires[5][12] ),
    .A1(\C_out[172] ),
    .S(_11297_),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_1 _25697_ (.A0(\systolic_inst.acc_wires[5][13] ),
    .A1(\C_out[173] ),
    .S(_11297_),
    .X(_02999_));
 sky130_fd_sc_hd__mux2_1 _25698_ (.A0(\systolic_inst.acc_wires[5][14] ),
    .A1(\C_out[174] ),
    .S(_11297_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _25699_ (.A0(\systolic_inst.acc_wires[5][15] ),
    .A1(\C_out[175] ),
    .S(_11297_),
    .X(_03001_));
 sky130_fd_sc_hd__mux2_1 _25700_ (.A0(\systolic_inst.acc_wires[5][16] ),
    .A1(\C_out[176] ),
    .S(_11297_),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_1 _25701_ (.A0(\systolic_inst.acc_wires[5][17] ),
    .A1(\C_out[177] ),
    .S(_11297_),
    .X(_03003_));
 sky130_fd_sc_hd__mux2_1 _25702_ (.A0(\systolic_inst.acc_wires[5][18] ),
    .A1(\C_out[178] ),
    .S(_11297_),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_1 _25703_ (.A0(\systolic_inst.acc_wires[5][19] ),
    .A1(\C_out[179] ),
    .S(_11297_),
    .X(_03005_));
 sky130_fd_sc_hd__mux2_1 _25704_ (.A0(\systolic_inst.acc_wires[5][20] ),
    .A1(\C_out[180] ),
    .S(_11297_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _25705_ (.A0(\systolic_inst.acc_wires[5][21] ),
    .A1(\C_out[181] ),
    .S(_11297_),
    .X(_03007_));
 sky130_fd_sc_hd__mux2_1 _25706_ (.A0(\systolic_inst.acc_wires[5][22] ),
    .A1(\C_out[182] ),
    .S(_11297_),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_1 _25707_ (.A0(\systolic_inst.acc_wires[5][23] ),
    .A1(\C_out[183] ),
    .S(_11297_),
    .X(_03009_));
 sky130_fd_sc_hd__mux2_1 _25708_ (.A0(\systolic_inst.acc_wires[5][24] ),
    .A1(\C_out[184] ),
    .S(_11297_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_1 _25709_ (.A0(\systolic_inst.acc_wires[5][25] ),
    .A1(\C_out[185] ),
    .S(_11297_),
    .X(_03011_));
 sky130_fd_sc_hd__mux2_1 _25710_ (.A0(\systolic_inst.acc_wires[5][26] ),
    .A1(\C_out[186] ),
    .S(_11297_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_1 _25711_ (.A0(\systolic_inst.acc_wires[5][27] ),
    .A1(\C_out[187] ),
    .S(_11297_),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_1 _25712_ (.A0(\systolic_inst.acc_wires[5][28] ),
    .A1(\C_out[188] ),
    .S(_11297_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _25713_ (.A0(\systolic_inst.acc_wires[5][29] ),
    .A1(\C_out[189] ),
    .S(_11297_),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _25714_ (.A0(\systolic_inst.acc_wires[5][30] ),
    .A1(\C_out[190] ),
    .S(_11297_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _25715_ (.A0(\systolic_inst.acc_wires[5][31] ),
    .A1(\C_out[191] ),
    .S(_11297_),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_1 _25716_ (.A0(\systolic_inst.acc_wires[6][0] ),
    .A1(\C_out[192] ),
    .S(_11297_),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_1 _25717_ (.A0(\systolic_inst.acc_wires[6][1] ),
    .A1(\C_out[193] ),
    .S(_11297_),
    .X(_03019_));
 sky130_fd_sc_hd__mux2_1 _25718_ (.A0(\systolic_inst.acc_wires[6][2] ),
    .A1(\C_out[194] ),
    .S(_11297_),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_1 _25719_ (.A0(\systolic_inst.acc_wires[6][3] ),
    .A1(\C_out[195] ),
    .S(_11297_),
    .X(_03021_));
 sky130_fd_sc_hd__mux2_1 _25720_ (.A0(\systolic_inst.acc_wires[6][4] ),
    .A1(\C_out[196] ),
    .S(_11297_),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_1 _25721_ (.A0(\systolic_inst.acc_wires[6][5] ),
    .A1(\C_out[197] ),
    .S(_11297_),
    .X(_03023_));
 sky130_fd_sc_hd__mux2_1 _25722_ (.A0(\systolic_inst.acc_wires[6][6] ),
    .A1(\C_out[198] ),
    .S(_11297_),
    .X(_03024_));
 sky130_fd_sc_hd__mux2_1 _25723_ (.A0(\systolic_inst.acc_wires[6][7] ),
    .A1(\C_out[199] ),
    .S(_11297_),
    .X(_03025_));
 sky130_fd_sc_hd__mux2_1 _25724_ (.A0(\systolic_inst.acc_wires[6][8] ),
    .A1(\C_out[200] ),
    .S(_11297_),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_1 _25725_ (.A0(\systolic_inst.acc_wires[6][9] ),
    .A1(\C_out[201] ),
    .S(_11297_),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _25726_ (.A0(\systolic_inst.acc_wires[6][10] ),
    .A1(\C_out[202] ),
    .S(_11297_),
    .X(_03028_));
 sky130_fd_sc_hd__mux2_1 _25727_ (.A0(\systolic_inst.acc_wires[6][11] ),
    .A1(\C_out[203] ),
    .S(_11297_),
    .X(_03029_));
 sky130_fd_sc_hd__mux2_1 _25728_ (.A0(\systolic_inst.acc_wires[6][12] ),
    .A1(\C_out[204] ),
    .S(_11297_),
    .X(_03030_));
 sky130_fd_sc_hd__mux2_1 _25729_ (.A0(\systolic_inst.acc_wires[6][13] ),
    .A1(\C_out[205] ),
    .S(_11297_),
    .X(_03031_));
 sky130_fd_sc_hd__mux2_1 _25730_ (.A0(\systolic_inst.acc_wires[6][14] ),
    .A1(\C_out[206] ),
    .S(_11297_),
    .X(_03032_));
 sky130_fd_sc_hd__mux2_1 _25731_ (.A0(\systolic_inst.acc_wires[6][15] ),
    .A1(\C_out[207] ),
    .S(_11297_),
    .X(_03033_));
 sky130_fd_sc_hd__mux2_1 _25732_ (.A0(\systolic_inst.acc_wires[6][16] ),
    .A1(\C_out[208] ),
    .S(_11297_),
    .X(_03034_));
 sky130_fd_sc_hd__mux2_1 _25733_ (.A0(\systolic_inst.acc_wires[6][17] ),
    .A1(\C_out[209] ),
    .S(_11297_),
    .X(_03035_));
 sky130_fd_sc_hd__mux2_1 _25734_ (.A0(\systolic_inst.acc_wires[6][18] ),
    .A1(\C_out[210] ),
    .S(_11297_),
    .X(_03036_));
 sky130_fd_sc_hd__mux2_1 _25735_ (.A0(\systolic_inst.acc_wires[6][19] ),
    .A1(\C_out[211] ),
    .S(_11297_),
    .X(_03037_));
 sky130_fd_sc_hd__mux2_1 _25736_ (.A0(\systolic_inst.acc_wires[6][20] ),
    .A1(\C_out[212] ),
    .S(_11297_),
    .X(_03038_));
 sky130_fd_sc_hd__mux2_1 _25737_ (.A0(\systolic_inst.acc_wires[6][21] ),
    .A1(\C_out[213] ),
    .S(_11297_),
    .X(_03039_));
 sky130_fd_sc_hd__mux2_1 _25738_ (.A0(\systolic_inst.acc_wires[6][22] ),
    .A1(\C_out[214] ),
    .S(_11297_),
    .X(_03040_));
 sky130_fd_sc_hd__mux2_1 _25739_ (.A0(\systolic_inst.acc_wires[6][23] ),
    .A1(\C_out[215] ),
    .S(_11297_),
    .X(_03041_));
 sky130_fd_sc_hd__mux2_1 _25740_ (.A0(\systolic_inst.acc_wires[6][24] ),
    .A1(\C_out[216] ),
    .S(_11297_),
    .X(_03042_));
 sky130_fd_sc_hd__mux2_1 _25741_ (.A0(\systolic_inst.acc_wires[6][25] ),
    .A1(\C_out[217] ),
    .S(_11297_),
    .X(_03043_));
 sky130_fd_sc_hd__mux2_1 _25742_ (.A0(\systolic_inst.acc_wires[6][26] ),
    .A1(\C_out[218] ),
    .S(_11297_),
    .X(_03044_));
 sky130_fd_sc_hd__mux2_1 _25743_ (.A0(\systolic_inst.acc_wires[6][27] ),
    .A1(\C_out[219] ),
    .S(_11297_),
    .X(_03045_));
 sky130_fd_sc_hd__mux2_1 _25744_ (.A0(\systolic_inst.acc_wires[6][28] ),
    .A1(\C_out[220] ),
    .S(_11297_),
    .X(_03046_));
 sky130_fd_sc_hd__mux2_1 _25745_ (.A0(\systolic_inst.acc_wires[6][29] ),
    .A1(\C_out[221] ),
    .S(_11297_),
    .X(_03047_));
 sky130_fd_sc_hd__mux2_1 _25746_ (.A0(\systolic_inst.acc_wires[6][30] ),
    .A1(\C_out[222] ),
    .S(_11297_),
    .X(_03048_));
 sky130_fd_sc_hd__mux2_1 _25747_ (.A0(\systolic_inst.acc_wires[6][31] ),
    .A1(\C_out[223] ),
    .S(_11297_),
    .X(_03049_));
 sky130_fd_sc_hd__mux2_1 _25748_ (.A0(\systolic_inst.acc_wires[7][0] ),
    .A1(\C_out[224] ),
    .S(_11297_),
    .X(_03050_));
 sky130_fd_sc_hd__mux2_1 _25749_ (.A0(\systolic_inst.acc_wires[7][1] ),
    .A1(\C_out[225] ),
    .S(_11297_),
    .X(_03051_));
 sky130_fd_sc_hd__mux2_1 _25750_ (.A0(\systolic_inst.acc_wires[7][2] ),
    .A1(\C_out[226] ),
    .S(_11297_),
    .X(_03052_));
 sky130_fd_sc_hd__mux2_1 _25751_ (.A0(\systolic_inst.acc_wires[7][3] ),
    .A1(\C_out[227] ),
    .S(_11297_),
    .X(_03053_));
 sky130_fd_sc_hd__mux2_1 _25752_ (.A0(\systolic_inst.acc_wires[7][4] ),
    .A1(\C_out[228] ),
    .S(_11297_),
    .X(_03054_));
 sky130_fd_sc_hd__mux2_1 _25753_ (.A0(\systolic_inst.acc_wires[7][5] ),
    .A1(\C_out[229] ),
    .S(_11297_),
    .X(_03055_));
 sky130_fd_sc_hd__mux2_1 _25754_ (.A0(\systolic_inst.acc_wires[7][6] ),
    .A1(\C_out[230] ),
    .S(_11297_),
    .X(_03056_));
 sky130_fd_sc_hd__mux2_1 _25755_ (.A0(\systolic_inst.acc_wires[7][7] ),
    .A1(\C_out[231] ),
    .S(_11297_),
    .X(_03057_));
 sky130_fd_sc_hd__mux2_1 _25756_ (.A0(\systolic_inst.acc_wires[7][8] ),
    .A1(\C_out[232] ),
    .S(_11297_),
    .X(_03058_));
 sky130_fd_sc_hd__mux2_1 _25757_ (.A0(\systolic_inst.acc_wires[7][9] ),
    .A1(\C_out[233] ),
    .S(_11297_),
    .X(_03059_));
 sky130_fd_sc_hd__mux2_1 _25758_ (.A0(\systolic_inst.acc_wires[7][10] ),
    .A1(\C_out[234] ),
    .S(_11297_),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_1 _25759_ (.A0(\systolic_inst.acc_wires[7][11] ),
    .A1(\C_out[235] ),
    .S(_11297_),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_1 _25760_ (.A0(\systolic_inst.acc_wires[7][12] ),
    .A1(\C_out[236] ),
    .S(_11297_),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_1 _25761_ (.A0(\systolic_inst.acc_wires[7][13] ),
    .A1(\C_out[237] ),
    .S(_11297_),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_1 _25762_ (.A0(\systolic_inst.acc_wires[7][14] ),
    .A1(\C_out[238] ),
    .S(_11297_),
    .X(_03064_));
 sky130_fd_sc_hd__mux2_1 _25763_ (.A0(\systolic_inst.acc_wires[7][15] ),
    .A1(\C_out[239] ),
    .S(_11297_),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_1 _25764_ (.A0(\systolic_inst.acc_wires[7][16] ),
    .A1(\C_out[240] ),
    .S(_11297_),
    .X(_03066_));
 sky130_fd_sc_hd__mux2_1 _25765_ (.A0(\systolic_inst.acc_wires[7][17] ),
    .A1(\C_out[241] ),
    .S(_11297_),
    .X(_03067_));
 sky130_fd_sc_hd__mux2_1 _25766_ (.A0(\systolic_inst.acc_wires[7][18] ),
    .A1(\C_out[242] ),
    .S(_11297_),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_1 _25767_ (.A0(\systolic_inst.acc_wires[7][19] ),
    .A1(\C_out[243] ),
    .S(_11297_),
    .X(_03069_));
 sky130_fd_sc_hd__mux2_1 _25768_ (.A0(\systolic_inst.acc_wires[7][20] ),
    .A1(\C_out[244] ),
    .S(_11297_),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _25769_ (.A0(\systolic_inst.acc_wires[7][21] ),
    .A1(\C_out[245] ),
    .S(_11297_),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_1 _25770_ (.A0(\systolic_inst.acc_wires[7][22] ),
    .A1(\C_out[246] ),
    .S(_11297_),
    .X(_03072_));
 sky130_fd_sc_hd__mux2_1 _25771_ (.A0(\systolic_inst.acc_wires[7][23] ),
    .A1(\C_out[247] ),
    .S(_11297_),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_1 _25772_ (.A0(\systolic_inst.acc_wires[7][24] ),
    .A1(\C_out[248] ),
    .S(_11297_),
    .X(_03074_));
 sky130_fd_sc_hd__mux2_1 _25773_ (.A0(\systolic_inst.acc_wires[7][25] ),
    .A1(\C_out[249] ),
    .S(_11297_),
    .X(_03075_));
 sky130_fd_sc_hd__mux2_1 _25774_ (.A0(\systolic_inst.acc_wires[7][26] ),
    .A1(\C_out[250] ),
    .S(_11297_),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_1 _25775_ (.A0(\systolic_inst.acc_wires[7][27] ),
    .A1(\C_out[251] ),
    .S(_11297_),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_1 _25776_ (.A0(\systolic_inst.acc_wires[7][28] ),
    .A1(\C_out[252] ),
    .S(_11297_),
    .X(_03078_));
 sky130_fd_sc_hd__mux2_1 _25777_ (.A0(\systolic_inst.acc_wires[7][29] ),
    .A1(\C_out[253] ),
    .S(_11297_),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_1 _25778_ (.A0(\systolic_inst.acc_wires[7][30] ),
    .A1(\C_out[254] ),
    .S(_11297_),
    .X(_03080_));
 sky130_fd_sc_hd__mux2_1 _25779_ (.A0(\systolic_inst.acc_wires[7][31] ),
    .A1(\C_out[255] ),
    .S(_11297_),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_1 _25780_ (.A0(\systolic_inst.acc_wires[8][0] ),
    .A1(\C_out[256] ),
    .S(_11297_),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_1 _25781_ (.A0(\systolic_inst.acc_wires[8][1] ),
    .A1(\C_out[257] ),
    .S(_11297_),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_1 _25782_ (.A0(\systolic_inst.acc_wires[8][2] ),
    .A1(\C_out[258] ),
    .S(_11297_),
    .X(_03084_));
 sky130_fd_sc_hd__mux2_1 _25783_ (.A0(\systolic_inst.acc_wires[8][3] ),
    .A1(\C_out[259] ),
    .S(_11297_),
    .X(_03085_));
 sky130_fd_sc_hd__mux2_1 _25784_ (.A0(\systolic_inst.acc_wires[8][4] ),
    .A1(\C_out[260] ),
    .S(_11297_),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_1 _25785_ (.A0(\systolic_inst.acc_wires[8][5] ),
    .A1(\C_out[261] ),
    .S(_11297_),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_1 _25786_ (.A0(\systolic_inst.acc_wires[8][6] ),
    .A1(\C_out[262] ),
    .S(_11297_),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_1 _25787_ (.A0(\systolic_inst.acc_wires[8][7] ),
    .A1(\C_out[263] ),
    .S(_11297_),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_1 _25788_ (.A0(\systolic_inst.acc_wires[8][8] ),
    .A1(\C_out[264] ),
    .S(_11297_),
    .X(_03090_));
 sky130_fd_sc_hd__mux2_1 _25789_ (.A0(\systolic_inst.acc_wires[8][9] ),
    .A1(\C_out[265] ),
    .S(_11297_),
    .X(_03091_));
 sky130_fd_sc_hd__mux2_1 _25790_ (.A0(\systolic_inst.acc_wires[8][10] ),
    .A1(\C_out[266] ),
    .S(_11297_),
    .X(_03092_));
 sky130_fd_sc_hd__mux2_1 _25791_ (.A0(\systolic_inst.acc_wires[8][11] ),
    .A1(\C_out[267] ),
    .S(_11297_),
    .X(_03093_));
 sky130_fd_sc_hd__mux2_1 _25792_ (.A0(\systolic_inst.acc_wires[8][12] ),
    .A1(\C_out[268] ),
    .S(_11297_),
    .X(_03094_));
 sky130_fd_sc_hd__mux2_1 _25793_ (.A0(\systolic_inst.acc_wires[8][13] ),
    .A1(\C_out[269] ),
    .S(_11297_),
    .X(_03095_));
 sky130_fd_sc_hd__mux2_1 _25794_ (.A0(\systolic_inst.acc_wires[8][14] ),
    .A1(\C_out[270] ),
    .S(_11297_),
    .X(_03096_));
 sky130_fd_sc_hd__mux2_1 _25795_ (.A0(\systolic_inst.acc_wires[8][15] ),
    .A1(\C_out[271] ),
    .S(_11297_),
    .X(_03097_));
 sky130_fd_sc_hd__mux2_1 _25796_ (.A0(\systolic_inst.acc_wires[8][16] ),
    .A1(\C_out[272] ),
    .S(_11297_),
    .X(_03098_));
 sky130_fd_sc_hd__mux2_1 _25797_ (.A0(\systolic_inst.acc_wires[8][17] ),
    .A1(\C_out[273] ),
    .S(_11297_),
    .X(_03099_));
 sky130_fd_sc_hd__mux2_1 _25798_ (.A0(\systolic_inst.acc_wires[8][18] ),
    .A1(\C_out[274] ),
    .S(_11297_),
    .X(_03100_));
 sky130_fd_sc_hd__mux2_1 _25799_ (.A0(\systolic_inst.acc_wires[8][19] ),
    .A1(\C_out[275] ),
    .S(_11297_),
    .X(_03101_));
 sky130_fd_sc_hd__mux2_1 _25800_ (.A0(\systolic_inst.acc_wires[8][20] ),
    .A1(\C_out[276] ),
    .S(_11297_),
    .X(_03102_));
 sky130_fd_sc_hd__mux2_1 _25801_ (.A0(\systolic_inst.acc_wires[8][21] ),
    .A1(\C_out[277] ),
    .S(_11297_),
    .X(_03103_));
 sky130_fd_sc_hd__mux2_1 _25802_ (.A0(\systolic_inst.acc_wires[8][22] ),
    .A1(\C_out[278] ),
    .S(_11297_),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _25803_ (.A0(\systolic_inst.acc_wires[8][23] ),
    .A1(\C_out[279] ),
    .S(_11297_),
    .X(_03105_));
 sky130_fd_sc_hd__mux2_1 _25804_ (.A0(\systolic_inst.acc_wires[8][24] ),
    .A1(\C_out[280] ),
    .S(_11297_),
    .X(_03106_));
 sky130_fd_sc_hd__mux2_1 _25805_ (.A0(\systolic_inst.acc_wires[8][25] ),
    .A1(\C_out[281] ),
    .S(_11297_),
    .X(_03107_));
 sky130_fd_sc_hd__mux2_1 _25806_ (.A0(\systolic_inst.acc_wires[8][26] ),
    .A1(\C_out[282] ),
    .S(_11297_),
    .X(_03108_));
 sky130_fd_sc_hd__mux2_1 _25807_ (.A0(\systolic_inst.acc_wires[8][27] ),
    .A1(\C_out[283] ),
    .S(_11297_),
    .X(_03109_));
 sky130_fd_sc_hd__mux2_1 _25808_ (.A0(\systolic_inst.acc_wires[8][28] ),
    .A1(\C_out[284] ),
    .S(_11297_),
    .X(_03110_));
 sky130_fd_sc_hd__mux2_1 _25809_ (.A0(\systolic_inst.acc_wires[8][29] ),
    .A1(\C_out[285] ),
    .S(_11297_),
    .X(_03111_));
 sky130_fd_sc_hd__mux2_1 _25810_ (.A0(\systolic_inst.acc_wires[8][30] ),
    .A1(\C_out[286] ),
    .S(_11297_),
    .X(_03112_));
 sky130_fd_sc_hd__mux2_1 _25811_ (.A0(\systolic_inst.acc_wires[8][31] ),
    .A1(\C_out[287] ),
    .S(_11297_),
    .X(_03113_));
 sky130_fd_sc_hd__mux2_1 _25812_ (.A0(\systolic_inst.acc_wires[9][0] ),
    .A1(\C_out[288] ),
    .S(_11297_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_1 _25813_ (.A0(\systolic_inst.acc_wires[9][1] ),
    .A1(\C_out[289] ),
    .S(_11297_),
    .X(_03115_));
 sky130_fd_sc_hd__mux2_1 _25814_ (.A0(\systolic_inst.acc_wires[9][2] ),
    .A1(\C_out[290] ),
    .S(_11297_),
    .X(_03116_));
 sky130_fd_sc_hd__mux2_1 _25815_ (.A0(\systolic_inst.acc_wires[9][3] ),
    .A1(\C_out[291] ),
    .S(_11297_),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_1 _25816_ (.A0(\systolic_inst.acc_wires[9][4] ),
    .A1(\C_out[292] ),
    .S(_11297_),
    .X(_03118_));
 sky130_fd_sc_hd__mux2_1 _25817_ (.A0(\systolic_inst.acc_wires[9][5] ),
    .A1(\C_out[293] ),
    .S(_11297_),
    .X(_03119_));
 sky130_fd_sc_hd__mux2_1 _25818_ (.A0(\systolic_inst.acc_wires[9][6] ),
    .A1(\C_out[294] ),
    .S(_11297_),
    .X(_03120_));
 sky130_fd_sc_hd__mux2_1 _25819_ (.A0(\systolic_inst.acc_wires[9][7] ),
    .A1(\C_out[295] ),
    .S(_11297_),
    .X(_03121_));
 sky130_fd_sc_hd__mux2_1 _25820_ (.A0(\systolic_inst.acc_wires[9][8] ),
    .A1(\C_out[296] ),
    .S(_11297_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_1 _25821_ (.A0(\systolic_inst.acc_wires[9][9] ),
    .A1(\C_out[297] ),
    .S(_11297_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_1 _25822_ (.A0(\systolic_inst.acc_wires[9][10] ),
    .A1(\C_out[298] ),
    .S(_11297_),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_1 _25823_ (.A0(\systolic_inst.acc_wires[9][11] ),
    .A1(\C_out[299] ),
    .S(_11297_),
    .X(_03125_));
 sky130_fd_sc_hd__mux2_1 _25824_ (.A0(\systolic_inst.acc_wires[9][12] ),
    .A1(\C_out[300] ),
    .S(_11297_),
    .X(_03126_));
 sky130_fd_sc_hd__mux2_1 _25825_ (.A0(\systolic_inst.acc_wires[9][13] ),
    .A1(\C_out[301] ),
    .S(_11297_),
    .X(_03127_));
 sky130_fd_sc_hd__mux2_1 _25826_ (.A0(\systolic_inst.acc_wires[9][14] ),
    .A1(\C_out[302] ),
    .S(_11297_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_1 _25827_ (.A0(\systolic_inst.acc_wires[9][15] ),
    .A1(\C_out[303] ),
    .S(_11297_),
    .X(_03129_));
 sky130_fd_sc_hd__mux2_1 _25828_ (.A0(\systolic_inst.acc_wires[9][16] ),
    .A1(\C_out[304] ),
    .S(_11297_),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_1 _25829_ (.A0(\systolic_inst.acc_wires[9][17] ),
    .A1(\C_out[305] ),
    .S(_11297_),
    .X(_03131_));
 sky130_fd_sc_hd__mux2_1 _25830_ (.A0(\systolic_inst.acc_wires[9][18] ),
    .A1(\C_out[306] ),
    .S(_11297_),
    .X(_03132_));
 sky130_fd_sc_hd__mux2_1 _25831_ (.A0(\systolic_inst.acc_wires[9][19] ),
    .A1(\C_out[307] ),
    .S(_11297_),
    .X(_03133_));
 sky130_fd_sc_hd__mux2_1 _25832_ (.A0(\systolic_inst.acc_wires[9][20] ),
    .A1(\C_out[308] ),
    .S(_11297_),
    .X(_03134_));
 sky130_fd_sc_hd__mux2_1 _25833_ (.A0(\systolic_inst.acc_wires[9][21] ),
    .A1(\C_out[309] ),
    .S(_11297_),
    .X(_03135_));
 sky130_fd_sc_hd__mux2_1 _25834_ (.A0(\systolic_inst.acc_wires[9][22] ),
    .A1(\C_out[310] ),
    .S(_11297_),
    .X(_03136_));
 sky130_fd_sc_hd__mux2_1 _25835_ (.A0(\systolic_inst.acc_wires[9][23] ),
    .A1(\C_out[311] ),
    .S(_11297_),
    .X(_03137_));
 sky130_fd_sc_hd__mux2_1 _25836_ (.A0(\systolic_inst.acc_wires[9][24] ),
    .A1(\C_out[312] ),
    .S(_11297_),
    .X(_03138_));
 sky130_fd_sc_hd__mux2_1 _25837_ (.A0(\systolic_inst.acc_wires[9][25] ),
    .A1(\C_out[313] ),
    .S(_11297_),
    .X(_03139_));
 sky130_fd_sc_hd__mux2_1 _25838_ (.A0(\systolic_inst.acc_wires[9][26] ),
    .A1(\C_out[314] ),
    .S(_11297_),
    .X(_03140_));
 sky130_fd_sc_hd__mux2_1 _25839_ (.A0(\systolic_inst.acc_wires[9][27] ),
    .A1(\C_out[315] ),
    .S(_11297_),
    .X(_03141_));
 sky130_fd_sc_hd__mux2_1 _25840_ (.A0(\systolic_inst.acc_wires[9][28] ),
    .A1(\C_out[316] ),
    .S(_11297_),
    .X(_03142_));
 sky130_fd_sc_hd__mux2_1 _25841_ (.A0(\systolic_inst.acc_wires[9][29] ),
    .A1(\C_out[317] ),
    .S(_11297_),
    .X(_03143_));
 sky130_fd_sc_hd__mux2_1 _25842_ (.A0(\systolic_inst.acc_wires[9][30] ),
    .A1(\C_out[318] ),
    .S(_11297_),
    .X(_03144_));
 sky130_fd_sc_hd__mux2_1 _25843_ (.A0(\systolic_inst.acc_wires[9][31] ),
    .A1(\C_out[319] ),
    .S(_11297_),
    .X(_03145_));
 sky130_fd_sc_hd__mux2_1 _25844_ (.A0(\systolic_inst.acc_wires[10][0] ),
    .A1(\C_out[320] ),
    .S(_11297_),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_1 _25845_ (.A0(\systolic_inst.acc_wires[10][1] ),
    .A1(\C_out[321] ),
    .S(_11297_),
    .X(_03147_));
 sky130_fd_sc_hd__mux2_1 _25846_ (.A0(\systolic_inst.acc_wires[10][2] ),
    .A1(\C_out[322] ),
    .S(_11297_),
    .X(_03148_));
 sky130_fd_sc_hd__mux2_1 _25847_ (.A0(\systolic_inst.acc_wires[10][3] ),
    .A1(\C_out[323] ),
    .S(_11297_),
    .X(_03149_));
 sky130_fd_sc_hd__mux2_1 _25848_ (.A0(\systolic_inst.acc_wires[10][4] ),
    .A1(\C_out[324] ),
    .S(_11297_),
    .X(_03150_));
 sky130_fd_sc_hd__mux2_1 _25849_ (.A0(\systolic_inst.acc_wires[10][5] ),
    .A1(\C_out[325] ),
    .S(_11297_),
    .X(_03151_));
 sky130_fd_sc_hd__mux2_1 _25850_ (.A0(\systolic_inst.acc_wires[10][6] ),
    .A1(\C_out[326] ),
    .S(_11297_),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_1 _25851_ (.A0(\systolic_inst.acc_wires[10][7] ),
    .A1(\C_out[327] ),
    .S(_11297_),
    .X(_03153_));
 sky130_fd_sc_hd__mux2_1 _25852_ (.A0(\systolic_inst.acc_wires[10][8] ),
    .A1(\C_out[328] ),
    .S(_11297_),
    .X(_03154_));
 sky130_fd_sc_hd__mux2_1 _25853_ (.A0(\systolic_inst.acc_wires[10][9] ),
    .A1(\C_out[329] ),
    .S(_11297_),
    .X(_03155_));
 sky130_fd_sc_hd__mux2_1 _25854_ (.A0(\systolic_inst.acc_wires[10][10] ),
    .A1(\C_out[330] ),
    .S(_11297_),
    .X(_03156_));
 sky130_fd_sc_hd__mux2_1 _25855_ (.A0(\systolic_inst.acc_wires[10][11] ),
    .A1(\C_out[331] ),
    .S(_11297_),
    .X(_03157_));
 sky130_fd_sc_hd__mux2_1 _25856_ (.A0(\systolic_inst.acc_wires[10][12] ),
    .A1(\C_out[332] ),
    .S(_11297_),
    .X(_03158_));
 sky130_fd_sc_hd__mux2_1 _25857_ (.A0(\systolic_inst.acc_wires[10][13] ),
    .A1(\C_out[333] ),
    .S(_11297_),
    .X(_03159_));
 sky130_fd_sc_hd__mux2_1 _25858_ (.A0(\systolic_inst.acc_wires[10][14] ),
    .A1(\C_out[334] ),
    .S(_11297_),
    .X(_03160_));
 sky130_fd_sc_hd__mux2_1 _25859_ (.A0(\systolic_inst.acc_wires[10][15] ),
    .A1(\C_out[335] ),
    .S(_11297_),
    .X(_03161_));
 sky130_fd_sc_hd__mux2_1 _25860_ (.A0(\systolic_inst.acc_wires[10][16] ),
    .A1(\C_out[336] ),
    .S(_11297_),
    .X(_03162_));
 sky130_fd_sc_hd__mux2_1 _25861_ (.A0(\systolic_inst.acc_wires[10][17] ),
    .A1(\C_out[337] ),
    .S(_11297_),
    .X(_03163_));
 sky130_fd_sc_hd__mux2_1 _25862_ (.A0(\systolic_inst.acc_wires[10][18] ),
    .A1(\C_out[338] ),
    .S(_11297_),
    .X(_03164_));
 sky130_fd_sc_hd__mux2_1 _25863_ (.A0(\systolic_inst.acc_wires[10][19] ),
    .A1(\C_out[339] ),
    .S(_11297_),
    .X(_03165_));
 sky130_fd_sc_hd__mux2_1 _25864_ (.A0(\systolic_inst.acc_wires[10][20] ),
    .A1(\C_out[340] ),
    .S(_11297_),
    .X(_03166_));
 sky130_fd_sc_hd__mux2_1 _25865_ (.A0(\systolic_inst.acc_wires[10][21] ),
    .A1(\C_out[341] ),
    .S(_11297_),
    .X(_03167_));
 sky130_fd_sc_hd__mux2_1 _25866_ (.A0(\systolic_inst.acc_wires[10][22] ),
    .A1(\C_out[342] ),
    .S(_11297_),
    .X(_03168_));
 sky130_fd_sc_hd__mux2_1 _25867_ (.A0(\systolic_inst.acc_wires[10][23] ),
    .A1(\C_out[343] ),
    .S(_11297_),
    .X(_03169_));
 sky130_fd_sc_hd__mux2_1 _25868_ (.A0(\systolic_inst.acc_wires[10][24] ),
    .A1(\C_out[344] ),
    .S(_11297_),
    .X(_03170_));
 sky130_fd_sc_hd__mux2_1 _25869_ (.A0(\systolic_inst.acc_wires[10][25] ),
    .A1(\C_out[345] ),
    .S(_11297_),
    .X(_03171_));
 sky130_fd_sc_hd__mux2_1 _25870_ (.A0(\systolic_inst.acc_wires[10][26] ),
    .A1(\C_out[346] ),
    .S(_11297_),
    .X(_03172_));
 sky130_fd_sc_hd__mux2_1 _25871_ (.A0(\systolic_inst.acc_wires[10][27] ),
    .A1(\C_out[347] ),
    .S(_11297_),
    .X(_03173_));
 sky130_fd_sc_hd__mux2_1 _25872_ (.A0(\systolic_inst.acc_wires[10][28] ),
    .A1(\C_out[348] ),
    .S(_11297_),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_1 _25873_ (.A0(\systolic_inst.acc_wires[10][29] ),
    .A1(\C_out[349] ),
    .S(_11297_),
    .X(_03175_));
 sky130_fd_sc_hd__mux2_1 _25874_ (.A0(\systolic_inst.acc_wires[10][30] ),
    .A1(\C_out[350] ),
    .S(_11297_),
    .X(_03176_));
 sky130_fd_sc_hd__mux2_1 _25875_ (.A0(\systolic_inst.acc_wires[10][31] ),
    .A1(\C_out[351] ),
    .S(_11297_),
    .X(_03177_));
 sky130_fd_sc_hd__mux2_1 _25876_ (.A0(\systolic_inst.acc_wires[11][0] ),
    .A1(\C_out[352] ),
    .S(_11297_),
    .X(_03178_));
 sky130_fd_sc_hd__mux2_1 _25877_ (.A0(\systolic_inst.acc_wires[11][1] ),
    .A1(\C_out[353] ),
    .S(_11297_),
    .X(_03179_));
 sky130_fd_sc_hd__mux2_1 _25878_ (.A0(\systolic_inst.acc_wires[11][2] ),
    .A1(\C_out[354] ),
    .S(_11297_),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_1 _25879_ (.A0(\systolic_inst.acc_wires[11][3] ),
    .A1(\C_out[355] ),
    .S(_11297_),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_1 _25880_ (.A0(\systolic_inst.acc_wires[11][4] ),
    .A1(\C_out[356] ),
    .S(_11297_),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_1 _25881_ (.A0(\systolic_inst.acc_wires[11][5] ),
    .A1(\C_out[357] ),
    .S(_11297_),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_1 _25882_ (.A0(\systolic_inst.acc_wires[11][6] ),
    .A1(\C_out[358] ),
    .S(_11297_),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_1 _25883_ (.A0(\systolic_inst.acc_wires[11][7] ),
    .A1(\C_out[359] ),
    .S(_11297_),
    .X(_03185_));
 sky130_fd_sc_hd__mux2_1 _25884_ (.A0(\systolic_inst.acc_wires[11][8] ),
    .A1(\C_out[360] ),
    .S(_11297_),
    .X(_03186_));
 sky130_fd_sc_hd__mux2_1 _25885_ (.A0(\systolic_inst.acc_wires[11][9] ),
    .A1(\C_out[361] ),
    .S(_11297_),
    .X(_03187_));
 sky130_fd_sc_hd__mux2_1 _25886_ (.A0(\systolic_inst.acc_wires[11][10] ),
    .A1(\C_out[362] ),
    .S(_11297_),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_1 _25887_ (.A0(\systolic_inst.acc_wires[11][11] ),
    .A1(\C_out[363] ),
    .S(_11297_),
    .X(_03189_));
 sky130_fd_sc_hd__mux2_1 _25888_ (.A0(\systolic_inst.acc_wires[11][12] ),
    .A1(\C_out[364] ),
    .S(_11297_),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_1 _25889_ (.A0(\systolic_inst.acc_wires[11][13] ),
    .A1(\C_out[365] ),
    .S(_11297_),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_1 _25890_ (.A0(\systolic_inst.acc_wires[11][14] ),
    .A1(\C_out[366] ),
    .S(_11297_),
    .X(_03192_));
 sky130_fd_sc_hd__mux2_1 _25891_ (.A0(\systolic_inst.acc_wires[11][15] ),
    .A1(\C_out[367] ),
    .S(_11297_),
    .X(_03193_));
 sky130_fd_sc_hd__mux2_1 _25892_ (.A0(\systolic_inst.acc_wires[11][16] ),
    .A1(\C_out[368] ),
    .S(_11297_),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_1 _25893_ (.A0(\systolic_inst.acc_wires[11][17] ),
    .A1(\C_out[369] ),
    .S(_11297_),
    .X(_03195_));
 sky130_fd_sc_hd__mux2_1 _25894_ (.A0(\systolic_inst.acc_wires[11][18] ),
    .A1(\C_out[370] ),
    .S(_11297_),
    .X(_03196_));
 sky130_fd_sc_hd__mux2_1 _25895_ (.A0(\systolic_inst.acc_wires[11][19] ),
    .A1(\C_out[371] ),
    .S(_11297_),
    .X(_03197_));
 sky130_fd_sc_hd__mux2_1 _25896_ (.A0(\systolic_inst.acc_wires[11][20] ),
    .A1(\C_out[372] ),
    .S(_11297_),
    .X(_03198_));
 sky130_fd_sc_hd__mux2_1 _25897_ (.A0(\systolic_inst.acc_wires[11][21] ),
    .A1(\C_out[373] ),
    .S(_11297_),
    .X(_03199_));
 sky130_fd_sc_hd__mux2_1 _25898_ (.A0(\systolic_inst.acc_wires[11][22] ),
    .A1(\C_out[374] ),
    .S(_11297_),
    .X(_03200_));
 sky130_fd_sc_hd__mux2_1 _25899_ (.A0(\systolic_inst.acc_wires[11][23] ),
    .A1(\C_out[375] ),
    .S(_11297_),
    .X(_03201_));
 sky130_fd_sc_hd__mux2_1 _25900_ (.A0(\systolic_inst.acc_wires[11][24] ),
    .A1(\C_out[376] ),
    .S(_11297_),
    .X(_03202_));
 sky130_fd_sc_hd__mux2_1 _25901_ (.A0(\systolic_inst.acc_wires[11][25] ),
    .A1(\C_out[377] ),
    .S(_11297_),
    .X(_03203_));
 sky130_fd_sc_hd__mux2_1 _25902_ (.A0(\systolic_inst.acc_wires[11][26] ),
    .A1(\C_out[378] ),
    .S(_11297_),
    .X(_03204_));
 sky130_fd_sc_hd__mux2_1 _25903_ (.A0(\systolic_inst.acc_wires[11][27] ),
    .A1(\C_out[379] ),
    .S(_11297_),
    .X(_03205_));
 sky130_fd_sc_hd__mux2_1 _25904_ (.A0(\systolic_inst.acc_wires[11][28] ),
    .A1(\C_out[380] ),
    .S(_11297_),
    .X(_03206_));
 sky130_fd_sc_hd__mux2_1 _25905_ (.A0(\systolic_inst.acc_wires[11][29] ),
    .A1(\C_out[381] ),
    .S(_11297_),
    .X(_03207_));
 sky130_fd_sc_hd__mux2_1 _25906_ (.A0(\systolic_inst.acc_wires[11][30] ),
    .A1(\C_out[382] ),
    .S(_11297_),
    .X(_03208_));
 sky130_fd_sc_hd__mux2_1 _25907_ (.A0(\systolic_inst.acc_wires[11][31] ),
    .A1(\C_out[383] ),
    .S(_11297_),
    .X(_03209_));
 sky130_fd_sc_hd__mux2_1 _25908_ (.A0(\systolic_inst.acc_wires[12][0] ),
    .A1(\C_out[384] ),
    .S(_11297_),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_1 _25909_ (.A0(\systolic_inst.acc_wires[12][1] ),
    .A1(\C_out[385] ),
    .S(_11297_),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_1 _25910_ (.A0(\systolic_inst.acc_wires[12][2] ),
    .A1(\C_out[386] ),
    .S(_11297_),
    .X(_03212_));
 sky130_fd_sc_hd__mux2_1 _25911_ (.A0(\systolic_inst.acc_wires[12][3] ),
    .A1(\C_out[387] ),
    .S(_11297_),
    .X(_03213_));
 sky130_fd_sc_hd__mux2_1 _25912_ (.A0(\systolic_inst.acc_wires[12][4] ),
    .A1(\C_out[388] ),
    .S(_11297_),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_1 _25913_ (.A0(\systolic_inst.acc_wires[12][5] ),
    .A1(\C_out[389] ),
    .S(_11297_),
    .X(_03215_));
 sky130_fd_sc_hd__mux2_1 _25914_ (.A0(\systolic_inst.acc_wires[12][6] ),
    .A1(\C_out[390] ),
    .S(_11297_),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_1 _25915_ (.A0(\systolic_inst.acc_wires[12][7] ),
    .A1(\C_out[391] ),
    .S(_11297_),
    .X(_03217_));
 sky130_fd_sc_hd__mux2_1 _25916_ (.A0(\systolic_inst.acc_wires[12][8] ),
    .A1(\C_out[392] ),
    .S(_11297_),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_1 _25917_ (.A0(\systolic_inst.acc_wires[12][9] ),
    .A1(\C_out[393] ),
    .S(_11297_),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_1 _25918_ (.A0(\systolic_inst.acc_wires[12][10] ),
    .A1(\C_out[394] ),
    .S(_11297_),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_1 _25919_ (.A0(\systolic_inst.acc_wires[12][11] ),
    .A1(\C_out[395] ),
    .S(_11297_),
    .X(_03221_));
 sky130_fd_sc_hd__mux2_1 _25920_ (.A0(\systolic_inst.acc_wires[12][12] ),
    .A1(\C_out[396] ),
    .S(_11297_),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_1 _25921_ (.A0(\systolic_inst.acc_wires[12][13] ),
    .A1(\C_out[397] ),
    .S(_11297_),
    .X(_03223_));
 sky130_fd_sc_hd__mux2_1 _25922_ (.A0(\systolic_inst.acc_wires[12][14] ),
    .A1(\C_out[398] ),
    .S(_11297_),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_1 _25923_ (.A0(\systolic_inst.acc_wires[12][15] ),
    .A1(\C_out[399] ),
    .S(_11297_),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_1 _25924_ (.A0(\systolic_inst.acc_wires[12][16] ),
    .A1(\C_out[400] ),
    .S(_11297_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_1 _25925_ (.A0(\systolic_inst.acc_wires[12][17] ),
    .A1(\C_out[401] ),
    .S(_11297_),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_1 _25926_ (.A0(\systolic_inst.acc_wires[12][18] ),
    .A1(\C_out[402] ),
    .S(_11297_),
    .X(_03228_));
 sky130_fd_sc_hd__mux2_1 _25927_ (.A0(\systolic_inst.acc_wires[12][19] ),
    .A1(\C_out[403] ),
    .S(_11297_),
    .X(_03229_));
 sky130_fd_sc_hd__mux2_1 _25928_ (.A0(\systolic_inst.acc_wires[12][20] ),
    .A1(\C_out[404] ),
    .S(_11297_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _25929_ (.A0(\systolic_inst.acc_wires[12][21] ),
    .A1(\C_out[405] ),
    .S(_11297_),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_1 _25930_ (.A0(\systolic_inst.acc_wires[12][22] ),
    .A1(\C_out[406] ),
    .S(_11297_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _25931_ (.A0(\systolic_inst.acc_wires[12][23] ),
    .A1(\C_out[407] ),
    .S(_11297_),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_1 _25932_ (.A0(\systolic_inst.acc_wires[12][24] ),
    .A1(\C_out[408] ),
    .S(_11297_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _25933_ (.A0(\systolic_inst.acc_wires[12][25] ),
    .A1(\C_out[409] ),
    .S(_11297_),
    .X(_03235_));
 sky130_fd_sc_hd__mux2_1 _25934_ (.A0(\systolic_inst.acc_wires[12][26] ),
    .A1(\C_out[410] ),
    .S(_11297_),
    .X(_03236_));
 sky130_fd_sc_hd__mux2_1 _25935_ (.A0(\systolic_inst.acc_wires[12][27] ),
    .A1(\C_out[411] ),
    .S(_11297_),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_1 _25936_ (.A0(\systolic_inst.acc_wires[12][28] ),
    .A1(\C_out[412] ),
    .S(_11297_),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_1 _25937_ (.A0(\systolic_inst.acc_wires[12][29] ),
    .A1(\C_out[413] ),
    .S(_11297_),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_1 _25938_ (.A0(\systolic_inst.acc_wires[12][30] ),
    .A1(\C_out[414] ),
    .S(_11297_),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_1 _25939_ (.A0(\systolic_inst.acc_wires[12][31] ),
    .A1(\C_out[415] ),
    .S(_11297_),
    .X(_03241_));
 sky130_fd_sc_hd__mux2_1 _25940_ (.A0(\systolic_inst.acc_wires[13][0] ),
    .A1(\C_out[416] ),
    .S(_11297_),
    .X(_03242_));
 sky130_fd_sc_hd__mux2_1 _25941_ (.A0(\systolic_inst.acc_wires[13][1] ),
    .A1(\C_out[417] ),
    .S(_11297_),
    .X(_03243_));
 sky130_fd_sc_hd__mux2_1 _25942_ (.A0(\systolic_inst.acc_wires[13][2] ),
    .A1(\C_out[418] ),
    .S(_11297_),
    .X(_03244_));
 sky130_fd_sc_hd__mux2_1 _25943_ (.A0(\systolic_inst.acc_wires[13][3] ),
    .A1(\C_out[419] ),
    .S(_11297_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_1 _25944_ (.A0(\systolic_inst.acc_wires[13][4] ),
    .A1(\C_out[420] ),
    .S(_11297_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _25945_ (.A0(\systolic_inst.acc_wires[13][5] ),
    .A1(\C_out[421] ),
    .S(_11297_),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_1 _25946_ (.A0(\systolic_inst.acc_wires[13][6] ),
    .A1(\C_out[422] ),
    .S(_11297_),
    .X(_03248_));
 sky130_fd_sc_hd__mux2_1 _25947_ (.A0(\systolic_inst.acc_wires[13][7] ),
    .A1(\C_out[423] ),
    .S(_11297_),
    .X(_03249_));
 sky130_fd_sc_hd__mux2_1 _25948_ (.A0(\systolic_inst.acc_wires[13][8] ),
    .A1(\C_out[424] ),
    .S(_11297_),
    .X(_03250_));
 sky130_fd_sc_hd__mux2_1 _25949_ (.A0(\systolic_inst.acc_wires[13][9] ),
    .A1(\C_out[425] ),
    .S(_11297_),
    .X(_03251_));
 sky130_fd_sc_hd__mux2_1 _25950_ (.A0(\systolic_inst.acc_wires[13][10] ),
    .A1(\C_out[426] ),
    .S(_11297_),
    .X(_03252_));
 sky130_fd_sc_hd__mux2_1 _25951_ (.A0(\systolic_inst.acc_wires[13][11] ),
    .A1(\C_out[427] ),
    .S(_11297_),
    .X(_03253_));
 sky130_fd_sc_hd__mux2_1 _25952_ (.A0(\systolic_inst.acc_wires[13][12] ),
    .A1(\C_out[428] ),
    .S(_11297_),
    .X(_03254_));
 sky130_fd_sc_hd__mux2_1 _25953_ (.A0(\systolic_inst.acc_wires[13][13] ),
    .A1(\C_out[429] ),
    .S(_11297_),
    .X(_03255_));
 sky130_fd_sc_hd__mux2_1 _25954_ (.A0(\systolic_inst.acc_wires[13][14] ),
    .A1(\C_out[430] ),
    .S(_11297_),
    .X(_03256_));
 sky130_fd_sc_hd__mux2_1 _25955_ (.A0(\systolic_inst.acc_wires[13][15] ),
    .A1(\C_out[431] ),
    .S(_11297_),
    .X(_03257_));
 sky130_fd_sc_hd__mux2_1 _25956_ (.A0(\systolic_inst.acc_wires[13][16] ),
    .A1(\C_out[432] ),
    .S(_11297_),
    .X(_03258_));
 sky130_fd_sc_hd__mux2_1 _25957_ (.A0(\systolic_inst.acc_wires[13][17] ),
    .A1(\C_out[433] ),
    .S(_11297_),
    .X(_03259_));
 sky130_fd_sc_hd__mux2_1 _25958_ (.A0(\systolic_inst.acc_wires[13][18] ),
    .A1(\C_out[434] ),
    .S(_11297_),
    .X(_03260_));
 sky130_fd_sc_hd__mux2_1 _25959_ (.A0(\systolic_inst.acc_wires[13][19] ),
    .A1(\C_out[435] ),
    .S(_11297_),
    .X(_03261_));
 sky130_fd_sc_hd__mux2_1 _25960_ (.A0(\systolic_inst.acc_wires[13][20] ),
    .A1(\C_out[436] ),
    .S(_11297_),
    .X(_03262_));
 sky130_fd_sc_hd__mux2_1 _25961_ (.A0(\systolic_inst.acc_wires[13][21] ),
    .A1(\C_out[437] ),
    .S(_11297_),
    .X(_03263_));
 sky130_fd_sc_hd__mux2_1 _25962_ (.A0(\systolic_inst.acc_wires[13][22] ),
    .A1(\C_out[438] ),
    .S(_11297_),
    .X(_03264_));
 sky130_fd_sc_hd__mux2_1 _25963_ (.A0(\systolic_inst.acc_wires[13][23] ),
    .A1(\C_out[439] ),
    .S(_11297_),
    .X(_03265_));
 sky130_fd_sc_hd__mux2_1 _25964_ (.A0(\systolic_inst.acc_wires[13][24] ),
    .A1(\ser_C.parallel_data[440] ),
    .S(_11297_),
    .X(_03266_));
 sky130_fd_sc_hd__mux2_1 _25965_ (.A0(\systolic_inst.acc_wires[13][25] ),
    .A1(\ser_C.parallel_data[441] ),
    .S(_11297_),
    .X(_03267_));
 sky130_fd_sc_hd__mux2_1 _25966_ (.A0(\systolic_inst.acc_wires[13][26] ),
    .A1(\ser_C.parallel_data[442] ),
    .S(_11297_),
    .X(_03268_));
 sky130_fd_sc_hd__mux2_1 _25967_ (.A0(\systolic_inst.acc_wires[13][27] ),
    .A1(\ser_C.parallel_data[443] ),
    .S(_11297_),
    .X(_03269_));
 sky130_fd_sc_hd__mux2_1 _25968_ (.A0(\systolic_inst.acc_wires[13][28] ),
    .A1(\ser_C.parallel_data[444] ),
    .S(_11297_),
    .X(_03270_));
 sky130_fd_sc_hd__mux2_1 _25969_ (.A0(\systolic_inst.acc_wires[13][29] ),
    .A1(\ser_C.parallel_data[445] ),
    .S(_11297_),
    .X(_03271_));
 sky130_fd_sc_hd__mux2_1 _25970_ (.A0(\systolic_inst.acc_wires[13][30] ),
    .A1(\ser_C.parallel_data[446] ),
    .S(_11297_),
    .X(_03272_));
 sky130_fd_sc_hd__mux2_1 _25971_ (.A0(\systolic_inst.acc_wires[13][31] ),
    .A1(\ser_C.parallel_data[447] ),
    .S(_11297_),
    .X(_03273_));
 sky130_fd_sc_hd__mux2_1 _25972_ (.A0(\systolic_inst.acc_wires[14][0] ),
    .A1(\ser_C.parallel_data[448] ),
    .S(_11297_),
    .X(_03274_));
 sky130_fd_sc_hd__mux2_1 _25973_ (.A0(\systolic_inst.acc_wires[14][1] ),
    .A1(\ser_C.parallel_data[449] ),
    .S(_11297_),
    .X(_03275_));
 sky130_fd_sc_hd__mux2_1 _25974_ (.A0(\systolic_inst.acc_wires[14][2] ),
    .A1(\ser_C.parallel_data[450] ),
    .S(_11297_),
    .X(_03276_));
 sky130_fd_sc_hd__mux2_1 _25975_ (.A0(\systolic_inst.acc_wires[14][3] ),
    .A1(\ser_C.parallel_data[451] ),
    .S(_11297_),
    .X(_03277_));
 sky130_fd_sc_hd__mux2_1 _25976_ (.A0(\systolic_inst.acc_wires[14][4] ),
    .A1(\ser_C.parallel_data[452] ),
    .S(_11297_),
    .X(_03278_));
 sky130_fd_sc_hd__mux2_1 _25977_ (.A0(\systolic_inst.acc_wires[14][5] ),
    .A1(\ser_C.parallel_data[453] ),
    .S(_11297_),
    .X(_03279_));
 sky130_fd_sc_hd__mux2_1 _25978_ (.A0(\systolic_inst.acc_wires[14][6] ),
    .A1(\ser_C.parallel_data[454] ),
    .S(_11297_),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_1 _25979_ (.A0(\systolic_inst.acc_wires[14][7] ),
    .A1(\ser_C.parallel_data[455] ),
    .S(_11297_),
    .X(_03281_));
 sky130_fd_sc_hd__mux2_1 _25980_ (.A0(\systolic_inst.acc_wires[14][8] ),
    .A1(\ser_C.parallel_data[456] ),
    .S(_11297_),
    .X(_03282_));
 sky130_fd_sc_hd__mux2_1 _25981_ (.A0(\systolic_inst.acc_wires[14][9] ),
    .A1(\ser_C.parallel_data[457] ),
    .S(_11297_),
    .X(_03283_));
 sky130_fd_sc_hd__mux2_1 _25982_ (.A0(\systolic_inst.acc_wires[14][10] ),
    .A1(\ser_C.parallel_data[458] ),
    .S(_11297_),
    .X(_03284_));
 sky130_fd_sc_hd__mux2_1 _25983_ (.A0(\systolic_inst.acc_wires[14][11] ),
    .A1(\ser_C.parallel_data[459] ),
    .S(_11297_),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_1 _25984_ (.A0(\systolic_inst.acc_wires[14][12] ),
    .A1(\ser_C.parallel_data[460] ),
    .S(_11297_),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_1 _25985_ (.A0(\systolic_inst.acc_wires[14][13] ),
    .A1(\ser_C.parallel_data[461] ),
    .S(_11297_),
    .X(_03287_));
 sky130_fd_sc_hd__mux2_1 _25986_ (.A0(\systolic_inst.acc_wires[14][14] ),
    .A1(\ser_C.parallel_data[462] ),
    .S(_11297_),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_1 _25987_ (.A0(\systolic_inst.acc_wires[14][15] ),
    .A1(\ser_C.parallel_data[463] ),
    .S(_11297_),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_1 _25988_ (.A0(\systolic_inst.acc_wires[14][16] ),
    .A1(\ser_C.parallel_data[464] ),
    .S(_11297_),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _25989_ (.A0(\systolic_inst.acc_wires[14][17] ),
    .A1(\ser_C.parallel_data[465] ),
    .S(_11297_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _25990_ (.A0(\systolic_inst.acc_wires[14][18] ),
    .A1(\ser_C.parallel_data[466] ),
    .S(_11297_),
    .X(_03292_));
 sky130_fd_sc_hd__mux2_1 _25991_ (.A0(\systolic_inst.acc_wires[14][19] ),
    .A1(\ser_C.parallel_data[467] ),
    .S(_11297_),
    .X(_03293_));
 sky130_fd_sc_hd__mux2_1 _25992_ (.A0(\systolic_inst.acc_wires[14][20] ),
    .A1(\ser_C.parallel_data[468] ),
    .S(_11297_),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_1 _25993_ (.A0(\systolic_inst.acc_wires[14][21] ),
    .A1(\ser_C.parallel_data[469] ),
    .S(_11297_),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_1 _25994_ (.A0(\systolic_inst.acc_wires[14][22] ),
    .A1(\ser_C.parallel_data[470] ),
    .S(_11297_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _25995_ (.A0(\systolic_inst.acc_wires[14][23] ),
    .A1(\ser_C.parallel_data[471] ),
    .S(_11297_),
    .X(_03297_));
 sky130_fd_sc_hd__mux2_1 _25996_ (.A0(\systolic_inst.acc_wires[14][24] ),
    .A1(\ser_C.parallel_data[472] ),
    .S(_11297_),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_1 _25997_ (.A0(\systolic_inst.acc_wires[14][25] ),
    .A1(\ser_C.parallel_data[473] ),
    .S(_11297_),
    .X(_03299_));
 sky130_fd_sc_hd__mux2_1 _25998_ (.A0(\systolic_inst.acc_wires[14][26] ),
    .A1(\ser_C.parallel_data[474] ),
    .S(_11297_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_1 _25999_ (.A0(\systolic_inst.acc_wires[14][27] ),
    .A1(\ser_C.parallel_data[475] ),
    .S(_11297_),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_1 _26000_ (.A0(\systolic_inst.acc_wires[14][28] ),
    .A1(\ser_C.parallel_data[476] ),
    .S(_11297_),
    .X(_03302_));
 sky130_fd_sc_hd__mux2_1 _26001_ (.A0(\systolic_inst.acc_wires[14][29] ),
    .A1(\ser_C.parallel_data[477] ),
    .S(_11297_),
    .X(_03303_));
 sky130_fd_sc_hd__mux2_1 _26002_ (.A0(\systolic_inst.acc_wires[14][30] ),
    .A1(\ser_C.parallel_data[478] ),
    .S(_11297_),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_1 _26003_ (.A0(\systolic_inst.acc_wires[14][31] ),
    .A1(\ser_C.parallel_data[479] ),
    .S(_11297_),
    .X(_03305_));
 sky130_fd_sc_hd__mux2_1 _26004_ (.A0(\systolic_inst.acc_wires[15][0] ),
    .A1(\ser_C.parallel_data[480] ),
    .S(_11297_),
    .X(_03306_));
 sky130_fd_sc_hd__mux2_1 _26005_ (.A0(\systolic_inst.acc_wires[15][1] ),
    .A1(\ser_C.parallel_data[481] ),
    .S(_11297_),
    .X(_03307_));
 sky130_fd_sc_hd__mux2_1 _26006_ (.A0(\systolic_inst.acc_wires[15][2] ),
    .A1(\ser_C.parallel_data[482] ),
    .S(_11297_),
    .X(_03308_));
 sky130_fd_sc_hd__mux2_1 _26007_ (.A0(\systolic_inst.acc_wires[15][3] ),
    .A1(\ser_C.parallel_data[483] ),
    .S(_11297_),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_1 _26008_ (.A0(\systolic_inst.acc_wires[15][4] ),
    .A1(\ser_C.parallel_data[484] ),
    .S(_11297_),
    .X(_03310_));
 sky130_fd_sc_hd__mux2_1 _26009_ (.A0(\systolic_inst.acc_wires[15][5] ),
    .A1(\ser_C.parallel_data[485] ),
    .S(_11297_),
    .X(_03311_));
 sky130_fd_sc_hd__mux2_1 _26010_ (.A0(\systolic_inst.acc_wires[15][6] ),
    .A1(\ser_C.parallel_data[486] ),
    .S(_11297_),
    .X(_03312_));
 sky130_fd_sc_hd__mux2_1 _26011_ (.A0(\systolic_inst.acc_wires[15][7] ),
    .A1(\ser_C.parallel_data[487] ),
    .S(_11297_),
    .X(_03313_));
 sky130_fd_sc_hd__mux2_1 _26012_ (.A0(\systolic_inst.acc_wires[15][8] ),
    .A1(\ser_C.parallel_data[488] ),
    .S(_11297_),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_1 _26013_ (.A0(\systolic_inst.acc_wires[15][9] ),
    .A1(\ser_C.parallel_data[489] ),
    .S(_11297_),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_1 _26014_ (.A0(\systolic_inst.acc_wires[15][10] ),
    .A1(\ser_C.parallel_data[490] ),
    .S(_11297_),
    .X(_03316_));
 sky130_fd_sc_hd__mux2_1 _26015_ (.A0(\systolic_inst.acc_wires[15][11] ),
    .A1(\ser_C.parallel_data[491] ),
    .S(_11297_),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_1 _26016_ (.A0(\systolic_inst.acc_wires[15][12] ),
    .A1(\ser_C.parallel_data[492] ),
    .S(_11297_),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_1 _26017_ (.A0(\systolic_inst.acc_wires[15][13] ),
    .A1(\ser_C.parallel_data[493] ),
    .S(_11297_),
    .X(_03319_));
 sky130_fd_sc_hd__mux2_1 _26018_ (.A0(\systolic_inst.acc_wires[15][14] ),
    .A1(\ser_C.parallel_data[494] ),
    .S(_11297_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _26019_ (.A0(\systolic_inst.acc_wires[15][15] ),
    .A1(\ser_C.parallel_data[495] ),
    .S(_11297_),
    .X(_03321_));
 sky130_fd_sc_hd__mux2_1 _26020_ (.A0(\systolic_inst.acc_wires[15][16] ),
    .A1(\ser_C.parallel_data[496] ),
    .S(_11297_),
    .X(_03322_));
 sky130_fd_sc_hd__mux2_1 _26021_ (.A0(\systolic_inst.acc_wires[15][17] ),
    .A1(\ser_C.parallel_data[497] ),
    .S(_11297_),
    .X(_03323_));
 sky130_fd_sc_hd__mux2_1 _26022_ (.A0(\systolic_inst.acc_wires[15][18] ),
    .A1(\ser_C.parallel_data[498] ),
    .S(_11297_),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_1 _26023_ (.A0(\systolic_inst.acc_wires[15][19] ),
    .A1(\ser_C.parallel_data[499] ),
    .S(_11297_),
    .X(_03325_));
 sky130_fd_sc_hd__mux2_1 _26024_ (.A0(\systolic_inst.acc_wires[15][20] ),
    .A1(\ser_C.parallel_data[500] ),
    .S(_11297_),
    .X(_03326_));
 sky130_fd_sc_hd__mux2_1 _26025_ (.A0(\systolic_inst.acc_wires[15][21] ),
    .A1(\ser_C.parallel_data[501] ),
    .S(_11297_),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_1 _26026_ (.A0(\systolic_inst.acc_wires[15][22] ),
    .A1(\ser_C.parallel_data[502] ),
    .S(_11297_),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_1 _26027_ (.A0(\systolic_inst.acc_wires[15][23] ),
    .A1(\ser_C.parallel_data[503] ),
    .S(_11297_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_1 _26028_ (.A0(\systolic_inst.acc_wires[15][24] ),
    .A1(\ser_C.parallel_data[504] ),
    .S(_11297_),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_1 _26029_ (.A0(\systolic_inst.acc_wires[15][25] ),
    .A1(\ser_C.parallel_data[505] ),
    .S(_11297_),
    .X(_03331_));
 sky130_fd_sc_hd__mux2_1 _26030_ (.A0(\systolic_inst.acc_wires[15][26] ),
    .A1(\ser_C.parallel_data[506] ),
    .S(_11297_),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_1 _26031_ (.A0(\systolic_inst.acc_wires[15][27] ),
    .A1(\ser_C.parallel_data[507] ),
    .S(_11297_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _26032_ (.A0(\systolic_inst.acc_wires[15][28] ),
    .A1(\ser_C.parallel_data[508] ),
    .S(_11297_),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_1 _26033_ (.A0(\systolic_inst.acc_wires[15][29] ),
    .A1(\ser_C.parallel_data[509] ),
    .S(_11297_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _26034_ (.A0(\systolic_inst.acc_wires[15][30] ),
    .A1(\ser_C.parallel_data[510] ),
    .S(_11297_),
    .X(_03336_));
 sky130_fd_sc_hd__mux2_1 _26035_ (.A0(\systolic_inst.acc_wires[15][31] ),
    .A1(\ser_C.parallel_data[511] ),
    .S(_11297_),
    .X(_03337_));
 sky130_fd_sc_hd__mux2_1 _26036_ (.A0(\systolic_inst.B_outs[15][0] ),
    .A1(\systolic_inst.B_outs[11][0] ),
    .S(\systolic_inst.ce_local ),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_1 _26037_ (.A0(\systolic_inst.B_outs[15][1] ),
    .A1(\systolic_inst.B_outs[11][1] ),
    .S(\systolic_inst.ce_local ),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _26038_ (.A0(\systolic_inst.B_outs[15][2] ),
    .A1(\systolic_inst.B_outs[11][2] ),
    .S(\systolic_inst.ce_local ),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_1 _26039_ (.A0(\systolic_inst.B_outs[15][3] ),
    .A1(\systolic_inst.B_outs[11][3] ),
    .S(\systolic_inst.ce_local ),
    .X(_03341_));
 sky130_fd_sc_hd__mux2_1 _26040_ (.A0(\systolic_inst.B_outs[15][4] ),
    .A1(\systolic_inst.B_outs[11][4] ),
    .S(\systolic_inst.ce_local ),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_1 _26041_ (.A0(\systolic_inst.B_outs[15][5] ),
    .A1(\systolic_inst.B_outs[11][5] ),
    .S(\systolic_inst.ce_local ),
    .X(_03343_));
 sky130_fd_sc_hd__mux2_1 _26042_ (.A0(\systolic_inst.B_outs[15][6] ),
    .A1(\systolic_inst.B_outs[11][6] ),
    .S(\systolic_inst.ce_local ),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_1 _26043_ (.A0(\systolic_inst.B_outs[15][7] ),
    .A1(\systolic_inst.B_outs[11][7] ),
    .S(\systolic_inst.ce_local ),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _26044_ (.A0(C_out_serial_data),
    .A1(\ser_C.shift_reg[0] ),
    .S(C_out_frame_sync),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_1 _26045_ (.A0(\deser_B.serial_word[0] ),
    .A1(\deser_B.shift_reg[0] ),
    .S(_00001_),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_1 _26046_ (.A0(\deser_B.serial_word[1] ),
    .A1(\deser_B.shift_reg[1] ),
    .S(_00001_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _26047_ (.A0(\deser_B.serial_word[2] ),
    .A1(\deser_B.shift_reg[2] ),
    .S(_00001_),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_1 _26048_ (.A0(\deser_B.serial_word[3] ),
    .A1(\deser_B.shift_reg[3] ),
    .S(_00001_),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_1 _26049_ (.A0(\deser_B.serial_word[4] ),
    .A1(\deser_B.shift_reg[4] ),
    .S(_00001_),
    .X(_03351_));
 sky130_fd_sc_hd__mux2_1 _26050_ (.A0(\deser_B.serial_word[5] ),
    .A1(\deser_B.shift_reg[5] ),
    .S(_00001_),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_1 _26051_ (.A0(\deser_B.serial_word[6] ),
    .A1(\deser_B.shift_reg[6] ),
    .S(_00001_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_1 _26052_ (.A0(\deser_B.serial_word[7] ),
    .A1(\deser_B.shift_reg[7] ),
    .S(_00001_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_1 _26053_ (.A0(\deser_B.serial_word[8] ),
    .A1(\deser_B.shift_reg[8] ),
    .S(_00001_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _26054_ (.A0(\deser_B.serial_word[9] ),
    .A1(\deser_B.shift_reg[9] ),
    .S(_00001_),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_1 _26055_ (.A0(\deser_B.serial_word[10] ),
    .A1(\deser_B.shift_reg[10] ),
    .S(_00001_),
    .X(_03357_));
 sky130_fd_sc_hd__mux2_1 _26056_ (.A0(\deser_B.serial_word[11] ),
    .A1(\deser_B.shift_reg[11] ),
    .S(_00001_),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_1 _26057_ (.A0(\deser_B.serial_word[12] ),
    .A1(\deser_B.shift_reg[12] ),
    .S(_00001_),
    .X(_03359_));
 sky130_fd_sc_hd__mux2_1 _26058_ (.A0(\deser_B.serial_word[13] ),
    .A1(\deser_B.shift_reg[13] ),
    .S(_00001_),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_1 _26059_ (.A0(\deser_B.serial_word[14] ),
    .A1(\deser_B.shift_reg[14] ),
    .S(_00001_),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_1 _26060_ (.A0(\deser_B.serial_word[15] ),
    .A1(\deser_B.shift_reg[15] ),
    .S(_00001_),
    .X(_03362_));
 sky130_fd_sc_hd__mux2_1 _26061_ (.A0(\deser_B.serial_word[16] ),
    .A1(\deser_B.shift_reg[16] ),
    .S(_00001_),
    .X(_03363_));
 sky130_fd_sc_hd__mux2_1 _26062_ (.A0(\deser_B.serial_word[17] ),
    .A1(\deser_B.shift_reg[17] ),
    .S(_00001_),
    .X(_03364_));
 sky130_fd_sc_hd__mux2_1 _26063_ (.A0(\deser_B.serial_word[18] ),
    .A1(\deser_B.shift_reg[18] ),
    .S(_00001_),
    .X(_03365_));
 sky130_fd_sc_hd__mux2_1 _26064_ (.A0(\deser_B.serial_word[19] ),
    .A1(\deser_B.shift_reg[19] ),
    .S(_00001_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_1 _26065_ (.A0(\deser_B.serial_word[20] ),
    .A1(\deser_B.shift_reg[20] ),
    .S(_00001_),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_1 _26066_ (.A0(\deser_B.serial_word[21] ),
    .A1(\deser_B.shift_reg[21] ),
    .S(_00001_),
    .X(_03368_));
 sky130_fd_sc_hd__mux2_1 _26067_ (.A0(\deser_B.serial_word[22] ),
    .A1(\deser_B.shift_reg[22] ),
    .S(_00001_),
    .X(_03369_));
 sky130_fd_sc_hd__mux2_1 _26068_ (.A0(\deser_B.serial_word[23] ),
    .A1(\deser_B.shift_reg[23] ),
    .S(_00001_),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_1 _26069_ (.A0(\deser_B.serial_word[24] ),
    .A1(\deser_B.shift_reg[24] ),
    .S(_00001_),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_1 _26070_ (.A0(\deser_B.serial_word[25] ),
    .A1(\deser_B.shift_reg[25] ),
    .S(_00001_),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_1 _26071_ (.A0(\deser_B.serial_word[26] ),
    .A1(\deser_B.shift_reg[26] ),
    .S(_00001_),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_1 _26072_ (.A0(\deser_B.serial_word[27] ),
    .A1(\deser_B.shift_reg[27] ),
    .S(_00001_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _26073_ (.A0(\deser_B.serial_word[28] ),
    .A1(\deser_B.shift_reg[28] ),
    .S(_00001_),
    .X(_03375_));
 sky130_fd_sc_hd__mux2_1 _26074_ (.A0(\deser_B.serial_word[29] ),
    .A1(\deser_B.shift_reg[29] ),
    .S(_00001_),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_1 _26075_ (.A0(\deser_B.serial_word[30] ),
    .A1(\deser_B.shift_reg[30] ),
    .S(_00001_),
    .X(_03377_));
 sky130_fd_sc_hd__mux2_1 _26076_ (.A0(\deser_B.serial_word[31] ),
    .A1(\deser_B.shift_reg[31] ),
    .S(_00001_),
    .X(_03378_));
 sky130_fd_sc_hd__mux2_1 _26077_ (.A0(\deser_B.serial_word[32] ),
    .A1(\deser_B.shift_reg[32] ),
    .S(_00001_),
    .X(_03379_));
 sky130_fd_sc_hd__mux2_1 _26078_ (.A0(\deser_B.serial_word[33] ),
    .A1(\deser_B.shift_reg[33] ),
    .S(_00001_),
    .X(_03380_));
 sky130_fd_sc_hd__mux2_1 _26079_ (.A0(\deser_B.serial_word[34] ),
    .A1(\deser_B.shift_reg[34] ),
    .S(_00001_),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_1 _26080_ (.A0(\deser_B.serial_word[35] ),
    .A1(\deser_B.shift_reg[35] ),
    .S(_00001_),
    .X(_03382_));
 sky130_fd_sc_hd__mux2_1 _26081_ (.A0(\deser_B.serial_word[36] ),
    .A1(\deser_B.shift_reg[36] ),
    .S(_00001_),
    .X(_03383_));
 sky130_fd_sc_hd__mux2_1 _26082_ (.A0(\deser_B.serial_word[37] ),
    .A1(\deser_B.shift_reg[37] ),
    .S(_00001_),
    .X(_03384_));
 sky130_fd_sc_hd__mux2_1 _26083_ (.A0(\deser_B.serial_word[38] ),
    .A1(\deser_B.shift_reg[38] ),
    .S(_00001_),
    .X(_03385_));
 sky130_fd_sc_hd__mux2_1 _26084_ (.A0(\deser_B.serial_word[39] ),
    .A1(\deser_B.shift_reg[39] ),
    .S(_00001_),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_1 _26085_ (.A0(\deser_B.serial_word[40] ),
    .A1(\deser_B.shift_reg[40] ),
    .S(_00001_),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _26086_ (.A0(\deser_B.serial_word[41] ),
    .A1(\deser_B.shift_reg[41] ),
    .S(_00001_),
    .X(_03388_));
 sky130_fd_sc_hd__mux2_1 _26087_ (.A0(\deser_B.serial_word[42] ),
    .A1(\deser_B.shift_reg[42] ),
    .S(_00001_),
    .X(_03389_));
 sky130_fd_sc_hd__mux2_1 _26088_ (.A0(\deser_B.serial_word[43] ),
    .A1(\deser_B.shift_reg[43] ),
    .S(_00001_),
    .X(_03390_));
 sky130_fd_sc_hd__mux2_1 _26089_ (.A0(\deser_B.serial_word[44] ),
    .A1(\deser_B.shift_reg[44] ),
    .S(_00001_),
    .X(_03391_));
 sky130_fd_sc_hd__mux2_1 _26090_ (.A0(\deser_B.serial_word[45] ),
    .A1(\deser_B.shift_reg[45] ),
    .S(_00001_),
    .X(_03392_));
 sky130_fd_sc_hd__mux2_1 _26091_ (.A0(\deser_B.serial_word[46] ),
    .A1(\deser_B.shift_reg[46] ),
    .S(_00001_),
    .X(_03393_));
 sky130_fd_sc_hd__mux2_1 _26092_ (.A0(\deser_B.serial_word[47] ),
    .A1(\deser_B.shift_reg[47] ),
    .S(_00001_),
    .X(_03394_));
 sky130_fd_sc_hd__mux2_1 _26093_ (.A0(\deser_B.serial_word[48] ),
    .A1(\deser_B.shift_reg[48] ),
    .S(_00001_),
    .X(_03395_));
 sky130_fd_sc_hd__mux2_1 _26094_ (.A0(\deser_B.serial_word[49] ),
    .A1(\deser_B.shift_reg[49] ),
    .S(_00001_),
    .X(_03396_));
 sky130_fd_sc_hd__mux2_1 _26095_ (.A0(\deser_B.serial_word[50] ),
    .A1(\deser_B.shift_reg[50] ),
    .S(_00001_),
    .X(_03397_));
 sky130_fd_sc_hd__mux2_1 _26096_ (.A0(\deser_B.serial_word[51] ),
    .A1(\deser_B.shift_reg[51] ),
    .S(_00001_),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_1 _26097_ (.A0(\deser_B.serial_word[52] ),
    .A1(\deser_B.shift_reg[52] ),
    .S(_00001_),
    .X(_03399_));
 sky130_fd_sc_hd__mux2_1 _26098_ (.A0(\deser_B.serial_word[53] ),
    .A1(\deser_B.shift_reg[53] ),
    .S(_00001_),
    .X(_03400_));
 sky130_fd_sc_hd__mux2_1 _26099_ (.A0(\deser_B.serial_word[54] ),
    .A1(\deser_B.shift_reg[54] ),
    .S(_00001_),
    .X(_03401_));
 sky130_fd_sc_hd__mux2_1 _26100_ (.A0(\deser_B.serial_word[55] ),
    .A1(\deser_B.shift_reg[55] ),
    .S(_00001_),
    .X(_03402_));
 sky130_fd_sc_hd__mux2_1 _26101_ (.A0(\deser_B.serial_word[56] ),
    .A1(\deser_B.shift_reg[56] ),
    .S(_00001_),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _26102_ (.A0(\deser_B.serial_word[57] ),
    .A1(\deser_B.shift_reg[57] ),
    .S(_00001_),
    .X(_03404_));
 sky130_fd_sc_hd__mux2_1 _26103_ (.A0(\deser_B.serial_word[58] ),
    .A1(\deser_B.shift_reg[58] ),
    .S(_00001_),
    .X(_03405_));
 sky130_fd_sc_hd__mux2_1 _26104_ (.A0(\deser_B.serial_word[59] ),
    .A1(\deser_B.shift_reg[59] ),
    .S(_00001_),
    .X(_03406_));
 sky130_fd_sc_hd__mux2_1 _26105_ (.A0(\deser_B.serial_word[60] ),
    .A1(\deser_B.shift_reg[60] ),
    .S(_00001_),
    .X(_03407_));
 sky130_fd_sc_hd__mux2_1 _26106_ (.A0(\deser_B.serial_word[61] ),
    .A1(\deser_B.shift_reg[61] ),
    .S(_00001_),
    .X(_03408_));
 sky130_fd_sc_hd__mux2_1 _26107_ (.A0(\deser_B.serial_word[62] ),
    .A1(\deser_B.shift_reg[62] ),
    .S(_00001_),
    .X(_03409_));
 sky130_fd_sc_hd__mux2_1 _26108_ (.A0(\deser_B.serial_word[63] ),
    .A1(\deser_B.shift_reg[63] ),
    .S(_00001_),
    .X(_03410_));
 sky130_fd_sc_hd__mux2_1 _26109_ (.A0(\deser_B.serial_word[64] ),
    .A1(\deser_B.shift_reg[64] ),
    .S(_00001_),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_1 _26110_ (.A0(\deser_B.serial_word[65] ),
    .A1(\deser_B.shift_reg[65] ),
    .S(_00001_),
    .X(_03412_));
 sky130_fd_sc_hd__mux2_1 _26111_ (.A0(\deser_B.serial_word[66] ),
    .A1(\deser_B.shift_reg[66] ),
    .S(_00001_),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_1 _26112_ (.A0(\deser_B.serial_word[67] ),
    .A1(\deser_B.shift_reg[67] ),
    .S(_00001_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _26113_ (.A0(\deser_B.serial_word[68] ),
    .A1(\deser_B.shift_reg[68] ),
    .S(_00001_),
    .X(_03415_));
 sky130_fd_sc_hd__mux2_1 _26114_ (.A0(\deser_B.serial_word[69] ),
    .A1(\deser_B.shift_reg[69] ),
    .S(_00001_),
    .X(_03416_));
 sky130_fd_sc_hd__mux2_1 _26115_ (.A0(\deser_B.serial_word[70] ),
    .A1(\deser_B.shift_reg[70] ),
    .S(_00001_),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_1 _26116_ (.A0(\deser_B.serial_word[71] ),
    .A1(\deser_B.shift_reg[71] ),
    .S(_00001_),
    .X(_03418_));
 sky130_fd_sc_hd__mux2_1 _26117_ (.A0(\deser_B.serial_word[72] ),
    .A1(\deser_B.shift_reg[72] ),
    .S(_00001_),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_1 _26118_ (.A0(\deser_B.serial_word[73] ),
    .A1(\deser_B.shift_reg[73] ),
    .S(_00001_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _26119_ (.A0(\deser_B.serial_word[74] ),
    .A1(\deser_B.shift_reg[74] ),
    .S(_00001_),
    .X(_03421_));
 sky130_fd_sc_hd__mux2_1 _26120_ (.A0(\deser_B.serial_word[75] ),
    .A1(\deser_B.shift_reg[75] ),
    .S(_00001_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_1 _26121_ (.A0(\deser_B.serial_word[76] ),
    .A1(\deser_B.shift_reg[76] ),
    .S(_00001_),
    .X(_03423_));
 sky130_fd_sc_hd__mux2_1 _26122_ (.A0(\deser_B.serial_word[77] ),
    .A1(\deser_B.shift_reg[77] ),
    .S(_00001_),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_1 _26123_ (.A0(\deser_B.serial_word[78] ),
    .A1(\deser_B.shift_reg[78] ),
    .S(_00001_),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_1 _26124_ (.A0(\deser_B.serial_word[79] ),
    .A1(\deser_B.shift_reg[79] ),
    .S(_00001_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _26125_ (.A0(\deser_B.serial_word[80] ),
    .A1(\deser_B.shift_reg[80] ),
    .S(_00001_),
    .X(_03427_));
 sky130_fd_sc_hd__mux2_1 _26126_ (.A0(\deser_B.serial_word[81] ),
    .A1(\deser_B.shift_reg[81] ),
    .S(_00001_),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_1 _26127_ (.A0(\deser_B.serial_word[82] ),
    .A1(\deser_B.shift_reg[82] ),
    .S(_00001_),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_1 _26128_ (.A0(\deser_B.serial_word[83] ),
    .A1(\deser_B.shift_reg[83] ),
    .S(_00001_),
    .X(_03430_));
 sky130_fd_sc_hd__mux2_1 _26129_ (.A0(\deser_B.serial_word[84] ),
    .A1(\deser_B.shift_reg[84] ),
    .S(_00001_),
    .X(_03431_));
 sky130_fd_sc_hd__mux2_1 _26130_ (.A0(\deser_B.serial_word[85] ),
    .A1(\deser_B.shift_reg[85] ),
    .S(_00001_),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_1 _26131_ (.A0(\deser_B.serial_word[86] ),
    .A1(\deser_B.shift_reg[86] ),
    .S(_00001_),
    .X(_03433_));
 sky130_fd_sc_hd__mux2_1 _26132_ (.A0(\deser_B.serial_word[87] ),
    .A1(\deser_B.shift_reg[87] ),
    .S(_00001_),
    .X(_03434_));
 sky130_fd_sc_hd__mux2_1 _26133_ (.A0(\deser_B.serial_word[88] ),
    .A1(\deser_B.shift_reg[88] ),
    .S(_00001_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _26134_ (.A0(\deser_B.serial_word[89] ),
    .A1(\deser_B.shift_reg[89] ),
    .S(_00001_),
    .X(_03436_));
 sky130_fd_sc_hd__mux2_1 _26135_ (.A0(\deser_B.serial_word[90] ),
    .A1(\deser_B.shift_reg[90] ),
    .S(_00001_),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_1 _26136_ (.A0(\deser_B.serial_word[91] ),
    .A1(\deser_B.shift_reg[91] ),
    .S(_00001_),
    .X(_03438_));
 sky130_fd_sc_hd__mux2_1 _26137_ (.A0(\deser_B.serial_word[92] ),
    .A1(\deser_B.shift_reg[92] ),
    .S(_00001_),
    .X(_03439_));
 sky130_fd_sc_hd__mux2_1 _26138_ (.A0(\deser_B.serial_word[93] ),
    .A1(\deser_B.shift_reg[93] ),
    .S(_00001_),
    .X(_03440_));
 sky130_fd_sc_hd__mux2_1 _26139_ (.A0(\deser_B.serial_word[94] ),
    .A1(\deser_B.shift_reg[94] ),
    .S(_00001_),
    .X(_03441_));
 sky130_fd_sc_hd__mux2_1 _26140_ (.A0(\deser_B.serial_word[95] ),
    .A1(\deser_B.shift_reg[95] ),
    .S(_00001_),
    .X(_03442_));
 sky130_fd_sc_hd__mux2_1 _26141_ (.A0(\deser_B.serial_word[96] ),
    .A1(\deser_B.shift_reg[96] ),
    .S(_00001_),
    .X(_03443_));
 sky130_fd_sc_hd__mux2_1 _26142_ (.A0(\deser_B.serial_word[97] ),
    .A1(\deser_B.shift_reg[97] ),
    .S(_00001_),
    .X(_03444_));
 sky130_fd_sc_hd__mux2_1 _26143_ (.A0(\deser_B.serial_word[98] ),
    .A1(\deser_B.shift_reg[98] ),
    .S(_00001_),
    .X(_03445_));
 sky130_fd_sc_hd__mux2_1 _26144_ (.A0(\deser_B.serial_word[99] ),
    .A1(\deser_B.shift_reg[99] ),
    .S(_00001_),
    .X(_03446_));
 sky130_fd_sc_hd__mux2_1 _26145_ (.A0(\deser_B.serial_word[100] ),
    .A1(\deser_B.shift_reg[100] ),
    .S(_00001_),
    .X(_03447_));
 sky130_fd_sc_hd__mux2_1 _26146_ (.A0(\deser_B.serial_word[101] ),
    .A1(\deser_B.shift_reg[101] ),
    .S(_00001_),
    .X(_03448_));
 sky130_fd_sc_hd__mux2_1 _26147_ (.A0(\deser_B.serial_word[102] ),
    .A1(\deser_B.shift_reg[102] ),
    .S(_00001_),
    .X(_03449_));
 sky130_fd_sc_hd__mux2_1 _26148_ (.A0(\deser_B.serial_word[103] ),
    .A1(\deser_B.shift_reg[103] ),
    .S(_00001_),
    .X(_03450_));
 sky130_fd_sc_hd__mux2_1 _26149_ (.A0(\deser_B.serial_word[104] ),
    .A1(\deser_B.shift_reg[104] ),
    .S(_00001_),
    .X(_03451_));
 sky130_fd_sc_hd__mux2_1 _26150_ (.A0(\deser_B.serial_word[105] ),
    .A1(\deser_B.shift_reg[105] ),
    .S(_00001_),
    .X(_03452_));
 sky130_fd_sc_hd__mux2_1 _26151_ (.A0(\deser_B.serial_word[106] ),
    .A1(\deser_B.shift_reg[106] ),
    .S(_00001_),
    .X(_03453_));
 sky130_fd_sc_hd__mux2_1 _26152_ (.A0(\deser_B.serial_word[107] ),
    .A1(\deser_B.shift_reg[107] ),
    .S(_00001_),
    .X(_03454_));
 sky130_fd_sc_hd__mux2_1 _26153_ (.A0(\deser_B.serial_word[108] ),
    .A1(\deser_B.shift_reg[108] ),
    .S(_00001_),
    .X(_03455_));
 sky130_fd_sc_hd__mux2_1 _26154_ (.A0(\deser_B.serial_word[109] ),
    .A1(\deser_B.shift_reg[109] ),
    .S(_00001_),
    .X(_03456_));
 sky130_fd_sc_hd__mux2_1 _26155_ (.A0(\deser_B.serial_word[110] ),
    .A1(\deser_B.shift_reg[110] ),
    .S(_00001_),
    .X(_03457_));
 sky130_fd_sc_hd__mux2_1 _26156_ (.A0(\deser_B.serial_word[111] ),
    .A1(\deser_B.shift_reg[111] ),
    .S(_00001_),
    .X(_03458_));
 sky130_fd_sc_hd__mux2_1 _26157_ (.A0(\deser_B.serial_word[112] ),
    .A1(\deser_B.shift_reg[112] ),
    .S(_00001_),
    .X(_03459_));
 sky130_fd_sc_hd__mux2_1 _26158_ (.A0(\deser_B.serial_word[113] ),
    .A1(\deser_B.shift_reg[113] ),
    .S(_00001_),
    .X(_03460_));
 sky130_fd_sc_hd__mux2_1 _26159_ (.A0(\deser_B.serial_word[114] ),
    .A1(\deser_B.shift_reg[114] ),
    .S(_00001_),
    .X(_03461_));
 sky130_fd_sc_hd__mux2_1 _26160_ (.A0(\deser_B.serial_word[115] ),
    .A1(\deser_B.shift_reg[115] ),
    .S(_00001_),
    .X(_03462_));
 sky130_fd_sc_hd__mux2_1 _26161_ (.A0(\deser_B.serial_word[116] ),
    .A1(\deser_B.shift_reg[116] ),
    .S(_00001_),
    .X(_03463_));
 sky130_fd_sc_hd__mux2_1 _26162_ (.A0(\deser_B.serial_word[117] ),
    .A1(\deser_B.shift_reg[117] ),
    .S(_00001_),
    .X(_03464_));
 sky130_fd_sc_hd__mux2_1 _26163_ (.A0(\deser_B.serial_word[118] ),
    .A1(\deser_B.shift_reg[118] ),
    .S(_00001_),
    .X(_03465_));
 sky130_fd_sc_hd__mux2_1 _26164_ (.A0(\deser_B.serial_word[119] ),
    .A1(\deser_B.shift_reg[119] ),
    .S(_00001_),
    .X(_03466_));
 sky130_fd_sc_hd__mux2_1 _26165_ (.A0(\deser_B.serial_word[120] ),
    .A1(\deser_B.shift_reg[120] ),
    .S(_00001_),
    .X(_03467_));
 sky130_fd_sc_hd__mux2_1 _26166_ (.A0(\deser_B.serial_word[121] ),
    .A1(\deser_B.shift_reg[121] ),
    .S(_00001_),
    .X(_03468_));
 sky130_fd_sc_hd__mux2_1 _26167_ (.A0(\deser_B.serial_word[122] ),
    .A1(\deser_B.shift_reg[122] ),
    .S(_00001_),
    .X(_03469_));
 sky130_fd_sc_hd__mux2_1 _26168_ (.A0(\deser_B.serial_word[123] ),
    .A1(\deser_B.shift_reg[123] ),
    .S(_00001_),
    .X(_03470_));
 sky130_fd_sc_hd__mux2_1 _26169_ (.A0(\deser_B.serial_word[124] ),
    .A1(\deser_B.shift_reg[124] ),
    .S(_00001_),
    .X(_03471_));
 sky130_fd_sc_hd__mux2_1 _26170_ (.A0(\deser_B.serial_word[125] ),
    .A1(\deser_B.shift_reg[125] ),
    .S(_00001_),
    .X(_03472_));
 sky130_fd_sc_hd__mux2_1 _26171_ (.A0(\deser_B.serial_word[126] ),
    .A1(\deser_B.shift_reg[126] ),
    .S(_00001_),
    .X(_03473_));
 sky130_fd_sc_hd__mux2_1 _26172_ (.A0(\deser_B.serial_word[127] ),
    .A1(\deser_B.shift_reg[127] ),
    .S(_00001_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_1 _26173_ (.A0(C_out_frame_sync),
    .A1(_10643_),
    .S(\ser_C.bit_idx[0] ),
    .X(_03475_));
 sky130_fd_sc_hd__and3_2 _26174_ (.A(C_out_frame_sync),
    .B(\ser_C.bit_idx[0] ),
    .C(\ser_C.bit_idx[1] ),
    .X(_11245_));
 sky130_fd_sc_hd__a21oi_2 _26175_ (.A1(C_out_frame_sync),
    .A2(\ser_C.bit_idx[0] ),
    .B1(\ser_C.bit_idx[1] ),
    .Y(_11246_));
 sky130_fd_sc_hd__nor3_2 _26176_ (.A(_11302_),
    .B(_11245_),
    .C(_11246_),
    .Y(_03476_));
 sky130_fd_sc_hd__and2_2 _26177_ (.A(\ser_C.bit_idx[2] ),
    .B(_11245_),
    .X(_11247_));
 sky130_fd_sc_hd__o21ai_2 _26178_ (.A1(\ser_C.bit_idx[2] ),
    .A2(_11245_),
    .B1(_11303_),
    .Y(_11248_));
 sky130_fd_sc_hd__nor2_2 _26179_ (.A(_11247_),
    .B(_11248_),
    .Y(_03477_));
 sky130_fd_sc_hd__a21oi_2 _26180_ (.A1(\ser_C.bit_idx[3] ),
    .A2(_11303_),
    .B1(_11247_),
    .Y(_11249_));
 sky130_fd_sc_hd__a21oi_2 _26181_ (.A1(\ser_C.bit_idx[3] ),
    .A2(_11247_),
    .B1(_11249_),
    .Y(_03478_));
 sky130_fd_sc_hd__and3_2 _26182_ (.A(\ser_C.bit_idx[3] ),
    .B(\ser_C.bit_idx[4] ),
    .C(_11247_),
    .X(_11250_));
 sky130_fd_sc_hd__a22oi_2 _26183_ (.A1(\ser_C.bit_idx[4] ),
    .A2(_11303_),
    .B1(_11247_),
    .B2(\ser_C.bit_idx[3] ),
    .Y(_11251_));
 sky130_fd_sc_hd__nor2_2 _26184_ (.A(_11250_),
    .B(_11251_),
    .Y(_03479_));
 sky130_fd_sc_hd__and2_2 _26185_ (.A(\ser_C.bit_idx[5] ),
    .B(_11250_),
    .X(_11252_));
 sky130_fd_sc_hd__o21ai_2 _26186_ (.A1(\ser_C.bit_idx[5] ),
    .A2(_11250_),
    .B1(_11303_),
    .Y(_11253_));
 sky130_fd_sc_hd__nor2_2 _26187_ (.A(_11252_),
    .B(_11253_),
    .Y(_03480_));
 sky130_fd_sc_hd__and3_2 _26188_ (.A(\ser_C.bit_idx[5] ),
    .B(\ser_C.bit_idx[6] ),
    .C(_11250_),
    .X(_11254_));
 sky130_fd_sc_hd__nor2_2 _26189_ (.A(_11302_),
    .B(_11254_),
    .Y(_11255_));
 sky130_fd_sc_hd__mux2_1 _26190_ (.A0(_11252_),
    .A1(_11255_),
    .S(\ser_C.bit_idx[6] ),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_1 _26191_ (.A0(_11254_),
    .A1(_11255_),
    .S(\ser_C.bit_idx[7] ),
    .X(_03482_));
 sky130_fd_sc_hd__nor2_2 _26192_ (.A(\ser_C.bit_idx[8] ),
    .B(_11300_),
    .Y(_11256_));
 sky130_fd_sc_hd__a2bb2o_2 _26193_ (.A1_N(_11301_),
    .A2_N(_11256_),
    .B1(_10643_),
    .B2(\ser_C.bit_idx[8] ),
    .X(_03483_));
 sky130_fd_sc_hd__a22o_2 _26194_ (.A1(\systolic_inst.A_shift[30][0] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[120] ),
    .X(_03484_));
 sky130_fd_sc_hd__a22o_2 _26195_ (.A1(\systolic_inst.A_shift[30][1] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[121] ),
    .X(_03485_));
 sky130_fd_sc_hd__a22o_2 _26196_ (.A1(\systolic_inst.A_shift[30][2] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[122] ),
    .X(_03486_));
 sky130_fd_sc_hd__a22o_2 _26197_ (.A1(\systolic_inst.A_shift[30][3] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[123] ),
    .X(_03487_));
 sky130_fd_sc_hd__a22o_2 _26198_ (.A1(\systolic_inst.A_shift[30][4] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[124] ),
    .X(_03488_));
 sky130_fd_sc_hd__a22o_2 _26199_ (.A1(\systolic_inst.A_shift[30][5] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[125] ),
    .X(_03489_));
 sky130_fd_sc_hd__a22o_2 _26200_ (.A1(\systolic_inst.A_shift[30][6] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[126] ),
    .X(_03490_));
 sky130_fd_sc_hd__a22o_2 _26201_ (.A1(\systolic_inst.A_shift[30][7] ),
    .A2(_11332_),
    .B1(_11333_),
    .B2(\A_in[127] ),
    .X(_03491_));
 sky130_fd_sc_hd__dfrtp_2 _26202_ (.CLK(A_in_serial_clk),
    .D(_00010_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26203_ (.CLK(A_in_serial_clk),
    .D(_00011_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26204_ (.CLK(A_in_serial_clk),
    .D(_00012_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26205_ (.CLK(A_in_serial_clk),
    .D(_00013_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26206_ (.CLK(A_in_serial_clk),
    .D(_00014_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26207_ (.CLK(A_in_serial_clk),
    .D(_00015_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26208_ (.CLK(A_in_serial_clk),
    .D(_00016_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26209_ (.CLK(A_in_serial_clk),
    .D(_00017_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26210_ (.CLK(A_in_serial_clk),
    .D(_00018_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26211_ (.CLK(A_in_serial_clk),
    .D(_00019_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26212_ (.CLK(A_in_serial_clk),
    .D(_00020_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[10] ));
 sky130_fd_sc_hd__dfrtp_2 _26213_ (.CLK(A_in_serial_clk),
    .D(_00021_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26214_ (.CLK(A_in_serial_clk),
    .D(_00022_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[12] ));
 sky130_fd_sc_hd__dfrtp_2 _26215_ (.CLK(A_in_serial_clk),
    .D(_00023_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26216_ (.CLK(A_in_serial_clk),
    .D(_00024_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26217_ (.CLK(A_in_serial_clk),
    .D(_00025_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26218_ (.CLK(A_in_serial_clk),
    .D(_00026_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[16] ));
 sky130_fd_sc_hd__dfrtp_2 _26219_ (.CLK(A_in_serial_clk),
    .D(_00027_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[17] ));
 sky130_fd_sc_hd__dfrtp_2 _26220_ (.CLK(A_in_serial_clk),
    .D(_00028_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[18] ));
 sky130_fd_sc_hd__dfrtp_2 _26221_ (.CLK(A_in_serial_clk),
    .D(_00029_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[19] ));
 sky130_fd_sc_hd__dfrtp_2 _26222_ (.CLK(A_in_serial_clk),
    .D(_00030_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[20] ));
 sky130_fd_sc_hd__dfrtp_2 _26223_ (.CLK(A_in_serial_clk),
    .D(_00031_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[21] ));
 sky130_fd_sc_hd__dfrtp_2 _26224_ (.CLK(A_in_serial_clk),
    .D(_00032_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[22] ));
 sky130_fd_sc_hd__dfrtp_2 _26225_ (.CLK(A_in_serial_clk),
    .D(_00033_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[23] ));
 sky130_fd_sc_hd__dfrtp_2 _26226_ (.CLK(A_in_serial_clk),
    .D(_00034_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[24] ));
 sky130_fd_sc_hd__dfrtp_2 _26227_ (.CLK(A_in_serial_clk),
    .D(_00035_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[25] ));
 sky130_fd_sc_hd__dfrtp_2 _26228_ (.CLK(A_in_serial_clk),
    .D(_00036_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[26] ));
 sky130_fd_sc_hd__dfrtp_2 _26229_ (.CLK(A_in_serial_clk),
    .D(_00037_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[27] ));
 sky130_fd_sc_hd__dfrtp_2 _26230_ (.CLK(A_in_serial_clk),
    .D(_00038_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[28] ));
 sky130_fd_sc_hd__dfrtp_2 _26231_ (.CLK(A_in_serial_clk),
    .D(_00039_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[29] ));
 sky130_fd_sc_hd__dfrtp_2 _26232_ (.CLK(A_in_serial_clk),
    .D(_00040_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[30] ));
 sky130_fd_sc_hd__dfrtp_2 _26233_ (.CLK(A_in_serial_clk),
    .D(_00041_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[31] ));
 sky130_fd_sc_hd__dfrtp_2 _26234_ (.CLK(A_in_serial_clk),
    .D(_00042_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[32] ));
 sky130_fd_sc_hd__dfrtp_2 _26235_ (.CLK(A_in_serial_clk),
    .D(_00043_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[33] ));
 sky130_fd_sc_hd__dfrtp_2 _26236_ (.CLK(A_in_serial_clk),
    .D(_00044_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[34] ));
 sky130_fd_sc_hd__dfrtp_2 _26237_ (.CLK(A_in_serial_clk),
    .D(_00045_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[35] ));
 sky130_fd_sc_hd__dfrtp_2 _26238_ (.CLK(A_in_serial_clk),
    .D(_00046_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[36] ));
 sky130_fd_sc_hd__dfrtp_2 _26239_ (.CLK(A_in_serial_clk),
    .D(_00047_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[37] ));
 sky130_fd_sc_hd__dfrtp_2 _26240_ (.CLK(A_in_serial_clk),
    .D(_00048_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[38] ));
 sky130_fd_sc_hd__dfrtp_2 _26241_ (.CLK(A_in_serial_clk),
    .D(_00049_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[39] ));
 sky130_fd_sc_hd__dfrtp_2 _26242_ (.CLK(A_in_serial_clk),
    .D(_00050_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[40] ));
 sky130_fd_sc_hd__dfrtp_2 _26243_ (.CLK(A_in_serial_clk),
    .D(_00051_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[41] ));
 sky130_fd_sc_hd__dfrtp_2 _26244_ (.CLK(A_in_serial_clk),
    .D(_00052_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[42] ));
 sky130_fd_sc_hd__dfrtp_2 _26245_ (.CLK(A_in_serial_clk),
    .D(_00053_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[43] ));
 sky130_fd_sc_hd__dfrtp_2 _26246_ (.CLK(A_in_serial_clk),
    .D(_00054_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[44] ));
 sky130_fd_sc_hd__dfrtp_2 _26247_ (.CLK(A_in_serial_clk),
    .D(_00055_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[45] ));
 sky130_fd_sc_hd__dfrtp_2 _26248_ (.CLK(A_in_serial_clk),
    .D(_00056_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[46] ));
 sky130_fd_sc_hd__dfrtp_2 _26249_ (.CLK(A_in_serial_clk),
    .D(_00057_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[47] ));
 sky130_fd_sc_hd__dfrtp_2 _26250_ (.CLK(A_in_serial_clk),
    .D(_00058_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[48] ));
 sky130_fd_sc_hd__dfrtp_2 _26251_ (.CLK(A_in_serial_clk),
    .D(_00059_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[49] ));
 sky130_fd_sc_hd__dfrtp_2 _26252_ (.CLK(A_in_serial_clk),
    .D(_00060_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[50] ));
 sky130_fd_sc_hd__dfrtp_2 _26253_ (.CLK(A_in_serial_clk),
    .D(_00061_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[51] ));
 sky130_fd_sc_hd__dfrtp_2 _26254_ (.CLK(A_in_serial_clk),
    .D(_00062_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[52] ));
 sky130_fd_sc_hd__dfrtp_2 _26255_ (.CLK(A_in_serial_clk),
    .D(_00063_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[53] ));
 sky130_fd_sc_hd__dfrtp_2 _26256_ (.CLK(A_in_serial_clk),
    .D(_00064_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[54] ));
 sky130_fd_sc_hd__dfrtp_2 _26257_ (.CLK(A_in_serial_clk),
    .D(_00065_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[55] ));
 sky130_fd_sc_hd__dfrtp_2 _26258_ (.CLK(A_in_serial_clk),
    .D(_00066_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[56] ));
 sky130_fd_sc_hd__dfrtp_2 _26259_ (.CLK(A_in_serial_clk),
    .D(_00067_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[57] ));
 sky130_fd_sc_hd__dfrtp_2 _26260_ (.CLK(A_in_serial_clk),
    .D(_00068_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[58] ));
 sky130_fd_sc_hd__dfrtp_2 _26261_ (.CLK(A_in_serial_clk),
    .D(_00069_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[59] ));
 sky130_fd_sc_hd__dfrtp_2 _26262_ (.CLK(A_in_serial_clk),
    .D(_00070_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[60] ));
 sky130_fd_sc_hd__dfrtp_2 _26263_ (.CLK(A_in_serial_clk),
    .D(_00071_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[61] ));
 sky130_fd_sc_hd__dfrtp_2 _26264_ (.CLK(A_in_serial_clk),
    .D(_00072_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[62] ));
 sky130_fd_sc_hd__dfrtp_2 _26265_ (.CLK(A_in_serial_clk),
    .D(_00073_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[63] ));
 sky130_fd_sc_hd__dfrtp_2 _26266_ (.CLK(A_in_serial_clk),
    .D(_00074_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[64] ));
 sky130_fd_sc_hd__dfrtp_2 _26267_ (.CLK(A_in_serial_clk),
    .D(_00075_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[65] ));
 sky130_fd_sc_hd__dfrtp_2 _26268_ (.CLK(A_in_serial_clk),
    .D(_00076_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[66] ));
 sky130_fd_sc_hd__dfrtp_2 _26269_ (.CLK(A_in_serial_clk),
    .D(_00077_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[67] ));
 sky130_fd_sc_hd__dfrtp_2 _26270_ (.CLK(A_in_serial_clk),
    .D(_00078_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[68] ));
 sky130_fd_sc_hd__dfrtp_2 _26271_ (.CLK(A_in_serial_clk),
    .D(_00079_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[69] ));
 sky130_fd_sc_hd__dfrtp_2 _26272_ (.CLK(A_in_serial_clk),
    .D(_00080_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[70] ));
 sky130_fd_sc_hd__dfrtp_2 _26273_ (.CLK(A_in_serial_clk),
    .D(_00081_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[71] ));
 sky130_fd_sc_hd__dfrtp_2 _26274_ (.CLK(A_in_serial_clk),
    .D(_00082_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[72] ));
 sky130_fd_sc_hd__dfrtp_2 _26275_ (.CLK(A_in_serial_clk),
    .D(_00083_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[73] ));
 sky130_fd_sc_hd__dfrtp_2 _26276_ (.CLK(A_in_serial_clk),
    .D(_00084_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[74] ));
 sky130_fd_sc_hd__dfrtp_2 _26277_ (.CLK(A_in_serial_clk),
    .D(_00085_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[75] ));
 sky130_fd_sc_hd__dfrtp_2 _26278_ (.CLK(A_in_serial_clk),
    .D(_00086_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[76] ));
 sky130_fd_sc_hd__dfrtp_2 _26279_ (.CLK(A_in_serial_clk),
    .D(_00087_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[77] ));
 sky130_fd_sc_hd__dfrtp_2 _26280_ (.CLK(A_in_serial_clk),
    .D(_00088_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[78] ));
 sky130_fd_sc_hd__dfrtp_2 _26281_ (.CLK(A_in_serial_clk),
    .D(_00089_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[79] ));
 sky130_fd_sc_hd__dfrtp_2 _26282_ (.CLK(A_in_serial_clk),
    .D(_00090_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[80] ));
 sky130_fd_sc_hd__dfrtp_2 _26283_ (.CLK(A_in_serial_clk),
    .D(_00091_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[81] ));
 sky130_fd_sc_hd__dfrtp_2 _26284_ (.CLK(A_in_serial_clk),
    .D(_00092_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[82] ));
 sky130_fd_sc_hd__dfrtp_2 _26285_ (.CLK(A_in_serial_clk),
    .D(_00093_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[83] ));
 sky130_fd_sc_hd__dfrtp_2 _26286_ (.CLK(A_in_serial_clk),
    .D(_00094_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[84] ));
 sky130_fd_sc_hd__dfrtp_2 _26287_ (.CLK(A_in_serial_clk),
    .D(_00095_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[85] ));
 sky130_fd_sc_hd__dfrtp_2 _26288_ (.CLK(A_in_serial_clk),
    .D(_00096_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[86] ));
 sky130_fd_sc_hd__dfrtp_2 _26289_ (.CLK(A_in_serial_clk),
    .D(_00097_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[87] ));
 sky130_fd_sc_hd__dfrtp_2 _26290_ (.CLK(A_in_serial_clk),
    .D(_00098_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[88] ));
 sky130_fd_sc_hd__dfrtp_2 _26291_ (.CLK(A_in_serial_clk),
    .D(_00099_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[89] ));
 sky130_fd_sc_hd__dfrtp_2 _26292_ (.CLK(A_in_serial_clk),
    .D(_00100_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[90] ));
 sky130_fd_sc_hd__dfrtp_2 _26293_ (.CLK(A_in_serial_clk),
    .D(_00101_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[91] ));
 sky130_fd_sc_hd__dfrtp_2 _26294_ (.CLK(A_in_serial_clk),
    .D(_00102_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[92] ));
 sky130_fd_sc_hd__dfrtp_2 _26295_ (.CLK(A_in_serial_clk),
    .D(_00103_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[93] ));
 sky130_fd_sc_hd__dfrtp_2 _26296_ (.CLK(A_in_serial_clk),
    .D(_00104_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[94] ));
 sky130_fd_sc_hd__dfrtp_2 _26297_ (.CLK(A_in_serial_clk),
    .D(_00105_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[95] ));
 sky130_fd_sc_hd__dfrtp_2 _26298_ (.CLK(A_in_serial_clk),
    .D(_00106_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[96] ));
 sky130_fd_sc_hd__dfrtp_2 _26299_ (.CLK(A_in_serial_clk),
    .D(_00107_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[97] ));
 sky130_fd_sc_hd__dfrtp_2 _26300_ (.CLK(A_in_serial_clk),
    .D(_00108_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[98] ));
 sky130_fd_sc_hd__dfrtp_2 _26301_ (.CLK(A_in_serial_clk),
    .D(_00109_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[99] ));
 sky130_fd_sc_hd__dfrtp_2 _26302_ (.CLK(A_in_serial_clk),
    .D(_00110_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[100] ));
 sky130_fd_sc_hd__dfrtp_2 _26303_ (.CLK(A_in_serial_clk),
    .D(_00111_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[101] ));
 sky130_fd_sc_hd__dfrtp_2 _26304_ (.CLK(A_in_serial_clk),
    .D(_00112_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[102] ));
 sky130_fd_sc_hd__dfrtp_2 _26305_ (.CLK(A_in_serial_clk),
    .D(_00113_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[103] ));
 sky130_fd_sc_hd__dfrtp_2 _26306_ (.CLK(A_in_serial_clk),
    .D(_00114_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[104] ));
 sky130_fd_sc_hd__dfrtp_2 _26307_ (.CLK(A_in_serial_clk),
    .D(_00115_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[105] ));
 sky130_fd_sc_hd__dfrtp_2 _26308_ (.CLK(A_in_serial_clk),
    .D(_00116_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[106] ));
 sky130_fd_sc_hd__dfrtp_2 _26309_ (.CLK(A_in_serial_clk),
    .D(_00117_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[107] ));
 sky130_fd_sc_hd__dfrtp_2 _26310_ (.CLK(A_in_serial_clk),
    .D(_00118_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[108] ));
 sky130_fd_sc_hd__dfrtp_2 _26311_ (.CLK(A_in_serial_clk),
    .D(_00119_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[109] ));
 sky130_fd_sc_hd__dfrtp_2 _26312_ (.CLK(A_in_serial_clk),
    .D(_00120_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[110] ));
 sky130_fd_sc_hd__dfrtp_2 _26313_ (.CLK(A_in_serial_clk),
    .D(_00121_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[111] ));
 sky130_fd_sc_hd__dfrtp_2 _26314_ (.CLK(A_in_serial_clk),
    .D(_00122_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[112] ));
 sky130_fd_sc_hd__dfrtp_2 _26315_ (.CLK(A_in_serial_clk),
    .D(_00123_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[113] ));
 sky130_fd_sc_hd__dfrtp_2 _26316_ (.CLK(A_in_serial_clk),
    .D(_00124_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[114] ));
 sky130_fd_sc_hd__dfrtp_2 _26317_ (.CLK(A_in_serial_clk),
    .D(_00125_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[115] ));
 sky130_fd_sc_hd__dfrtp_2 _26318_ (.CLK(A_in_serial_clk),
    .D(_00126_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[116] ));
 sky130_fd_sc_hd__dfrtp_2 _26319_ (.CLK(A_in_serial_clk),
    .D(_00127_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[117] ));
 sky130_fd_sc_hd__dfrtp_2 _26320_ (.CLK(A_in_serial_clk),
    .D(_00128_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[118] ));
 sky130_fd_sc_hd__dfrtp_2 _26321_ (.CLK(A_in_serial_clk),
    .D(_00129_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[119] ));
 sky130_fd_sc_hd__dfrtp_2 _26322_ (.CLK(A_in_serial_clk),
    .D(_00130_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[120] ));
 sky130_fd_sc_hd__dfrtp_2 _26323_ (.CLK(A_in_serial_clk),
    .D(_00131_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[121] ));
 sky130_fd_sc_hd__dfrtp_2 _26324_ (.CLK(A_in_serial_clk),
    .D(_00132_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[122] ));
 sky130_fd_sc_hd__dfrtp_2 _26325_ (.CLK(A_in_serial_clk),
    .D(_00133_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[123] ));
 sky130_fd_sc_hd__dfrtp_2 _26326_ (.CLK(A_in_serial_clk),
    .D(_00134_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[124] ));
 sky130_fd_sc_hd__dfrtp_2 _26327_ (.CLK(A_in_serial_clk),
    .D(_00135_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[125] ));
 sky130_fd_sc_hd__dfrtp_2 _26328_ (.CLK(A_in_serial_clk),
    .D(_00136_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[126] ));
 sky130_fd_sc_hd__dfrtp_2 _26329_ (.CLK(A_in_serial_clk),
    .D(_00137_),
    .RESET_B(rst_n),
    .Q(\deser_A.word_buffer[127] ));
 sky130_fd_sc_hd__dfrtp_2 _26330_ (.CLK(A_in_serial_clk),
    .D(_00004_),
    .RESET_B(rst_n),
    .Q(\deser_A.receiving ));
 sky130_fd_sc_hd__dfrtp_2 _26331_ (.CLK(A_in_serial_clk),
    .D(_00138_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_toggle ));
 sky130_fd_sc_hd__dfrtp_2 _26332_ (.CLK(clk),
    .D(_00139_),
    .RESET_B(rst_n),
    .Q(\A_in[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26333_ (.CLK(clk),
    .D(_00140_),
    .RESET_B(rst_n),
    .Q(\A_in[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26334_ (.CLK(clk),
    .D(_00141_),
    .RESET_B(rst_n),
    .Q(\A_in[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26335_ (.CLK(clk),
    .D(_00142_),
    .RESET_B(rst_n),
    .Q(\A_in[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26336_ (.CLK(clk),
    .D(_00143_),
    .RESET_B(rst_n),
    .Q(\A_in[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26337_ (.CLK(clk),
    .D(_00144_),
    .RESET_B(rst_n),
    .Q(\A_in[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26338_ (.CLK(clk),
    .D(_00145_),
    .RESET_B(rst_n),
    .Q(\A_in[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26339_ (.CLK(clk),
    .D(_00146_),
    .RESET_B(rst_n),
    .Q(\A_in[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26340_ (.CLK(clk),
    .D(_00147_),
    .RESET_B(rst_n),
    .Q(\A_in[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26341_ (.CLK(clk),
    .D(_00148_),
    .RESET_B(rst_n),
    .Q(\A_in[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26342_ (.CLK(clk),
    .D(_00149_),
    .RESET_B(rst_n),
    .Q(\A_in[10] ));
 sky130_fd_sc_hd__dfrtp_2 _26343_ (.CLK(clk),
    .D(_00150_),
    .RESET_B(rst_n),
    .Q(\A_in[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26344_ (.CLK(clk),
    .D(_00151_),
    .RESET_B(rst_n),
    .Q(\A_in[12] ));
 sky130_fd_sc_hd__dfrtp_2 _26345_ (.CLK(clk),
    .D(_00152_),
    .RESET_B(rst_n),
    .Q(\A_in[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26346_ (.CLK(clk),
    .D(_00153_),
    .RESET_B(rst_n),
    .Q(\A_in[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26347_ (.CLK(clk),
    .D(_00154_),
    .RESET_B(rst_n),
    .Q(\A_in[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26348_ (.CLK(clk),
    .D(_00155_),
    .RESET_B(rst_n),
    .Q(\A_in[16] ));
 sky130_fd_sc_hd__dfrtp_2 _26349_ (.CLK(clk),
    .D(_00156_),
    .RESET_B(rst_n),
    .Q(\A_in[17] ));
 sky130_fd_sc_hd__dfrtp_2 _26350_ (.CLK(clk),
    .D(_00157_),
    .RESET_B(rst_n),
    .Q(\A_in[18] ));
 sky130_fd_sc_hd__dfrtp_2 _26351_ (.CLK(clk),
    .D(_00158_),
    .RESET_B(rst_n),
    .Q(\A_in[19] ));
 sky130_fd_sc_hd__dfrtp_2 _26352_ (.CLK(clk),
    .D(_00159_),
    .RESET_B(rst_n),
    .Q(\A_in[20] ));
 sky130_fd_sc_hd__dfrtp_2 _26353_ (.CLK(clk),
    .D(_00160_),
    .RESET_B(rst_n),
    .Q(\A_in[21] ));
 sky130_fd_sc_hd__dfrtp_2 _26354_ (.CLK(clk),
    .D(_00161_),
    .RESET_B(rst_n),
    .Q(\A_in[22] ));
 sky130_fd_sc_hd__dfrtp_2 _26355_ (.CLK(clk),
    .D(_00162_),
    .RESET_B(rst_n),
    .Q(\A_in[23] ));
 sky130_fd_sc_hd__dfrtp_2 _26356_ (.CLK(clk),
    .D(_00163_),
    .RESET_B(rst_n),
    .Q(\A_in[24] ));
 sky130_fd_sc_hd__dfrtp_2 _26357_ (.CLK(clk),
    .D(_00164_),
    .RESET_B(rst_n),
    .Q(\A_in[25] ));
 sky130_fd_sc_hd__dfrtp_2 _26358_ (.CLK(clk),
    .D(_00165_),
    .RESET_B(rst_n),
    .Q(\A_in[26] ));
 sky130_fd_sc_hd__dfrtp_2 _26359_ (.CLK(clk),
    .D(_00166_),
    .RESET_B(rst_n),
    .Q(\A_in[27] ));
 sky130_fd_sc_hd__dfrtp_2 _26360_ (.CLK(clk),
    .D(_00167_),
    .RESET_B(rst_n),
    .Q(\A_in[28] ));
 sky130_fd_sc_hd__dfrtp_2 _26361_ (.CLK(clk),
    .D(_00168_),
    .RESET_B(rst_n),
    .Q(\A_in[29] ));
 sky130_fd_sc_hd__dfrtp_2 _26362_ (.CLK(clk),
    .D(_00169_),
    .RESET_B(rst_n),
    .Q(\A_in[30] ));
 sky130_fd_sc_hd__dfrtp_2 _26363_ (.CLK(clk),
    .D(_00170_),
    .RESET_B(rst_n),
    .Q(\A_in[31] ));
 sky130_fd_sc_hd__dfrtp_2 _26364_ (.CLK(clk),
    .D(_00171_),
    .RESET_B(rst_n),
    .Q(\A_in[32] ));
 sky130_fd_sc_hd__dfrtp_2 _26365_ (.CLK(clk),
    .D(_00172_),
    .RESET_B(rst_n),
    .Q(\A_in[33] ));
 sky130_fd_sc_hd__dfrtp_2 _26366_ (.CLK(clk),
    .D(_00173_),
    .RESET_B(rst_n),
    .Q(\A_in[34] ));
 sky130_fd_sc_hd__dfrtp_2 _26367_ (.CLK(clk),
    .D(_00174_),
    .RESET_B(rst_n),
    .Q(\A_in[35] ));
 sky130_fd_sc_hd__dfrtp_2 _26368_ (.CLK(clk),
    .D(_00175_),
    .RESET_B(rst_n),
    .Q(\A_in[36] ));
 sky130_fd_sc_hd__dfrtp_2 _26369_ (.CLK(clk),
    .D(_00176_),
    .RESET_B(rst_n),
    .Q(\A_in[37] ));
 sky130_fd_sc_hd__dfrtp_2 _26370_ (.CLK(clk),
    .D(_00177_),
    .RESET_B(rst_n),
    .Q(\A_in[38] ));
 sky130_fd_sc_hd__dfrtp_2 _26371_ (.CLK(clk),
    .D(_00178_),
    .RESET_B(rst_n),
    .Q(\A_in[39] ));
 sky130_fd_sc_hd__dfrtp_2 _26372_ (.CLK(clk),
    .D(_00179_),
    .RESET_B(rst_n),
    .Q(\A_in[40] ));
 sky130_fd_sc_hd__dfrtp_2 _26373_ (.CLK(clk),
    .D(_00180_),
    .RESET_B(rst_n),
    .Q(\A_in[41] ));
 sky130_fd_sc_hd__dfrtp_2 _26374_ (.CLK(clk),
    .D(_00181_),
    .RESET_B(rst_n),
    .Q(\A_in[42] ));
 sky130_fd_sc_hd__dfrtp_2 _26375_ (.CLK(clk),
    .D(_00182_),
    .RESET_B(rst_n),
    .Q(\A_in[43] ));
 sky130_fd_sc_hd__dfrtp_2 _26376_ (.CLK(clk),
    .D(_00183_),
    .RESET_B(rst_n),
    .Q(\A_in[44] ));
 sky130_fd_sc_hd__dfrtp_2 _26377_ (.CLK(clk),
    .D(_00184_),
    .RESET_B(rst_n),
    .Q(\A_in[45] ));
 sky130_fd_sc_hd__dfrtp_2 _26378_ (.CLK(clk),
    .D(_00185_),
    .RESET_B(rst_n),
    .Q(\A_in[46] ));
 sky130_fd_sc_hd__dfrtp_2 _26379_ (.CLK(clk),
    .D(_00186_),
    .RESET_B(rst_n),
    .Q(\A_in[47] ));
 sky130_fd_sc_hd__dfrtp_2 _26380_ (.CLK(clk),
    .D(_00187_),
    .RESET_B(rst_n),
    .Q(\A_in[48] ));
 sky130_fd_sc_hd__dfrtp_2 _26381_ (.CLK(clk),
    .D(_00188_),
    .RESET_B(rst_n),
    .Q(\A_in[49] ));
 sky130_fd_sc_hd__dfrtp_2 _26382_ (.CLK(clk),
    .D(_00189_),
    .RESET_B(rst_n),
    .Q(\A_in[50] ));
 sky130_fd_sc_hd__dfrtp_2 _26383_ (.CLK(clk),
    .D(_00190_),
    .RESET_B(rst_n),
    .Q(\A_in[51] ));
 sky130_fd_sc_hd__dfrtp_2 _26384_ (.CLK(clk),
    .D(_00191_),
    .RESET_B(rst_n),
    .Q(\A_in[52] ));
 sky130_fd_sc_hd__dfrtp_2 _26385_ (.CLK(clk),
    .D(_00192_),
    .RESET_B(rst_n),
    .Q(\A_in[53] ));
 sky130_fd_sc_hd__dfrtp_2 _26386_ (.CLK(clk),
    .D(_00193_),
    .RESET_B(rst_n),
    .Q(\A_in[54] ));
 sky130_fd_sc_hd__dfrtp_2 _26387_ (.CLK(clk),
    .D(_00194_),
    .RESET_B(rst_n),
    .Q(\A_in[55] ));
 sky130_fd_sc_hd__dfrtp_2 _26388_ (.CLK(clk),
    .D(_00195_),
    .RESET_B(rst_n),
    .Q(\A_in[56] ));
 sky130_fd_sc_hd__dfrtp_2 _26389_ (.CLK(clk),
    .D(_00196_),
    .RESET_B(rst_n),
    .Q(\A_in[57] ));
 sky130_fd_sc_hd__dfrtp_2 _26390_ (.CLK(clk),
    .D(_00197_),
    .RESET_B(rst_n),
    .Q(\A_in[58] ));
 sky130_fd_sc_hd__dfrtp_2 _26391_ (.CLK(clk),
    .D(_00198_),
    .RESET_B(rst_n),
    .Q(\A_in[59] ));
 sky130_fd_sc_hd__dfrtp_2 _26392_ (.CLK(clk),
    .D(_00199_),
    .RESET_B(rst_n),
    .Q(\A_in[60] ));
 sky130_fd_sc_hd__dfrtp_2 _26393_ (.CLK(clk),
    .D(_00200_),
    .RESET_B(rst_n),
    .Q(\A_in[61] ));
 sky130_fd_sc_hd__dfrtp_2 _26394_ (.CLK(clk),
    .D(_00201_),
    .RESET_B(rst_n),
    .Q(\A_in[62] ));
 sky130_fd_sc_hd__dfrtp_2 _26395_ (.CLK(clk),
    .D(_00202_),
    .RESET_B(rst_n),
    .Q(\A_in[63] ));
 sky130_fd_sc_hd__dfrtp_2 _26396_ (.CLK(clk),
    .D(_00203_),
    .RESET_B(rst_n),
    .Q(\A_in[64] ));
 sky130_fd_sc_hd__dfrtp_2 _26397_ (.CLK(clk),
    .D(_00204_),
    .RESET_B(rst_n),
    .Q(\A_in[65] ));
 sky130_fd_sc_hd__dfrtp_2 _26398_ (.CLK(clk),
    .D(_00205_),
    .RESET_B(rst_n),
    .Q(\A_in[66] ));
 sky130_fd_sc_hd__dfrtp_2 _26399_ (.CLK(clk),
    .D(_00206_),
    .RESET_B(rst_n),
    .Q(\A_in[67] ));
 sky130_fd_sc_hd__dfrtp_2 _26400_ (.CLK(clk),
    .D(_00207_),
    .RESET_B(rst_n),
    .Q(\A_in[68] ));
 sky130_fd_sc_hd__dfrtp_2 _26401_ (.CLK(clk),
    .D(_00208_),
    .RESET_B(rst_n),
    .Q(\A_in[69] ));
 sky130_fd_sc_hd__dfrtp_2 _26402_ (.CLK(clk),
    .D(_00209_),
    .RESET_B(rst_n),
    .Q(\A_in[70] ));
 sky130_fd_sc_hd__dfrtp_2 _26403_ (.CLK(clk),
    .D(_00210_),
    .RESET_B(rst_n),
    .Q(\A_in[71] ));
 sky130_fd_sc_hd__dfrtp_2 _26404_ (.CLK(clk),
    .D(_00211_),
    .RESET_B(rst_n),
    .Q(\A_in[72] ));
 sky130_fd_sc_hd__dfrtp_2 _26405_ (.CLK(clk),
    .D(_00212_),
    .RESET_B(rst_n),
    .Q(\A_in[73] ));
 sky130_fd_sc_hd__dfrtp_2 _26406_ (.CLK(clk),
    .D(_00213_),
    .RESET_B(rst_n),
    .Q(\A_in[74] ));
 sky130_fd_sc_hd__dfrtp_2 _26407_ (.CLK(clk),
    .D(_00214_),
    .RESET_B(rst_n),
    .Q(\A_in[75] ));
 sky130_fd_sc_hd__dfrtp_2 _26408_ (.CLK(clk),
    .D(_00215_),
    .RESET_B(rst_n),
    .Q(\A_in[76] ));
 sky130_fd_sc_hd__dfrtp_2 _26409_ (.CLK(clk),
    .D(_00216_),
    .RESET_B(rst_n),
    .Q(\A_in[77] ));
 sky130_fd_sc_hd__dfrtp_2 _26410_ (.CLK(clk),
    .D(_00217_),
    .RESET_B(rst_n),
    .Q(\A_in[78] ));
 sky130_fd_sc_hd__dfrtp_2 _26411_ (.CLK(clk),
    .D(_00218_),
    .RESET_B(rst_n),
    .Q(\A_in[79] ));
 sky130_fd_sc_hd__dfrtp_2 _26412_ (.CLK(clk),
    .D(_00219_),
    .RESET_B(rst_n),
    .Q(\A_in[80] ));
 sky130_fd_sc_hd__dfrtp_2 _26413_ (.CLK(clk),
    .D(_00220_),
    .RESET_B(rst_n),
    .Q(\A_in[81] ));
 sky130_fd_sc_hd__dfrtp_2 _26414_ (.CLK(clk),
    .D(_00221_),
    .RESET_B(rst_n),
    .Q(\A_in[82] ));
 sky130_fd_sc_hd__dfrtp_2 _26415_ (.CLK(clk),
    .D(_00222_),
    .RESET_B(rst_n),
    .Q(\A_in[83] ));
 sky130_fd_sc_hd__dfrtp_2 _26416_ (.CLK(clk),
    .D(_00223_),
    .RESET_B(rst_n),
    .Q(\A_in[84] ));
 sky130_fd_sc_hd__dfrtp_2 _26417_ (.CLK(clk),
    .D(_00224_),
    .RESET_B(rst_n),
    .Q(\A_in[85] ));
 sky130_fd_sc_hd__dfrtp_2 _26418_ (.CLK(clk),
    .D(_00225_),
    .RESET_B(rst_n),
    .Q(\A_in[86] ));
 sky130_fd_sc_hd__dfrtp_2 _26419_ (.CLK(clk),
    .D(_00226_),
    .RESET_B(rst_n),
    .Q(\A_in[87] ));
 sky130_fd_sc_hd__dfrtp_2 _26420_ (.CLK(clk),
    .D(_00227_),
    .RESET_B(rst_n),
    .Q(\A_in[88] ));
 sky130_fd_sc_hd__dfrtp_2 _26421_ (.CLK(clk),
    .D(_00228_),
    .RESET_B(rst_n),
    .Q(\A_in[89] ));
 sky130_fd_sc_hd__dfrtp_2 _26422_ (.CLK(clk),
    .D(_00229_),
    .RESET_B(rst_n),
    .Q(\A_in[90] ));
 sky130_fd_sc_hd__dfrtp_2 _26423_ (.CLK(clk),
    .D(_00230_),
    .RESET_B(rst_n),
    .Q(\A_in[91] ));
 sky130_fd_sc_hd__dfrtp_2 _26424_ (.CLK(clk),
    .D(_00231_),
    .RESET_B(rst_n),
    .Q(\A_in[92] ));
 sky130_fd_sc_hd__dfrtp_2 _26425_ (.CLK(clk),
    .D(_00232_),
    .RESET_B(rst_n),
    .Q(\A_in[93] ));
 sky130_fd_sc_hd__dfrtp_2 _26426_ (.CLK(clk),
    .D(_00233_),
    .RESET_B(rst_n),
    .Q(\A_in[94] ));
 sky130_fd_sc_hd__dfrtp_2 _26427_ (.CLK(clk),
    .D(_00234_),
    .RESET_B(rst_n),
    .Q(\A_in[95] ));
 sky130_fd_sc_hd__dfrtp_2 _26428_ (.CLK(clk),
    .D(_00235_),
    .RESET_B(rst_n),
    .Q(\A_in[96] ));
 sky130_fd_sc_hd__dfrtp_2 _26429_ (.CLK(clk),
    .D(_00236_),
    .RESET_B(rst_n),
    .Q(\A_in[97] ));
 sky130_fd_sc_hd__dfrtp_2 _26430_ (.CLK(clk),
    .D(_00237_),
    .RESET_B(rst_n),
    .Q(\A_in[98] ));
 sky130_fd_sc_hd__dfrtp_2 _26431_ (.CLK(clk),
    .D(_00238_),
    .RESET_B(rst_n),
    .Q(\A_in[99] ));
 sky130_fd_sc_hd__dfrtp_2 _26432_ (.CLK(clk),
    .D(_00239_),
    .RESET_B(rst_n),
    .Q(\A_in[100] ));
 sky130_fd_sc_hd__dfrtp_2 _26433_ (.CLK(clk),
    .D(_00240_),
    .RESET_B(rst_n),
    .Q(\A_in[101] ));
 sky130_fd_sc_hd__dfrtp_2 _26434_ (.CLK(clk),
    .D(_00241_),
    .RESET_B(rst_n),
    .Q(\A_in[102] ));
 sky130_fd_sc_hd__dfrtp_2 _26435_ (.CLK(clk),
    .D(_00242_),
    .RESET_B(rst_n),
    .Q(\A_in[103] ));
 sky130_fd_sc_hd__dfrtp_2 _26436_ (.CLK(clk),
    .D(_00243_),
    .RESET_B(rst_n),
    .Q(\A_in[104] ));
 sky130_fd_sc_hd__dfrtp_2 _26437_ (.CLK(clk),
    .D(_00244_),
    .RESET_B(rst_n),
    .Q(\A_in[105] ));
 sky130_fd_sc_hd__dfrtp_2 _26438_ (.CLK(clk),
    .D(_00245_),
    .RESET_B(rst_n),
    .Q(\A_in[106] ));
 sky130_fd_sc_hd__dfrtp_2 _26439_ (.CLK(clk),
    .D(_00246_),
    .RESET_B(rst_n),
    .Q(\A_in[107] ));
 sky130_fd_sc_hd__dfrtp_2 _26440_ (.CLK(clk),
    .D(_00247_),
    .RESET_B(rst_n),
    .Q(\A_in[108] ));
 sky130_fd_sc_hd__dfrtp_2 _26441_ (.CLK(clk),
    .D(_00248_),
    .RESET_B(rst_n),
    .Q(\A_in[109] ));
 sky130_fd_sc_hd__dfrtp_2 _26442_ (.CLK(clk),
    .D(_00249_),
    .RESET_B(rst_n),
    .Q(\A_in[110] ));
 sky130_fd_sc_hd__dfrtp_2 _26443_ (.CLK(clk),
    .D(_00250_),
    .RESET_B(rst_n),
    .Q(\A_in[111] ));
 sky130_fd_sc_hd__dfrtp_2 _26444_ (.CLK(clk),
    .D(_00251_),
    .RESET_B(rst_n),
    .Q(\A_in[112] ));
 sky130_fd_sc_hd__dfrtp_2 _26445_ (.CLK(clk),
    .D(_00252_),
    .RESET_B(rst_n),
    .Q(\A_in[113] ));
 sky130_fd_sc_hd__dfrtp_2 _26446_ (.CLK(clk),
    .D(_00253_),
    .RESET_B(rst_n),
    .Q(\A_in[114] ));
 sky130_fd_sc_hd__dfrtp_2 _26447_ (.CLK(clk),
    .D(_00254_),
    .RESET_B(rst_n),
    .Q(\A_in[115] ));
 sky130_fd_sc_hd__dfrtp_2 _26448_ (.CLK(clk),
    .D(_00255_),
    .RESET_B(rst_n),
    .Q(\A_in[116] ));
 sky130_fd_sc_hd__dfrtp_2 _26449_ (.CLK(clk),
    .D(_00256_),
    .RESET_B(rst_n),
    .Q(\A_in[117] ));
 sky130_fd_sc_hd__dfrtp_2 _26450_ (.CLK(clk),
    .D(_00257_),
    .RESET_B(rst_n),
    .Q(\A_in[118] ));
 sky130_fd_sc_hd__dfrtp_2 _26451_ (.CLK(clk),
    .D(_00258_),
    .RESET_B(rst_n),
    .Q(\A_in[119] ));
 sky130_fd_sc_hd__dfrtp_2 _26452_ (.CLK(clk),
    .D(_00259_),
    .RESET_B(rst_n),
    .Q(\A_in[120] ));
 sky130_fd_sc_hd__dfrtp_2 _26453_ (.CLK(clk),
    .D(_00260_),
    .RESET_B(rst_n),
    .Q(\A_in[121] ));
 sky130_fd_sc_hd__dfrtp_2 _26454_ (.CLK(clk),
    .D(_00261_),
    .RESET_B(rst_n),
    .Q(\A_in[122] ));
 sky130_fd_sc_hd__dfrtp_2 _26455_ (.CLK(clk),
    .D(_00262_),
    .RESET_B(rst_n),
    .Q(\A_in[123] ));
 sky130_fd_sc_hd__dfrtp_2 _26456_ (.CLK(clk),
    .D(_00263_),
    .RESET_B(rst_n),
    .Q(\A_in[124] ));
 sky130_fd_sc_hd__dfrtp_2 _26457_ (.CLK(clk),
    .D(_00264_),
    .RESET_B(rst_n),
    .Q(\A_in[125] ));
 sky130_fd_sc_hd__dfrtp_2 _26458_ (.CLK(clk),
    .D(_00265_),
    .RESET_B(rst_n),
    .Q(\A_in[126] ));
 sky130_fd_sc_hd__dfrtp_2 _26459_ (.CLK(clk),
    .D(_00266_),
    .RESET_B(rst_n),
    .Q(\A_in[127] ));
 sky130_fd_sc_hd__dfrtp_2 _26460_ (.CLK(A_in_serial_clk),
    .D(_00267_),
    .RESET_B(rst_n),
    .Q(\deser_A.bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26461_ (.CLK(A_in_serial_clk),
    .D(_00268_),
    .RESET_B(rst_n),
    .Q(\deser_A.bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26462_ (.CLK(A_in_serial_clk),
    .D(_00269_),
    .RESET_B(rst_n),
    .Q(\deser_A.bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26463_ (.CLK(A_in_serial_clk),
    .D(_00270_),
    .RESET_B(rst_n),
    .Q(\deser_A.bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26464_ (.CLK(A_in_serial_clk),
    .D(_00271_),
    .RESET_B(rst_n),
    .Q(\deser_A.bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26465_ (.CLK(A_in_serial_clk),
    .D(_00272_),
    .RESET_B(rst_n),
    .Q(\deser_A.bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26466_ (.CLK(A_in_serial_clk),
    .D(_00273_),
    .RESET_B(rst_n),
    .Q(\deser_A.bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26467_ (.CLK(clk),
    .D(\deser_A.serial_toggle_sync1 ),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_toggle_sync2 ));
 sky130_fd_sc_hd__dfrtp_2 _26468_ (.CLK(A_in_serial_clk),
    .D(_00002_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word_ready ));
 sky130_fd_sc_hd__dfrtp_2 _26469_ (.CLK(clk),
    .D(\deser_A.serial_toggle ),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_toggle_sync1 ));
 sky130_fd_sc_hd__dfrtp_2 _26470_ (.CLK(clk),
    .D(_00003_),
    .RESET_B(rst_n),
    .Q(A_in_valid));
 sky130_fd_sc_hd__dfrtp_2 _26471_ (.CLK(A_in_serial_clk),
    .D(_00274_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26472_ (.CLK(A_in_serial_clk),
    .D(_00275_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26473_ (.CLK(A_in_serial_clk),
    .D(_00276_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26474_ (.CLK(A_in_serial_clk),
    .D(_00277_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26475_ (.CLK(A_in_serial_clk),
    .D(_00278_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26476_ (.CLK(A_in_serial_clk),
    .D(_00279_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26477_ (.CLK(A_in_serial_clk),
    .D(_00280_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26478_ (.CLK(A_in_serial_clk),
    .D(_00281_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26479_ (.CLK(A_in_serial_clk),
    .D(_00282_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26480_ (.CLK(A_in_serial_clk),
    .D(_00283_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _26481_ (.CLK(A_in_serial_clk),
    .D(_00284_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26482_ (.CLK(A_in_serial_clk),
    .D(_00285_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _26483_ (.CLK(A_in_serial_clk),
    .D(_00286_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26484_ (.CLK(A_in_serial_clk),
    .D(_00287_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26485_ (.CLK(A_in_serial_clk),
    .D(_00288_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26486_ (.CLK(A_in_serial_clk),
    .D(_00289_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[16] ));
 sky130_fd_sc_hd__dfrtp_2 _26487_ (.CLK(A_in_serial_clk),
    .D(_00290_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[17] ));
 sky130_fd_sc_hd__dfrtp_2 _26488_ (.CLK(A_in_serial_clk),
    .D(_00291_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[18] ));
 sky130_fd_sc_hd__dfrtp_2 _26489_ (.CLK(A_in_serial_clk),
    .D(_00292_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[19] ));
 sky130_fd_sc_hd__dfrtp_2 _26490_ (.CLK(A_in_serial_clk),
    .D(_00293_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[20] ));
 sky130_fd_sc_hd__dfrtp_2 _26491_ (.CLK(A_in_serial_clk),
    .D(_00294_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[21] ));
 sky130_fd_sc_hd__dfrtp_2 _26492_ (.CLK(A_in_serial_clk),
    .D(_00295_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[22] ));
 sky130_fd_sc_hd__dfrtp_2 _26493_ (.CLK(A_in_serial_clk),
    .D(_00296_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[23] ));
 sky130_fd_sc_hd__dfrtp_2 _26494_ (.CLK(A_in_serial_clk),
    .D(_00297_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[24] ));
 sky130_fd_sc_hd__dfrtp_2 _26495_ (.CLK(A_in_serial_clk),
    .D(_00298_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[25] ));
 sky130_fd_sc_hd__dfrtp_2 _26496_ (.CLK(A_in_serial_clk),
    .D(_00299_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[26] ));
 sky130_fd_sc_hd__dfrtp_2 _26497_ (.CLK(A_in_serial_clk),
    .D(_00300_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[27] ));
 sky130_fd_sc_hd__dfrtp_2 _26498_ (.CLK(A_in_serial_clk),
    .D(_00301_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[28] ));
 sky130_fd_sc_hd__dfrtp_2 _26499_ (.CLK(A_in_serial_clk),
    .D(_00302_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[29] ));
 sky130_fd_sc_hd__dfrtp_2 _26500_ (.CLK(A_in_serial_clk),
    .D(_00303_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[30] ));
 sky130_fd_sc_hd__dfrtp_2 _26501_ (.CLK(A_in_serial_clk),
    .D(_00304_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[31] ));
 sky130_fd_sc_hd__dfrtp_2 _26502_ (.CLK(A_in_serial_clk),
    .D(_00305_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[32] ));
 sky130_fd_sc_hd__dfrtp_2 _26503_ (.CLK(A_in_serial_clk),
    .D(_00306_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[33] ));
 sky130_fd_sc_hd__dfrtp_2 _26504_ (.CLK(A_in_serial_clk),
    .D(_00307_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[34] ));
 sky130_fd_sc_hd__dfrtp_2 _26505_ (.CLK(A_in_serial_clk),
    .D(_00308_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[35] ));
 sky130_fd_sc_hd__dfrtp_2 _26506_ (.CLK(A_in_serial_clk),
    .D(_00309_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[36] ));
 sky130_fd_sc_hd__dfrtp_2 _26507_ (.CLK(A_in_serial_clk),
    .D(_00310_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[37] ));
 sky130_fd_sc_hd__dfrtp_2 _26508_ (.CLK(A_in_serial_clk),
    .D(_00311_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[38] ));
 sky130_fd_sc_hd__dfrtp_2 _26509_ (.CLK(A_in_serial_clk),
    .D(_00312_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[39] ));
 sky130_fd_sc_hd__dfrtp_2 _26510_ (.CLK(A_in_serial_clk),
    .D(_00313_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[40] ));
 sky130_fd_sc_hd__dfrtp_2 _26511_ (.CLK(A_in_serial_clk),
    .D(_00314_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[41] ));
 sky130_fd_sc_hd__dfrtp_2 _26512_ (.CLK(A_in_serial_clk),
    .D(_00315_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[42] ));
 sky130_fd_sc_hd__dfrtp_2 _26513_ (.CLK(A_in_serial_clk),
    .D(_00316_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[43] ));
 sky130_fd_sc_hd__dfrtp_2 _26514_ (.CLK(A_in_serial_clk),
    .D(_00317_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[44] ));
 sky130_fd_sc_hd__dfrtp_2 _26515_ (.CLK(A_in_serial_clk),
    .D(_00318_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[45] ));
 sky130_fd_sc_hd__dfrtp_2 _26516_ (.CLK(A_in_serial_clk),
    .D(_00319_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[46] ));
 sky130_fd_sc_hd__dfrtp_2 _26517_ (.CLK(A_in_serial_clk),
    .D(_00320_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[47] ));
 sky130_fd_sc_hd__dfrtp_2 _26518_ (.CLK(A_in_serial_clk),
    .D(_00321_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[48] ));
 sky130_fd_sc_hd__dfrtp_2 _26519_ (.CLK(A_in_serial_clk),
    .D(_00322_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[49] ));
 sky130_fd_sc_hd__dfrtp_2 _26520_ (.CLK(A_in_serial_clk),
    .D(_00323_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[50] ));
 sky130_fd_sc_hd__dfrtp_2 _26521_ (.CLK(A_in_serial_clk),
    .D(_00324_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[51] ));
 sky130_fd_sc_hd__dfrtp_2 _26522_ (.CLK(A_in_serial_clk),
    .D(_00325_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[52] ));
 sky130_fd_sc_hd__dfrtp_2 _26523_ (.CLK(A_in_serial_clk),
    .D(_00326_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[53] ));
 sky130_fd_sc_hd__dfrtp_2 _26524_ (.CLK(A_in_serial_clk),
    .D(_00327_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[54] ));
 sky130_fd_sc_hd__dfrtp_2 _26525_ (.CLK(A_in_serial_clk),
    .D(_00328_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[55] ));
 sky130_fd_sc_hd__dfrtp_2 _26526_ (.CLK(A_in_serial_clk),
    .D(_00329_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[56] ));
 sky130_fd_sc_hd__dfrtp_2 _26527_ (.CLK(A_in_serial_clk),
    .D(_00330_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[57] ));
 sky130_fd_sc_hd__dfrtp_2 _26528_ (.CLK(A_in_serial_clk),
    .D(_00331_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[58] ));
 sky130_fd_sc_hd__dfrtp_2 _26529_ (.CLK(A_in_serial_clk),
    .D(_00332_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[59] ));
 sky130_fd_sc_hd__dfrtp_2 _26530_ (.CLK(A_in_serial_clk),
    .D(_00333_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[60] ));
 sky130_fd_sc_hd__dfrtp_2 _26531_ (.CLK(A_in_serial_clk),
    .D(_00334_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[61] ));
 sky130_fd_sc_hd__dfrtp_2 _26532_ (.CLK(A_in_serial_clk),
    .D(_00335_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[62] ));
 sky130_fd_sc_hd__dfrtp_2 _26533_ (.CLK(A_in_serial_clk),
    .D(_00336_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[63] ));
 sky130_fd_sc_hd__dfrtp_2 _26534_ (.CLK(A_in_serial_clk),
    .D(_00337_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[64] ));
 sky130_fd_sc_hd__dfrtp_2 _26535_ (.CLK(A_in_serial_clk),
    .D(_00338_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[65] ));
 sky130_fd_sc_hd__dfrtp_2 _26536_ (.CLK(A_in_serial_clk),
    .D(_00339_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[66] ));
 sky130_fd_sc_hd__dfrtp_2 _26537_ (.CLK(A_in_serial_clk),
    .D(_00340_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[67] ));
 sky130_fd_sc_hd__dfrtp_2 _26538_ (.CLK(A_in_serial_clk),
    .D(_00341_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[68] ));
 sky130_fd_sc_hd__dfrtp_2 _26539_ (.CLK(A_in_serial_clk),
    .D(_00342_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[69] ));
 sky130_fd_sc_hd__dfrtp_2 _26540_ (.CLK(A_in_serial_clk),
    .D(_00343_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[70] ));
 sky130_fd_sc_hd__dfrtp_2 _26541_ (.CLK(A_in_serial_clk),
    .D(_00344_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[71] ));
 sky130_fd_sc_hd__dfrtp_2 _26542_ (.CLK(A_in_serial_clk),
    .D(_00345_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[72] ));
 sky130_fd_sc_hd__dfrtp_2 _26543_ (.CLK(A_in_serial_clk),
    .D(_00346_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[73] ));
 sky130_fd_sc_hd__dfrtp_2 _26544_ (.CLK(A_in_serial_clk),
    .D(_00347_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[74] ));
 sky130_fd_sc_hd__dfrtp_2 _26545_ (.CLK(A_in_serial_clk),
    .D(_00348_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[75] ));
 sky130_fd_sc_hd__dfrtp_2 _26546_ (.CLK(A_in_serial_clk),
    .D(_00349_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[76] ));
 sky130_fd_sc_hd__dfrtp_2 _26547_ (.CLK(A_in_serial_clk),
    .D(_00350_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[77] ));
 sky130_fd_sc_hd__dfrtp_2 _26548_ (.CLK(A_in_serial_clk),
    .D(_00351_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[78] ));
 sky130_fd_sc_hd__dfrtp_2 _26549_ (.CLK(A_in_serial_clk),
    .D(_00352_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[79] ));
 sky130_fd_sc_hd__dfrtp_2 _26550_ (.CLK(A_in_serial_clk),
    .D(_00353_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[80] ));
 sky130_fd_sc_hd__dfrtp_2 _26551_ (.CLK(A_in_serial_clk),
    .D(_00354_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[81] ));
 sky130_fd_sc_hd__dfrtp_2 _26552_ (.CLK(A_in_serial_clk),
    .D(_00355_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[82] ));
 sky130_fd_sc_hd__dfrtp_2 _26553_ (.CLK(A_in_serial_clk),
    .D(_00356_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[83] ));
 sky130_fd_sc_hd__dfrtp_2 _26554_ (.CLK(A_in_serial_clk),
    .D(_00357_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[84] ));
 sky130_fd_sc_hd__dfrtp_2 _26555_ (.CLK(A_in_serial_clk),
    .D(_00358_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[85] ));
 sky130_fd_sc_hd__dfrtp_2 _26556_ (.CLK(A_in_serial_clk),
    .D(_00359_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[86] ));
 sky130_fd_sc_hd__dfrtp_2 _26557_ (.CLK(A_in_serial_clk),
    .D(_00360_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[87] ));
 sky130_fd_sc_hd__dfrtp_2 _26558_ (.CLK(A_in_serial_clk),
    .D(_00361_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[88] ));
 sky130_fd_sc_hd__dfrtp_2 _26559_ (.CLK(A_in_serial_clk),
    .D(_00362_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[89] ));
 sky130_fd_sc_hd__dfrtp_2 _26560_ (.CLK(A_in_serial_clk),
    .D(_00363_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[90] ));
 sky130_fd_sc_hd__dfrtp_2 _26561_ (.CLK(A_in_serial_clk),
    .D(_00364_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[91] ));
 sky130_fd_sc_hd__dfrtp_2 _26562_ (.CLK(A_in_serial_clk),
    .D(_00365_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[92] ));
 sky130_fd_sc_hd__dfrtp_2 _26563_ (.CLK(A_in_serial_clk),
    .D(_00366_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[93] ));
 sky130_fd_sc_hd__dfrtp_2 _26564_ (.CLK(A_in_serial_clk),
    .D(_00367_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[94] ));
 sky130_fd_sc_hd__dfrtp_2 _26565_ (.CLK(A_in_serial_clk),
    .D(_00368_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[95] ));
 sky130_fd_sc_hd__dfrtp_2 _26566_ (.CLK(A_in_serial_clk),
    .D(_00369_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[96] ));
 sky130_fd_sc_hd__dfrtp_2 _26567_ (.CLK(A_in_serial_clk),
    .D(_00370_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[97] ));
 sky130_fd_sc_hd__dfrtp_2 _26568_ (.CLK(A_in_serial_clk),
    .D(_00371_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[98] ));
 sky130_fd_sc_hd__dfrtp_2 _26569_ (.CLK(A_in_serial_clk),
    .D(_00372_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[99] ));
 sky130_fd_sc_hd__dfrtp_2 _26570_ (.CLK(A_in_serial_clk),
    .D(_00373_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[100] ));
 sky130_fd_sc_hd__dfrtp_2 _26571_ (.CLK(A_in_serial_clk),
    .D(_00374_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[101] ));
 sky130_fd_sc_hd__dfrtp_2 _26572_ (.CLK(A_in_serial_clk),
    .D(_00375_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[102] ));
 sky130_fd_sc_hd__dfrtp_2 _26573_ (.CLK(A_in_serial_clk),
    .D(_00376_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[103] ));
 sky130_fd_sc_hd__dfrtp_2 _26574_ (.CLK(A_in_serial_clk),
    .D(_00377_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[104] ));
 sky130_fd_sc_hd__dfrtp_2 _26575_ (.CLK(A_in_serial_clk),
    .D(_00378_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[105] ));
 sky130_fd_sc_hd__dfrtp_2 _26576_ (.CLK(A_in_serial_clk),
    .D(_00379_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[106] ));
 sky130_fd_sc_hd__dfrtp_2 _26577_ (.CLK(A_in_serial_clk),
    .D(_00380_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[107] ));
 sky130_fd_sc_hd__dfrtp_2 _26578_ (.CLK(A_in_serial_clk),
    .D(_00381_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[108] ));
 sky130_fd_sc_hd__dfrtp_2 _26579_ (.CLK(A_in_serial_clk),
    .D(_00382_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[109] ));
 sky130_fd_sc_hd__dfrtp_2 _26580_ (.CLK(A_in_serial_clk),
    .D(_00383_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[110] ));
 sky130_fd_sc_hd__dfrtp_2 _26581_ (.CLK(A_in_serial_clk),
    .D(_00384_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[111] ));
 sky130_fd_sc_hd__dfrtp_2 _26582_ (.CLK(A_in_serial_clk),
    .D(_00385_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[112] ));
 sky130_fd_sc_hd__dfrtp_2 _26583_ (.CLK(A_in_serial_clk),
    .D(_00386_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[113] ));
 sky130_fd_sc_hd__dfrtp_2 _26584_ (.CLK(A_in_serial_clk),
    .D(_00387_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[114] ));
 sky130_fd_sc_hd__dfrtp_2 _26585_ (.CLK(A_in_serial_clk),
    .D(_00388_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[115] ));
 sky130_fd_sc_hd__dfrtp_2 _26586_ (.CLK(A_in_serial_clk),
    .D(_00389_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[116] ));
 sky130_fd_sc_hd__dfrtp_2 _26587_ (.CLK(A_in_serial_clk),
    .D(_00390_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[117] ));
 sky130_fd_sc_hd__dfrtp_2 _26588_ (.CLK(A_in_serial_clk),
    .D(_00391_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[118] ));
 sky130_fd_sc_hd__dfrtp_2 _26589_ (.CLK(A_in_serial_clk),
    .D(_00392_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[119] ));
 sky130_fd_sc_hd__dfrtp_2 _26590_ (.CLK(A_in_serial_clk),
    .D(_00393_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[120] ));
 sky130_fd_sc_hd__dfrtp_2 _26591_ (.CLK(A_in_serial_clk),
    .D(_00394_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[121] ));
 sky130_fd_sc_hd__dfrtp_2 _26592_ (.CLK(A_in_serial_clk),
    .D(_00395_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[122] ));
 sky130_fd_sc_hd__dfrtp_2 _26593_ (.CLK(A_in_serial_clk),
    .D(_00396_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[123] ));
 sky130_fd_sc_hd__dfrtp_2 _26594_ (.CLK(A_in_serial_clk),
    .D(_00397_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[124] ));
 sky130_fd_sc_hd__dfrtp_2 _26595_ (.CLK(A_in_serial_clk),
    .D(_00398_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[125] ));
 sky130_fd_sc_hd__dfrtp_2 _26596_ (.CLK(A_in_serial_clk),
    .D(_00399_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[126] ));
 sky130_fd_sc_hd__dfrtp_2 _26597_ (.CLK(A_in_serial_clk),
    .D(_00400_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[127] ));
 sky130_fd_sc_hd__dfrtp_2 _26598_ (.CLK(B_in_serial_clk),
    .D(_00401_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26599_ (.CLK(B_in_serial_clk),
    .D(_00402_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26600_ (.CLK(B_in_serial_clk),
    .D(_00403_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26601_ (.CLK(B_in_serial_clk),
    .D(_00404_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26602_ (.CLK(B_in_serial_clk),
    .D(_00405_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26603_ (.CLK(B_in_serial_clk),
    .D(_00406_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26604_ (.CLK(B_in_serial_clk),
    .D(_00407_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26605_ (.CLK(B_in_serial_clk),
    .D(_00408_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26606_ (.CLK(B_in_serial_clk),
    .D(_00409_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26607_ (.CLK(B_in_serial_clk),
    .D(_00410_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26608_ (.CLK(B_in_serial_clk),
    .D(_00411_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[10] ));
 sky130_fd_sc_hd__dfrtp_2 _26609_ (.CLK(B_in_serial_clk),
    .D(_00412_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26610_ (.CLK(B_in_serial_clk),
    .D(_00413_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[12] ));
 sky130_fd_sc_hd__dfrtp_2 _26611_ (.CLK(B_in_serial_clk),
    .D(_00414_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26612_ (.CLK(B_in_serial_clk),
    .D(_00415_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26613_ (.CLK(B_in_serial_clk),
    .D(_00416_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26614_ (.CLK(B_in_serial_clk),
    .D(_00417_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[16] ));
 sky130_fd_sc_hd__dfrtp_2 _26615_ (.CLK(B_in_serial_clk),
    .D(_00418_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[17] ));
 sky130_fd_sc_hd__dfrtp_2 _26616_ (.CLK(B_in_serial_clk),
    .D(_00419_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[18] ));
 sky130_fd_sc_hd__dfrtp_2 _26617_ (.CLK(B_in_serial_clk),
    .D(_00420_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[19] ));
 sky130_fd_sc_hd__dfrtp_2 _26618_ (.CLK(B_in_serial_clk),
    .D(_00421_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[20] ));
 sky130_fd_sc_hd__dfrtp_2 _26619_ (.CLK(B_in_serial_clk),
    .D(_00422_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[21] ));
 sky130_fd_sc_hd__dfrtp_2 _26620_ (.CLK(B_in_serial_clk),
    .D(_00423_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[22] ));
 sky130_fd_sc_hd__dfrtp_2 _26621_ (.CLK(B_in_serial_clk),
    .D(_00424_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[23] ));
 sky130_fd_sc_hd__dfrtp_2 _26622_ (.CLK(B_in_serial_clk),
    .D(_00425_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[24] ));
 sky130_fd_sc_hd__dfrtp_2 _26623_ (.CLK(B_in_serial_clk),
    .D(_00426_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[25] ));
 sky130_fd_sc_hd__dfrtp_2 _26624_ (.CLK(B_in_serial_clk),
    .D(_00427_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[26] ));
 sky130_fd_sc_hd__dfrtp_2 _26625_ (.CLK(B_in_serial_clk),
    .D(_00428_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[27] ));
 sky130_fd_sc_hd__dfrtp_2 _26626_ (.CLK(B_in_serial_clk),
    .D(_00429_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[28] ));
 sky130_fd_sc_hd__dfrtp_2 _26627_ (.CLK(B_in_serial_clk),
    .D(_00430_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[29] ));
 sky130_fd_sc_hd__dfrtp_2 _26628_ (.CLK(B_in_serial_clk),
    .D(_00431_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[30] ));
 sky130_fd_sc_hd__dfrtp_2 _26629_ (.CLK(B_in_serial_clk),
    .D(_00432_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[31] ));
 sky130_fd_sc_hd__dfrtp_2 _26630_ (.CLK(B_in_serial_clk),
    .D(_00433_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[32] ));
 sky130_fd_sc_hd__dfrtp_2 _26631_ (.CLK(B_in_serial_clk),
    .D(_00434_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[33] ));
 sky130_fd_sc_hd__dfrtp_2 _26632_ (.CLK(B_in_serial_clk),
    .D(_00435_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[34] ));
 sky130_fd_sc_hd__dfrtp_2 _26633_ (.CLK(B_in_serial_clk),
    .D(_00436_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[35] ));
 sky130_fd_sc_hd__dfrtp_2 _26634_ (.CLK(B_in_serial_clk),
    .D(_00437_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[36] ));
 sky130_fd_sc_hd__dfrtp_2 _26635_ (.CLK(B_in_serial_clk),
    .D(_00438_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[37] ));
 sky130_fd_sc_hd__dfrtp_2 _26636_ (.CLK(B_in_serial_clk),
    .D(_00439_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[38] ));
 sky130_fd_sc_hd__dfrtp_2 _26637_ (.CLK(B_in_serial_clk),
    .D(_00440_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[39] ));
 sky130_fd_sc_hd__dfrtp_2 _26638_ (.CLK(B_in_serial_clk),
    .D(_00441_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[40] ));
 sky130_fd_sc_hd__dfrtp_2 _26639_ (.CLK(B_in_serial_clk),
    .D(_00442_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[41] ));
 sky130_fd_sc_hd__dfrtp_2 _26640_ (.CLK(B_in_serial_clk),
    .D(_00443_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[42] ));
 sky130_fd_sc_hd__dfrtp_2 _26641_ (.CLK(B_in_serial_clk),
    .D(_00444_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[43] ));
 sky130_fd_sc_hd__dfrtp_2 _26642_ (.CLK(B_in_serial_clk),
    .D(_00445_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[44] ));
 sky130_fd_sc_hd__dfrtp_2 _26643_ (.CLK(B_in_serial_clk),
    .D(_00446_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[45] ));
 sky130_fd_sc_hd__dfrtp_2 _26644_ (.CLK(B_in_serial_clk),
    .D(_00447_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[46] ));
 sky130_fd_sc_hd__dfrtp_2 _26645_ (.CLK(B_in_serial_clk),
    .D(_00448_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[47] ));
 sky130_fd_sc_hd__dfrtp_2 _26646_ (.CLK(B_in_serial_clk),
    .D(_00449_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[48] ));
 sky130_fd_sc_hd__dfrtp_2 _26647_ (.CLK(B_in_serial_clk),
    .D(_00450_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[49] ));
 sky130_fd_sc_hd__dfrtp_2 _26648_ (.CLK(B_in_serial_clk),
    .D(_00451_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[50] ));
 sky130_fd_sc_hd__dfrtp_2 _26649_ (.CLK(B_in_serial_clk),
    .D(_00452_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[51] ));
 sky130_fd_sc_hd__dfrtp_2 _26650_ (.CLK(B_in_serial_clk),
    .D(_00453_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[52] ));
 sky130_fd_sc_hd__dfrtp_2 _26651_ (.CLK(B_in_serial_clk),
    .D(_00454_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[53] ));
 sky130_fd_sc_hd__dfrtp_2 _26652_ (.CLK(B_in_serial_clk),
    .D(_00455_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[54] ));
 sky130_fd_sc_hd__dfrtp_2 _26653_ (.CLK(B_in_serial_clk),
    .D(_00456_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[55] ));
 sky130_fd_sc_hd__dfrtp_2 _26654_ (.CLK(B_in_serial_clk),
    .D(_00457_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[56] ));
 sky130_fd_sc_hd__dfrtp_2 _26655_ (.CLK(B_in_serial_clk),
    .D(_00458_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[57] ));
 sky130_fd_sc_hd__dfrtp_2 _26656_ (.CLK(B_in_serial_clk),
    .D(_00459_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[58] ));
 sky130_fd_sc_hd__dfrtp_2 _26657_ (.CLK(B_in_serial_clk),
    .D(_00460_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[59] ));
 sky130_fd_sc_hd__dfrtp_2 _26658_ (.CLK(B_in_serial_clk),
    .D(_00461_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[60] ));
 sky130_fd_sc_hd__dfrtp_2 _26659_ (.CLK(B_in_serial_clk),
    .D(_00462_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[61] ));
 sky130_fd_sc_hd__dfrtp_2 _26660_ (.CLK(B_in_serial_clk),
    .D(_00463_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[62] ));
 sky130_fd_sc_hd__dfrtp_2 _26661_ (.CLK(B_in_serial_clk),
    .D(_00464_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[63] ));
 sky130_fd_sc_hd__dfrtp_2 _26662_ (.CLK(B_in_serial_clk),
    .D(_00465_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[64] ));
 sky130_fd_sc_hd__dfrtp_2 _26663_ (.CLK(B_in_serial_clk),
    .D(_00466_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[65] ));
 sky130_fd_sc_hd__dfrtp_2 _26664_ (.CLK(B_in_serial_clk),
    .D(_00467_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[66] ));
 sky130_fd_sc_hd__dfrtp_2 _26665_ (.CLK(B_in_serial_clk),
    .D(_00468_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[67] ));
 sky130_fd_sc_hd__dfrtp_2 _26666_ (.CLK(B_in_serial_clk),
    .D(_00469_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[68] ));
 sky130_fd_sc_hd__dfrtp_2 _26667_ (.CLK(B_in_serial_clk),
    .D(_00470_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[69] ));
 sky130_fd_sc_hd__dfrtp_2 _26668_ (.CLK(B_in_serial_clk),
    .D(_00471_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[70] ));
 sky130_fd_sc_hd__dfrtp_2 _26669_ (.CLK(B_in_serial_clk),
    .D(_00472_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[71] ));
 sky130_fd_sc_hd__dfrtp_2 _26670_ (.CLK(B_in_serial_clk),
    .D(_00473_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[72] ));
 sky130_fd_sc_hd__dfrtp_2 _26671_ (.CLK(B_in_serial_clk),
    .D(_00474_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[73] ));
 sky130_fd_sc_hd__dfrtp_2 _26672_ (.CLK(B_in_serial_clk),
    .D(_00475_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[74] ));
 sky130_fd_sc_hd__dfrtp_2 _26673_ (.CLK(B_in_serial_clk),
    .D(_00476_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[75] ));
 sky130_fd_sc_hd__dfrtp_2 _26674_ (.CLK(B_in_serial_clk),
    .D(_00477_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[76] ));
 sky130_fd_sc_hd__dfrtp_2 _26675_ (.CLK(B_in_serial_clk),
    .D(_00478_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[77] ));
 sky130_fd_sc_hd__dfrtp_2 _26676_ (.CLK(B_in_serial_clk),
    .D(_00479_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[78] ));
 sky130_fd_sc_hd__dfrtp_2 _26677_ (.CLK(B_in_serial_clk),
    .D(_00480_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[79] ));
 sky130_fd_sc_hd__dfrtp_2 _26678_ (.CLK(B_in_serial_clk),
    .D(_00481_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[80] ));
 sky130_fd_sc_hd__dfrtp_2 _26679_ (.CLK(B_in_serial_clk),
    .D(_00482_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[81] ));
 sky130_fd_sc_hd__dfrtp_2 _26680_ (.CLK(B_in_serial_clk),
    .D(_00483_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[82] ));
 sky130_fd_sc_hd__dfrtp_2 _26681_ (.CLK(B_in_serial_clk),
    .D(_00484_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[83] ));
 sky130_fd_sc_hd__dfrtp_2 _26682_ (.CLK(B_in_serial_clk),
    .D(_00485_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[84] ));
 sky130_fd_sc_hd__dfrtp_2 _26683_ (.CLK(B_in_serial_clk),
    .D(_00486_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[85] ));
 sky130_fd_sc_hd__dfrtp_2 _26684_ (.CLK(B_in_serial_clk),
    .D(_00487_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[86] ));
 sky130_fd_sc_hd__dfrtp_2 _26685_ (.CLK(B_in_serial_clk),
    .D(_00488_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[87] ));
 sky130_fd_sc_hd__dfrtp_2 _26686_ (.CLK(B_in_serial_clk),
    .D(_00489_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[88] ));
 sky130_fd_sc_hd__dfrtp_2 _26687_ (.CLK(B_in_serial_clk),
    .D(_00490_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[89] ));
 sky130_fd_sc_hd__dfrtp_2 _26688_ (.CLK(B_in_serial_clk),
    .D(_00491_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[90] ));
 sky130_fd_sc_hd__dfrtp_2 _26689_ (.CLK(B_in_serial_clk),
    .D(_00492_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[91] ));
 sky130_fd_sc_hd__dfrtp_2 _26690_ (.CLK(B_in_serial_clk),
    .D(_00493_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[92] ));
 sky130_fd_sc_hd__dfrtp_2 _26691_ (.CLK(B_in_serial_clk),
    .D(_00494_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[93] ));
 sky130_fd_sc_hd__dfrtp_2 _26692_ (.CLK(B_in_serial_clk),
    .D(_00495_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[94] ));
 sky130_fd_sc_hd__dfrtp_2 _26693_ (.CLK(B_in_serial_clk),
    .D(_00496_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[95] ));
 sky130_fd_sc_hd__dfrtp_2 _26694_ (.CLK(B_in_serial_clk),
    .D(_00497_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[96] ));
 sky130_fd_sc_hd__dfrtp_2 _26695_ (.CLK(B_in_serial_clk),
    .D(_00498_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[97] ));
 sky130_fd_sc_hd__dfrtp_2 _26696_ (.CLK(B_in_serial_clk),
    .D(_00499_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[98] ));
 sky130_fd_sc_hd__dfrtp_2 _26697_ (.CLK(B_in_serial_clk),
    .D(_00500_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[99] ));
 sky130_fd_sc_hd__dfrtp_2 _26698_ (.CLK(B_in_serial_clk),
    .D(_00501_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[100] ));
 sky130_fd_sc_hd__dfrtp_2 _26699_ (.CLK(B_in_serial_clk),
    .D(_00502_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[101] ));
 sky130_fd_sc_hd__dfrtp_2 _26700_ (.CLK(B_in_serial_clk),
    .D(_00503_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[102] ));
 sky130_fd_sc_hd__dfrtp_2 _26701_ (.CLK(B_in_serial_clk),
    .D(_00504_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[103] ));
 sky130_fd_sc_hd__dfrtp_2 _26702_ (.CLK(B_in_serial_clk),
    .D(_00505_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[104] ));
 sky130_fd_sc_hd__dfrtp_2 _26703_ (.CLK(B_in_serial_clk),
    .D(_00506_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[105] ));
 sky130_fd_sc_hd__dfrtp_2 _26704_ (.CLK(B_in_serial_clk),
    .D(_00507_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[106] ));
 sky130_fd_sc_hd__dfrtp_2 _26705_ (.CLK(B_in_serial_clk),
    .D(_00508_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[107] ));
 sky130_fd_sc_hd__dfrtp_2 _26706_ (.CLK(B_in_serial_clk),
    .D(_00509_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[108] ));
 sky130_fd_sc_hd__dfrtp_2 _26707_ (.CLK(B_in_serial_clk),
    .D(_00510_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[109] ));
 sky130_fd_sc_hd__dfrtp_2 _26708_ (.CLK(B_in_serial_clk),
    .D(_00511_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[110] ));
 sky130_fd_sc_hd__dfrtp_2 _26709_ (.CLK(B_in_serial_clk),
    .D(_00512_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[111] ));
 sky130_fd_sc_hd__dfrtp_2 _26710_ (.CLK(B_in_serial_clk),
    .D(_00513_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[112] ));
 sky130_fd_sc_hd__dfrtp_2 _26711_ (.CLK(B_in_serial_clk),
    .D(_00514_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[113] ));
 sky130_fd_sc_hd__dfrtp_2 _26712_ (.CLK(B_in_serial_clk),
    .D(_00515_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[114] ));
 sky130_fd_sc_hd__dfrtp_2 _26713_ (.CLK(B_in_serial_clk),
    .D(_00516_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[115] ));
 sky130_fd_sc_hd__dfrtp_2 _26714_ (.CLK(B_in_serial_clk),
    .D(_00517_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[116] ));
 sky130_fd_sc_hd__dfrtp_2 _26715_ (.CLK(B_in_serial_clk),
    .D(_00518_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[117] ));
 sky130_fd_sc_hd__dfrtp_2 _26716_ (.CLK(B_in_serial_clk),
    .D(_00519_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[118] ));
 sky130_fd_sc_hd__dfrtp_2 _26717_ (.CLK(B_in_serial_clk),
    .D(_00520_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[119] ));
 sky130_fd_sc_hd__dfrtp_2 _26718_ (.CLK(B_in_serial_clk),
    .D(_00521_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[120] ));
 sky130_fd_sc_hd__dfrtp_2 _26719_ (.CLK(B_in_serial_clk),
    .D(_00522_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[121] ));
 sky130_fd_sc_hd__dfrtp_2 _26720_ (.CLK(B_in_serial_clk),
    .D(_00523_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[122] ));
 sky130_fd_sc_hd__dfrtp_2 _26721_ (.CLK(B_in_serial_clk),
    .D(_00524_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[123] ));
 sky130_fd_sc_hd__dfrtp_2 _26722_ (.CLK(B_in_serial_clk),
    .D(_00525_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[124] ));
 sky130_fd_sc_hd__dfrtp_2 _26723_ (.CLK(B_in_serial_clk),
    .D(_00526_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[125] ));
 sky130_fd_sc_hd__dfrtp_2 _26724_ (.CLK(B_in_serial_clk),
    .D(_00527_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[126] ));
 sky130_fd_sc_hd__dfrtp_2 _26725_ (.CLK(B_in_serial_clk),
    .D(_00528_),
    .RESET_B(rst_n),
    .Q(\deser_B.word_buffer[127] ));
 sky130_fd_sc_hd__dfrtp_2 _26726_ (.CLK(B_in_serial_clk),
    .D(_00006_),
    .RESET_B(rst_n),
    .Q(\deser_B.receiving ));
 sky130_fd_sc_hd__dfrtp_2 _26727_ (.CLK(B_in_serial_clk),
    .D(_00529_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_toggle ));
 sky130_fd_sc_hd__dfrtp_2 _26728_ (.CLK(clk),
    .D(_00530_),
    .RESET_B(rst_n),
    .Q(\B_in[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26729_ (.CLK(clk),
    .D(_00531_),
    .RESET_B(rst_n),
    .Q(\B_in[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26730_ (.CLK(clk),
    .D(_00532_),
    .RESET_B(rst_n),
    .Q(\B_in[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26731_ (.CLK(clk),
    .D(_00533_),
    .RESET_B(rst_n),
    .Q(\B_in[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26732_ (.CLK(clk),
    .D(_00534_),
    .RESET_B(rst_n),
    .Q(\B_in[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26733_ (.CLK(clk),
    .D(_00535_),
    .RESET_B(rst_n),
    .Q(\B_in[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26734_ (.CLK(clk),
    .D(_00536_),
    .RESET_B(rst_n),
    .Q(\B_in[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26735_ (.CLK(clk),
    .D(_00537_),
    .RESET_B(rst_n),
    .Q(\B_in[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26736_ (.CLK(clk),
    .D(_00538_),
    .RESET_B(rst_n),
    .Q(\B_in[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26737_ (.CLK(clk),
    .D(_00539_),
    .RESET_B(rst_n),
    .Q(\B_in[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26738_ (.CLK(clk),
    .D(_00540_),
    .RESET_B(rst_n),
    .Q(\B_in[10] ));
 sky130_fd_sc_hd__dfrtp_2 _26739_ (.CLK(clk),
    .D(_00541_),
    .RESET_B(rst_n),
    .Q(\B_in[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26740_ (.CLK(clk),
    .D(_00542_),
    .RESET_B(rst_n),
    .Q(\B_in[12] ));
 sky130_fd_sc_hd__dfrtp_2 _26741_ (.CLK(clk),
    .D(_00543_),
    .RESET_B(rst_n),
    .Q(\B_in[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26742_ (.CLK(clk),
    .D(_00544_),
    .RESET_B(rst_n),
    .Q(\B_in[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26743_ (.CLK(clk),
    .D(_00545_),
    .RESET_B(rst_n),
    .Q(\B_in[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26744_ (.CLK(clk),
    .D(_00546_),
    .RESET_B(rst_n),
    .Q(\B_in[16] ));
 sky130_fd_sc_hd__dfrtp_2 _26745_ (.CLK(clk),
    .D(_00547_),
    .RESET_B(rst_n),
    .Q(\B_in[17] ));
 sky130_fd_sc_hd__dfrtp_2 _26746_ (.CLK(clk),
    .D(_00548_),
    .RESET_B(rst_n),
    .Q(\B_in[18] ));
 sky130_fd_sc_hd__dfrtp_2 _26747_ (.CLK(clk),
    .D(_00549_),
    .RESET_B(rst_n),
    .Q(\B_in[19] ));
 sky130_fd_sc_hd__dfrtp_2 _26748_ (.CLK(clk),
    .D(_00550_),
    .RESET_B(rst_n),
    .Q(\B_in[20] ));
 sky130_fd_sc_hd__dfrtp_2 _26749_ (.CLK(clk),
    .D(_00551_),
    .RESET_B(rst_n),
    .Q(\B_in[21] ));
 sky130_fd_sc_hd__dfrtp_2 _26750_ (.CLK(clk),
    .D(_00552_),
    .RESET_B(rst_n),
    .Q(\B_in[22] ));
 sky130_fd_sc_hd__dfrtp_2 _26751_ (.CLK(clk),
    .D(_00553_),
    .RESET_B(rst_n),
    .Q(\B_in[23] ));
 sky130_fd_sc_hd__dfrtp_2 _26752_ (.CLK(clk),
    .D(_00554_),
    .RESET_B(rst_n),
    .Q(\B_in[24] ));
 sky130_fd_sc_hd__dfrtp_2 _26753_ (.CLK(clk),
    .D(_00555_),
    .RESET_B(rst_n),
    .Q(\B_in[25] ));
 sky130_fd_sc_hd__dfrtp_2 _26754_ (.CLK(clk),
    .D(_00556_),
    .RESET_B(rst_n),
    .Q(\B_in[26] ));
 sky130_fd_sc_hd__dfrtp_2 _26755_ (.CLK(clk),
    .D(_00557_),
    .RESET_B(rst_n),
    .Q(\B_in[27] ));
 sky130_fd_sc_hd__dfrtp_2 _26756_ (.CLK(clk),
    .D(_00558_),
    .RESET_B(rst_n),
    .Q(\B_in[28] ));
 sky130_fd_sc_hd__dfrtp_2 _26757_ (.CLK(clk),
    .D(_00559_),
    .RESET_B(rst_n),
    .Q(\B_in[29] ));
 sky130_fd_sc_hd__dfrtp_2 _26758_ (.CLK(clk),
    .D(_00560_),
    .RESET_B(rst_n),
    .Q(\B_in[30] ));
 sky130_fd_sc_hd__dfrtp_2 _26759_ (.CLK(clk),
    .D(_00561_),
    .RESET_B(rst_n),
    .Q(\B_in[31] ));
 sky130_fd_sc_hd__dfrtp_2 _26760_ (.CLK(clk),
    .D(_00562_),
    .RESET_B(rst_n),
    .Q(\B_in[32] ));
 sky130_fd_sc_hd__dfrtp_2 _26761_ (.CLK(clk),
    .D(_00563_),
    .RESET_B(rst_n),
    .Q(\B_in[33] ));
 sky130_fd_sc_hd__dfrtp_2 _26762_ (.CLK(clk),
    .D(_00564_),
    .RESET_B(rst_n),
    .Q(\B_in[34] ));
 sky130_fd_sc_hd__dfrtp_2 _26763_ (.CLK(clk),
    .D(_00565_),
    .RESET_B(rst_n),
    .Q(\B_in[35] ));
 sky130_fd_sc_hd__dfrtp_2 _26764_ (.CLK(clk),
    .D(_00566_),
    .RESET_B(rst_n),
    .Q(\B_in[36] ));
 sky130_fd_sc_hd__dfrtp_2 _26765_ (.CLK(clk),
    .D(_00567_),
    .RESET_B(rst_n),
    .Q(\B_in[37] ));
 sky130_fd_sc_hd__dfrtp_2 _26766_ (.CLK(clk),
    .D(_00568_),
    .RESET_B(rst_n),
    .Q(\B_in[38] ));
 sky130_fd_sc_hd__dfrtp_2 _26767_ (.CLK(clk),
    .D(_00569_),
    .RESET_B(rst_n),
    .Q(\B_in[39] ));
 sky130_fd_sc_hd__dfrtp_2 _26768_ (.CLK(clk),
    .D(_00570_),
    .RESET_B(rst_n),
    .Q(\B_in[40] ));
 sky130_fd_sc_hd__dfrtp_2 _26769_ (.CLK(clk),
    .D(_00571_),
    .RESET_B(rst_n),
    .Q(\B_in[41] ));
 sky130_fd_sc_hd__dfrtp_2 _26770_ (.CLK(clk),
    .D(_00572_),
    .RESET_B(rst_n),
    .Q(\B_in[42] ));
 sky130_fd_sc_hd__dfrtp_2 _26771_ (.CLK(clk),
    .D(_00573_),
    .RESET_B(rst_n),
    .Q(\B_in[43] ));
 sky130_fd_sc_hd__dfrtp_2 _26772_ (.CLK(clk),
    .D(_00574_),
    .RESET_B(rst_n),
    .Q(\B_in[44] ));
 sky130_fd_sc_hd__dfrtp_2 _26773_ (.CLK(clk),
    .D(_00575_),
    .RESET_B(rst_n),
    .Q(\B_in[45] ));
 sky130_fd_sc_hd__dfrtp_2 _26774_ (.CLK(clk),
    .D(_00576_),
    .RESET_B(rst_n),
    .Q(\B_in[46] ));
 sky130_fd_sc_hd__dfrtp_2 _26775_ (.CLK(clk),
    .D(_00577_),
    .RESET_B(rst_n),
    .Q(\B_in[47] ));
 sky130_fd_sc_hd__dfrtp_2 _26776_ (.CLK(clk),
    .D(_00578_),
    .RESET_B(rst_n),
    .Q(\B_in[48] ));
 sky130_fd_sc_hd__dfrtp_2 _26777_ (.CLK(clk),
    .D(_00579_),
    .RESET_B(rst_n),
    .Q(\B_in[49] ));
 sky130_fd_sc_hd__dfrtp_2 _26778_ (.CLK(clk),
    .D(_00580_),
    .RESET_B(rst_n),
    .Q(\B_in[50] ));
 sky130_fd_sc_hd__dfrtp_2 _26779_ (.CLK(clk),
    .D(_00581_),
    .RESET_B(rst_n),
    .Q(\B_in[51] ));
 sky130_fd_sc_hd__dfrtp_2 _26780_ (.CLK(clk),
    .D(_00582_),
    .RESET_B(rst_n),
    .Q(\B_in[52] ));
 sky130_fd_sc_hd__dfrtp_2 _26781_ (.CLK(clk),
    .D(_00583_),
    .RESET_B(rst_n),
    .Q(\B_in[53] ));
 sky130_fd_sc_hd__dfrtp_2 _26782_ (.CLK(clk),
    .D(_00584_),
    .RESET_B(rst_n),
    .Q(\B_in[54] ));
 sky130_fd_sc_hd__dfrtp_2 _26783_ (.CLK(clk),
    .D(_00585_),
    .RESET_B(rst_n),
    .Q(\B_in[55] ));
 sky130_fd_sc_hd__dfrtp_2 _26784_ (.CLK(clk),
    .D(_00586_),
    .RESET_B(rst_n),
    .Q(\B_in[56] ));
 sky130_fd_sc_hd__dfrtp_2 _26785_ (.CLK(clk),
    .D(_00587_),
    .RESET_B(rst_n),
    .Q(\B_in[57] ));
 sky130_fd_sc_hd__dfrtp_2 _26786_ (.CLK(clk),
    .D(_00588_),
    .RESET_B(rst_n),
    .Q(\B_in[58] ));
 sky130_fd_sc_hd__dfrtp_2 _26787_ (.CLK(clk),
    .D(_00589_),
    .RESET_B(rst_n),
    .Q(\B_in[59] ));
 sky130_fd_sc_hd__dfrtp_2 _26788_ (.CLK(clk),
    .D(_00590_),
    .RESET_B(rst_n),
    .Q(\B_in[60] ));
 sky130_fd_sc_hd__dfrtp_2 _26789_ (.CLK(clk),
    .D(_00591_),
    .RESET_B(rst_n),
    .Q(\B_in[61] ));
 sky130_fd_sc_hd__dfrtp_2 _26790_ (.CLK(clk),
    .D(_00592_),
    .RESET_B(rst_n),
    .Q(\B_in[62] ));
 sky130_fd_sc_hd__dfrtp_2 _26791_ (.CLK(clk),
    .D(_00593_),
    .RESET_B(rst_n),
    .Q(\B_in[63] ));
 sky130_fd_sc_hd__dfrtp_2 _26792_ (.CLK(clk),
    .D(_00594_),
    .RESET_B(rst_n),
    .Q(\B_in[64] ));
 sky130_fd_sc_hd__dfrtp_2 _26793_ (.CLK(clk),
    .D(_00595_),
    .RESET_B(rst_n),
    .Q(\B_in[65] ));
 sky130_fd_sc_hd__dfrtp_2 _26794_ (.CLK(clk),
    .D(_00596_),
    .RESET_B(rst_n),
    .Q(\B_in[66] ));
 sky130_fd_sc_hd__dfrtp_2 _26795_ (.CLK(clk),
    .D(_00597_),
    .RESET_B(rst_n),
    .Q(\B_in[67] ));
 sky130_fd_sc_hd__dfrtp_2 _26796_ (.CLK(clk),
    .D(_00598_),
    .RESET_B(rst_n),
    .Q(\B_in[68] ));
 sky130_fd_sc_hd__dfrtp_2 _26797_ (.CLK(clk),
    .D(_00599_),
    .RESET_B(rst_n),
    .Q(\B_in[69] ));
 sky130_fd_sc_hd__dfrtp_2 _26798_ (.CLK(clk),
    .D(_00600_),
    .RESET_B(rst_n),
    .Q(\B_in[70] ));
 sky130_fd_sc_hd__dfrtp_2 _26799_ (.CLK(clk),
    .D(_00601_),
    .RESET_B(rst_n),
    .Q(\B_in[71] ));
 sky130_fd_sc_hd__dfrtp_2 _26800_ (.CLK(clk),
    .D(_00602_),
    .RESET_B(rst_n),
    .Q(\B_in[72] ));
 sky130_fd_sc_hd__dfrtp_2 _26801_ (.CLK(clk),
    .D(_00603_),
    .RESET_B(rst_n),
    .Q(\B_in[73] ));
 sky130_fd_sc_hd__dfrtp_2 _26802_ (.CLK(clk),
    .D(_00604_),
    .RESET_B(rst_n),
    .Q(\B_in[74] ));
 sky130_fd_sc_hd__dfrtp_2 _26803_ (.CLK(clk),
    .D(_00605_),
    .RESET_B(rst_n),
    .Q(\B_in[75] ));
 sky130_fd_sc_hd__dfrtp_2 _26804_ (.CLK(clk),
    .D(_00606_),
    .RESET_B(rst_n),
    .Q(\B_in[76] ));
 sky130_fd_sc_hd__dfrtp_2 _26805_ (.CLK(clk),
    .D(_00607_),
    .RESET_B(rst_n),
    .Q(\B_in[77] ));
 sky130_fd_sc_hd__dfrtp_2 _26806_ (.CLK(clk),
    .D(_00608_),
    .RESET_B(rst_n),
    .Q(\B_in[78] ));
 sky130_fd_sc_hd__dfrtp_2 _26807_ (.CLK(clk),
    .D(_00609_),
    .RESET_B(rst_n),
    .Q(\B_in[79] ));
 sky130_fd_sc_hd__dfrtp_2 _26808_ (.CLK(clk),
    .D(_00610_),
    .RESET_B(rst_n),
    .Q(\B_in[80] ));
 sky130_fd_sc_hd__dfrtp_2 _26809_ (.CLK(clk),
    .D(_00611_),
    .RESET_B(rst_n),
    .Q(\B_in[81] ));
 sky130_fd_sc_hd__dfrtp_2 _26810_ (.CLK(clk),
    .D(_00612_),
    .RESET_B(rst_n),
    .Q(\B_in[82] ));
 sky130_fd_sc_hd__dfrtp_2 _26811_ (.CLK(clk),
    .D(_00613_),
    .RESET_B(rst_n),
    .Q(\B_in[83] ));
 sky130_fd_sc_hd__dfrtp_2 _26812_ (.CLK(clk),
    .D(_00614_),
    .RESET_B(rst_n),
    .Q(\B_in[84] ));
 sky130_fd_sc_hd__dfrtp_2 _26813_ (.CLK(clk),
    .D(_00615_),
    .RESET_B(rst_n),
    .Q(\B_in[85] ));
 sky130_fd_sc_hd__dfrtp_2 _26814_ (.CLK(clk),
    .D(_00616_),
    .RESET_B(rst_n),
    .Q(\B_in[86] ));
 sky130_fd_sc_hd__dfrtp_2 _26815_ (.CLK(clk),
    .D(_00617_),
    .RESET_B(rst_n),
    .Q(\B_in[87] ));
 sky130_fd_sc_hd__dfrtp_2 _26816_ (.CLK(clk),
    .D(_00618_),
    .RESET_B(rst_n),
    .Q(\B_in[88] ));
 sky130_fd_sc_hd__dfrtp_2 _26817_ (.CLK(clk),
    .D(_00619_),
    .RESET_B(rst_n),
    .Q(\B_in[89] ));
 sky130_fd_sc_hd__dfrtp_2 _26818_ (.CLK(clk),
    .D(_00620_),
    .RESET_B(rst_n),
    .Q(\B_in[90] ));
 sky130_fd_sc_hd__dfrtp_2 _26819_ (.CLK(clk),
    .D(_00621_),
    .RESET_B(rst_n),
    .Q(\B_in[91] ));
 sky130_fd_sc_hd__dfrtp_2 _26820_ (.CLK(clk),
    .D(_00622_),
    .RESET_B(rst_n),
    .Q(\B_in[92] ));
 sky130_fd_sc_hd__dfrtp_2 _26821_ (.CLK(clk),
    .D(_00623_),
    .RESET_B(rst_n),
    .Q(\B_in[93] ));
 sky130_fd_sc_hd__dfrtp_2 _26822_ (.CLK(clk),
    .D(_00624_),
    .RESET_B(rst_n),
    .Q(\B_in[94] ));
 sky130_fd_sc_hd__dfrtp_2 _26823_ (.CLK(clk),
    .D(_00625_),
    .RESET_B(rst_n),
    .Q(\B_in[95] ));
 sky130_fd_sc_hd__dfrtp_2 _26824_ (.CLK(clk),
    .D(_00626_),
    .RESET_B(rst_n),
    .Q(\B_in[96] ));
 sky130_fd_sc_hd__dfrtp_2 _26825_ (.CLK(clk),
    .D(_00627_),
    .RESET_B(rst_n),
    .Q(\B_in[97] ));
 sky130_fd_sc_hd__dfrtp_2 _26826_ (.CLK(clk),
    .D(_00628_),
    .RESET_B(rst_n),
    .Q(\B_in[98] ));
 sky130_fd_sc_hd__dfrtp_2 _26827_ (.CLK(clk),
    .D(_00629_),
    .RESET_B(rst_n),
    .Q(\B_in[99] ));
 sky130_fd_sc_hd__dfrtp_2 _26828_ (.CLK(clk),
    .D(_00630_),
    .RESET_B(rst_n),
    .Q(\B_in[100] ));
 sky130_fd_sc_hd__dfrtp_2 _26829_ (.CLK(clk),
    .D(_00631_),
    .RESET_B(rst_n),
    .Q(\B_in[101] ));
 sky130_fd_sc_hd__dfrtp_2 _26830_ (.CLK(clk),
    .D(_00632_),
    .RESET_B(rst_n),
    .Q(\B_in[102] ));
 sky130_fd_sc_hd__dfrtp_2 _26831_ (.CLK(clk),
    .D(_00633_),
    .RESET_B(rst_n),
    .Q(\B_in[103] ));
 sky130_fd_sc_hd__dfrtp_2 _26832_ (.CLK(clk),
    .D(_00634_),
    .RESET_B(rst_n),
    .Q(\B_in[104] ));
 sky130_fd_sc_hd__dfrtp_2 _26833_ (.CLK(clk),
    .D(_00635_),
    .RESET_B(rst_n),
    .Q(\B_in[105] ));
 sky130_fd_sc_hd__dfrtp_2 _26834_ (.CLK(clk),
    .D(_00636_),
    .RESET_B(rst_n),
    .Q(\B_in[106] ));
 sky130_fd_sc_hd__dfrtp_2 _26835_ (.CLK(clk),
    .D(_00637_),
    .RESET_B(rst_n),
    .Q(\B_in[107] ));
 sky130_fd_sc_hd__dfrtp_2 _26836_ (.CLK(clk),
    .D(_00638_),
    .RESET_B(rst_n),
    .Q(\B_in[108] ));
 sky130_fd_sc_hd__dfrtp_2 _26837_ (.CLK(clk),
    .D(_00639_),
    .RESET_B(rst_n),
    .Q(\B_in[109] ));
 sky130_fd_sc_hd__dfrtp_2 _26838_ (.CLK(clk),
    .D(_00640_),
    .RESET_B(rst_n),
    .Q(\B_in[110] ));
 sky130_fd_sc_hd__dfrtp_2 _26839_ (.CLK(clk),
    .D(_00641_),
    .RESET_B(rst_n),
    .Q(\B_in[111] ));
 sky130_fd_sc_hd__dfrtp_2 _26840_ (.CLK(clk),
    .D(_00642_),
    .RESET_B(rst_n),
    .Q(\B_in[112] ));
 sky130_fd_sc_hd__dfrtp_2 _26841_ (.CLK(clk),
    .D(_00643_),
    .RESET_B(rst_n),
    .Q(\B_in[113] ));
 sky130_fd_sc_hd__dfrtp_2 _26842_ (.CLK(clk),
    .D(_00644_),
    .RESET_B(rst_n),
    .Q(\B_in[114] ));
 sky130_fd_sc_hd__dfrtp_2 _26843_ (.CLK(clk),
    .D(_00645_),
    .RESET_B(rst_n),
    .Q(\B_in[115] ));
 sky130_fd_sc_hd__dfrtp_2 _26844_ (.CLK(clk),
    .D(_00646_),
    .RESET_B(rst_n),
    .Q(\B_in[116] ));
 sky130_fd_sc_hd__dfrtp_2 _26845_ (.CLK(clk),
    .D(_00647_),
    .RESET_B(rst_n),
    .Q(\B_in[117] ));
 sky130_fd_sc_hd__dfrtp_2 _26846_ (.CLK(clk),
    .D(_00648_),
    .RESET_B(rst_n),
    .Q(\B_in[118] ));
 sky130_fd_sc_hd__dfrtp_2 _26847_ (.CLK(clk),
    .D(_00649_),
    .RESET_B(rst_n),
    .Q(\B_in[119] ));
 sky130_fd_sc_hd__dfrtp_2 _26848_ (.CLK(clk),
    .D(_00650_),
    .RESET_B(rst_n),
    .Q(\B_in[120] ));
 sky130_fd_sc_hd__dfrtp_2 _26849_ (.CLK(clk),
    .D(_00651_),
    .RESET_B(rst_n),
    .Q(\B_in[121] ));
 sky130_fd_sc_hd__dfrtp_2 _26850_ (.CLK(clk),
    .D(_00652_),
    .RESET_B(rst_n),
    .Q(\B_in[122] ));
 sky130_fd_sc_hd__dfrtp_2 _26851_ (.CLK(clk),
    .D(_00653_),
    .RESET_B(rst_n),
    .Q(\B_in[123] ));
 sky130_fd_sc_hd__dfrtp_2 _26852_ (.CLK(clk),
    .D(_00654_),
    .RESET_B(rst_n),
    .Q(\B_in[124] ));
 sky130_fd_sc_hd__dfrtp_2 _26853_ (.CLK(clk),
    .D(_00655_),
    .RESET_B(rst_n),
    .Q(\B_in[125] ));
 sky130_fd_sc_hd__dfrtp_2 _26854_ (.CLK(clk),
    .D(_00656_),
    .RESET_B(rst_n),
    .Q(\B_in[126] ));
 sky130_fd_sc_hd__dfrtp_2 _26855_ (.CLK(clk),
    .D(_00657_),
    .RESET_B(rst_n),
    .Q(\B_in[127] ));
 sky130_fd_sc_hd__dfrtp_2 _26856_ (.CLK(B_in_serial_clk),
    .D(_00658_),
    .RESET_B(rst_n),
    .Q(\deser_B.bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26857_ (.CLK(B_in_serial_clk),
    .D(_00659_),
    .RESET_B(rst_n),
    .Q(\deser_B.bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26858_ (.CLK(B_in_serial_clk),
    .D(_00660_),
    .RESET_B(rst_n),
    .Q(\deser_B.bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26859_ (.CLK(B_in_serial_clk),
    .D(_00661_),
    .RESET_B(rst_n),
    .Q(\deser_B.bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26860_ (.CLK(B_in_serial_clk),
    .D(_00662_),
    .RESET_B(rst_n),
    .Q(\deser_B.bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26861_ (.CLK(B_in_serial_clk),
    .D(_00663_),
    .RESET_B(rst_n),
    .Q(\deser_B.bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26862_ (.CLK(B_in_serial_clk),
    .D(_00664_),
    .RESET_B(rst_n),
    .Q(\deser_B.bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26863_ (.CLK(clk),
    .D(\deser_B.serial_toggle_sync1 ),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_toggle_sync2 ));
 sky130_fd_sc_hd__dfrtp_2 _26864_ (.CLK(B_in_serial_clk),
    .D(_00001_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word_ready ));
 sky130_fd_sc_hd__dfrtp_2 _26865_ (.CLK(clk),
    .D(\deser_B.serial_toggle ),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_toggle_sync1 ));
 sky130_fd_sc_hd__dfrtp_2 _26866_ (.CLK(clk),
    .D(_00005_),
    .RESET_B(rst_n),
    .Q(B_in_valid));
 sky130_fd_sc_hd__dfrtp_2 _26867_ (.CLK(A_in_serial_clk),
    .D(_00665_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26868_ (.CLK(A_in_serial_clk),
    .D(_00666_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26869_ (.CLK(A_in_serial_clk),
    .D(_00667_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26870_ (.CLK(A_in_serial_clk),
    .D(_00668_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26871_ (.CLK(A_in_serial_clk),
    .D(_00669_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26872_ (.CLK(A_in_serial_clk),
    .D(_00670_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26873_ (.CLK(A_in_serial_clk),
    .D(_00671_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26874_ (.CLK(A_in_serial_clk),
    .D(_00672_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26875_ (.CLK(A_in_serial_clk),
    .D(_00673_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26876_ (.CLK(A_in_serial_clk),
    .D(_00674_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26877_ (.CLK(A_in_serial_clk),
    .D(_00675_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[10] ));
 sky130_fd_sc_hd__dfrtp_2 _26878_ (.CLK(A_in_serial_clk),
    .D(_00676_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26879_ (.CLK(A_in_serial_clk),
    .D(_00677_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[12] ));
 sky130_fd_sc_hd__dfrtp_2 _26880_ (.CLK(A_in_serial_clk),
    .D(_00678_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26881_ (.CLK(A_in_serial_clk),
    .D(_00679_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26882_ (.CLK(A_in_serial_clk),
    .D(_00680_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26883_ (.CLK(A_in_serial_clk),
    .D(_00681_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[16] ));
 sky130_fd_sc_hd__dfrtp_2 _26884_ (.CLK(A_in_serial_clk),
    .D(_00682_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[17] ));
 sky130_fd_sc_hd__dfrtp_2 _26885_ (.CLK(A_in_serial_clk),
    .D(_00683_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[18] ));
 sky130_fd_sc_hd__dfrtp_2 _26886_ (.CLK(A_in_serial_clk),
    .D(_00684_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[19] ));
 sky130_fd_sc_hd__dfrtp_2 _26887_ (.CLK(A_in_serial_clk),
    .D(_00685_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[20] ));
 sky130_fd_sc_hd__dfrtp_2 _26888_ (.CLK(A_in_serial_clk),
    .D(_00686_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[21] ));
 sky130_fd_sc_hd__dfrtp_2 _26889_ (.CLK(A_in_serial_clk),
    .D(_00687_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[22] ));
 sky130_fd_sc_hd__dfrtp_2 _26890_ (.CLK(A_in_serial_clk),
    .D(_00688_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[23] ));
 sky130_fd_sc_hd__dfrtp_2 _26891_ (.CLK(A_in_serial_clk),
    .D(_00689_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[24] ));
 sky130_fd_sc_hd__dfrtp_2 _26892_ (.CLK(A_in_serial_clk),
    .D(_00690_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[25] ));
 sky130_fd_sc_hd__dfrtp_2 _26893_ (.CLK(A_in_serial_clk),
    .D(_00691_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[26] ));
 sky130_fd_sc_hd__dfrtp_2 _26894_ (.CLK(A_in_serial_clk),
    .D(_00692_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[27] ));
 sky130_fd_sc_hd__dfrtp_2 _26895_ (.CLK(A_in_serial_clk),
    .D(_00693_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[28] ));
 sky130_fd_sc_hd__dfrtp_2 _26896_ (.CLK(A_in_serial_clk),
    .D(_00694_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[29] ));
 sky130_fd_sc_hd__dfrtp_2 _26897_ (.CLK(A_in_serial_clk),
    .D(_00695_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[30] ));
 sky130_fd_sc_hd__dfrtp_2 _26898_ (.CLK(A_in_serial_clk),
    .D(_00696_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[31] ));
 sky130_fd_sc_hd__dfrtp_2 _26899_ (.CLK(A_in_serial_clk),
    .D(_00697_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[32] ));
 sky130_fd_sc_hd__dfrtp_2 _26900_ (.CLK(A_in_serial_clk),
    .D(_00698_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[33] ));
 sky130_fd_sc_hd__dfrtp_2 _26901_ (.CLK(A_in_serial_clk),
    .D(_00699_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[34] ));
 sky130_fd_sc_hd__dfrtp_2 _26902_ (.CLK(A_in_serial_clk),
    .D(_00700_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[35] ));
 sky130_fd_sc_hd__dfrtp_2 _26903_ (.CLK(A_in_serial_clk),
    .D(_00701_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[36] ));
 sky130_fd_sc_hd__dfrtp_2 _26904_ (.CLK(A_in_serial_clk),
    .D(_00702_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[37] ));
 sky130_fd_sc_hd__dfrtp_2 _26905_ (.CLK(A_in_serial_clk),
    .D(_00703_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[38] ));
 sky130_fd_sc_hd__dfrtp_2 _26906_ (.CLK(A_in_serial_clk),
    .D(_00704_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[39] ));
 sky130_fd_sc_hd__dfrtp_2 _26907_ (.CLK(A_in_serial_clk),
    .D(_00705_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[40] ));
 sky130_fd_sc_hd__dfrtp_2 _26908_ (.CLK(A_in_serial_clk),
    .D(_00706_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[41] ));
 sky130_fd_sc_hd__dfrtp_2 _26909_ (.CLK(A_in_serial_clk),
    .D(_00707_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[42] ));
 sky130_fd_sc_hd__dfrtp_2 _26910_ (.CLK(A_in_serial_clk),
    .D(_00708_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[43] ));
 sky130_fd_sc_hd__dfrtp_2 _26911_ (.CLK(A_in_serial_clk),
    .D(_00709_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[44] ));
 sky130_fd_sc_hd__dfrtp_2 _26912_ (.CLK(A_in_serial_clk),
    .D(_00710_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[45] ));
 sky130_fd_sc_hd__dfrtp_2 _26913_ (.CLK(A_in_serial_clk),
    .D(_00711_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[46] ));
 sky130_fd_sc_hd__dfrtp_2 _26914_ (.CLK(A_in_serial_clk),
    .D(_00712_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[47] ));
 sky130_fd_sc_hd__dfrtp_2 _26915_ (.CLK(A_in_serial_clk),
    .D(_00713_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[48] ));
 sky130_fd_sc_hd__dfrtp_2 _26916_ (.CLK(A_in_serial_clk),
    .D(_00714_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[49] ));
 sky130_fd_sc_hd__dfrtp_2 _26917_ (.CLK(A_in_serial_clk),
    .D(_00715_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[50] ));
 sky130_fd_sc_hd__dfrtp_2 _26918_ (.CLK(A_in_serial_clk),
    .D(_00716_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[51] ));
 sky130_fd_sc_hd__dfrtp_2 _26919_ (.CLK(A_in_serial_clk),
    .D(_00717_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[52] ));
 sky130_fd_sc_hd__dfrtp_2 _26920_ (.CLK(A_in_serial_clk),
    .D(_00718_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[53] ));
 sky130_fd_sc_hd__dfrtp_2 _26921_ (.CLK(A_in_serial_clk),
    .D(_00719_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[54] ));
 sky130_fd_sc_hd__dfrtp_2 _26922_ (.CLK(A_in_serial_clk),
    .D(_00720_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[55] ));
 sky130_fd_sc_hd__dfrtp_2 _26923_ (.CLK(A_in_serial_clk),
    .D(_00721_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[56] ));
 sky130_fd_sc_hd__dfrtp_2 _26924_ (.CLK(A_in_serial_clk),
    .D(_00722_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[57] ));
 sky130_fd_sc_hd__dfrtp_2 _26925_ (.CLK(A_in_serial_clk),
    .D(_00723_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[58] ));
 sky130_fd_sc_hd__dfrtp_2 _26926_ (.CLK(A_in_serial_clk),
    .D(_00724_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[59] ));
 sky130_fd_sc_hd__dfrtp_2 _26927_ (.CLK(A_in_serial_clk),
    .D(_00725_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[60] ));
 sky130_fd_sc_hd__dfrtp_2 _26928_ (.CLK(A_in_serial_clk),
    .D(_00726_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[61] ));
 sky130_fd_sc_hd__dfrtp_2 _26929_ (.CLK(A_in_serial_clk),
    .D(_00727_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[62] ));
 sky130_fd_sc_hd__dfrtp_2 _26930_ (.CLK(A_in_serial_clk),
    .D(_00728_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[63] ));
 sky130_fd_sc_hd__dfrtp_2 _26931_ (.CLK(A_in_serial_clk),
    .D(_00729_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[64] ));
 sky130_fd_sc_hd__dfrtp_2 _26932_ (.CLK(A_in_serial_clk),
    .D(_00730_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[65] ));
 sky130_fd_sc_hd__dfrtp_2 _26933_ (.CLK(A_in_serial_clk),
    .D(_00731_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[66] ));
 sky130_fd_sc_hd__dfrtp_2 _26934_ (.CLK(A_in_serial_clk),
    .D(_00732_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[67] ));
 sky130_fd_sc_hd__dfrtp_2 _26935_ (.CLK(A_in_serial_clk),
    .D(_00733_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[68] ));
 sky130_fd_sc_hd__dfrtp_2 _26936_ (.CLK(A_in_serial_clk),
    .D(_00734_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[69] ));
 sky130_fd_sc_hd__dfrtp_2 _26937_ (.CLK(A_in_serial_clk),
    .D(_00735_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[70] ));
 sky130_fd_sc_hd__dfrtp_2 _26938_ (.CLK(A_in_serial_clk),
    .D(_00736_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[71] ));
 sky130_fd_sc_hd__dfrtp_2 _26939_ (.CLK(A_in_serial_clk),
    .D(_00737_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[72] ));
 sky130_fd_sc_hd__dfrtp_2 _26940_ (.CLK(A_in_serial_clk),
    .D(_00738_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[73] ));
 sky130_fd_sc_hd__dfrtp_2 _26941_ (.CLK(A_in_serial_clk),
    .D(_00739_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[74] ));
 sky130_fd_sc_hd__dfrtp_2 _26942_ (.CLK(A_in_serial_clk),
    .D(_00740_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[75] ));
 sky130_fd_sc_hd__dfrtp_2 _26943_ (.CLK(A_in_serial_clk),
    .D(_00741_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[76] ));
 sky130_fd_sc_hd__dfrtp_2 _26944_ (.CLK(A_in_serial_clk),
    .D(_00742_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[77] ));
 sky130_fd_sc_hd__dfrtp_2 _26945_ (.CLK(A_in_serial_clk),
    .D(_00743_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[78] ));
 sky130_fd_sc_hd__dfrtp_2 _26946_ (.CLK(A_in_serial_clk),
    .D(_00744_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[79] ));
 sky130_fd_sc_hd__dfrtp_2 _26947_ (.CLK(A_in_serial_clk),
    .D(_00745_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[80] ));
 sky130_fd_sc_hd__dfrtp_2 _26948_ (.CLK(A_in_serial_clk),
    .D(_00746_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[81] ));
 sky130_fd_sc_hd__dfrtp_2 _26949_ (.CLK(A_in_serial_clk),
    .D(_00747_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[82] ));
 sky130_fd_sc_hd__dfrtp_2 _26950_ (.CLK(A_in_serial_clk),
    .D(_00748_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[83] ));
 sky130_fd_sc_hd__dfrtp_2 _26951_ (.CLK(A_in_serial_clk),
    .D(_00749_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[84] ));
 sky130_fd_sc_hd__dfrtp_2 _26952_ (.CLK(A_in_serial_clk),
    .D(_00750_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[85] ));
 sky130_fd_sc_hd__dfrtp_2 _26953_ (.CLK(A_in_serial_clk),
    .D(_00751_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[86] ));
 sky130_fd_sc_hd__dfrtp_2 _26954_ (.CLK(A_in_serial_clk),
    .D(_00752_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[87] ));
 sky130_fd_sc_hd__dfrtp_2 _26955_ (.CLK(A_in_serial_clk),
    .D(_00753_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[88] ));
 sky130_fd_sc_hd__dfrtp_2 _26956_ (.CLK(A_in_serial_clk),
    .D(_00754_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[89] ));
 sky130_fd_sc_hd__dfrtp_2 _26957_ (.CLK(A_in_serial_clk),
    .D(_00755_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[90] ));
 sky130_fd_sc_hd__dfrtp_2 _26958_ (.CLK(A_in_serial_clk),
    .D(_00756_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[91] ));
 sky130_fd_sc_hd__dfrtp_2 _26959_ (.CLK(A_in_serial_clk),
    .D(_00757_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[92] ));
 sky130_fd_sc_hd__dfrtp_2 _26960_ (.CLK(A_in_serial_clk),
    .D(_00758_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[93] ));
 sky130_fd_sc_hd__dfrtp_2 _26961_ (.CLK(A_in_serial_clk),
    .D(_00759_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[94] ));
 sky130_fd_sc_hd__dfrtp_2 _26962_ (.CLK(A_in_serial_clk),
    .D(_00760_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[95] ));
 sky130_fd_sc_hd__dfrtp_2 _26963_ (.CLK(A_in_serial_clk),
    .D(_00761_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[96] ));
 sky130_fd_sc_hd__dfrtp_2 _26964_ (.CLK(A_in_serial_clk),
    .D(_00762_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[97] ));
 sky130_fd_sc_hd__dfrtp_2 _26965_ (.CLK(A_in_serial_clk),
    .D(_00763_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[98] ));
 sky130_fd_sc_hd__dfrtp_2 _26966_ (.CLK(A_in_serial_clk),
    .D(_00764_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[99] ));
 sky130_fd_sc_hd__dfrtp_2 _26967_ (.CLK(A_in_serial_clk),
    .D(_00765_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[100] ));
 sky130_fd_sc_hd__dfrtp_2 _26968_ (.CLK(A_in_serial_clk),
    .D(_00766_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[101] ));
 sky130_fd_sc_hd__dfrtp_2 _26969_ (.CLK(A_in_serial_clk),
    .D(_00767_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[102] ));
 sky130_fd_sc_hd__dfrtp_2 _26970_ (.CLK(A_in_serial_clk),
    .D(_00768_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[103] ));
 sky130_fd_sc_hd__dfrtp_2 _26971_ (.CLK(A_in_serial_clk),
    .D(_00769_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[104] ));
 sky130_fd_sc_hd__dfrtp_2 _26972_ (.CLK(A_in_serial_clk),
    .D(_00770_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[105] ));
 sky130_fd_sc_hd__dfrtp_2 _26973_ (.CLK(A_in_serial_clk),
    .D(_00771_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[106] ));
 sky130_fd_sc_hd__dfrtp_2 _26974_ (.CLK(A_in_serial_clk),
    .D(_00772_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[107] ));
 sky130_fd_sc_hd__dfrtp_2 _26975_ (.CLK(A_in_serial_clk),
    .D(_00773_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[108] ));
 sky130_fd_sc_hd__dfrtp_2 _26976_ (.CLK(A_in_serial_clk),
    .D(_00774_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[109] ));
 sky130_fd_sc_hd__dfrtp_2 _26977_ (.CLK(A_in_serial_clk),
    .D(_00775_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[110] ));
 sky130_fd_sc_hd__dfrtp_2 _26978_ (.CLK(A_in_serial_clk),
    .D(_00776_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[111] ));
 sky130_fd_sc_hd__dfrtp_2 _26979_ (.CLK(A_in_serial_clk),
    .D(_00777_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[112] ));
 sky130_fd_sc_hd__dfrtp_2 _26980_ (.CLK(A_in_serial_clk),
    .D(_00778_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[113] ));
 sky130_fd_sc_hd__dfrtp_2 _26981_ (.CLK(A_in_serial_clk),
    .D(_00779_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[114] ));
 sky130_fd_sc_hd__dfrtp_2 _26982_ (.CLK(A_in_serial_clk),
    .D(_00780_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[115] ));
 sky130_fd_sc_hd__dfrtp_2 _26983_ (.CLK(A_in_serial_clk),
    .D(_00781_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[116] ));
 sky130_fd_sc_hd__dfrtp_2 _26984_ (.CLK(A_in_serial_clk),
    .D(_00782_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[117] ));
 sky130_fd_sc_hd__dfrtp_2 _26985_ (.CLK(A_in_serial_clk),
    .D(_00783_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[118] ));
 sky130_fd_sc_hd__dfrtp_2 _26986_ (.CLK(A_in_serial_clk),
    .D(_00784_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[119] ));
 sky130_fd_sc_hd__dfrtp_2 _26987_ (.CLK(A_in_serial_clk),
    .D(_00785_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[120] ));
 sky130_fd_sc_hd__dfrtp_2 _26988_ (.CLK(A_in_serial_clk),
    .D(_00786_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[121] ));
 sky130_fd_sc_hd__dfrtp_2 _26989_ (.CLK(A_in_serial_clk),
    .D(_00787_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[122] ));
 sky130_fd_sc_hd__dfrtp_2 _26990_ (.CLK(A_in_serial_clk),
    .D(_00788_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[123] ));
 sky130_fd_sc_hd__dfrtp_2 _26991_ (.CLK(A_in_serial_clk),
    .D(_00789_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[124] ));
 sky130_fd_sc_hd__dfrtp_2 _26992_ (.CLK(A_in_serial_clk),
    .D(_00790_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[125] ));
 sky130_fd_sc_hd__dfrtp_2 _26993_ (.CLK(A_in_serial_clk),
    .D(_00791_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[126] ));
 sky130_fd_sc_hd__dfrtp_2 _26994_ (.CLK(A_in_serial_clk),
    .D(_00792_),
    .RESET_B(rst_n),
    .Q(\deser_A.serial_word[127] ));
 sky130_fd_sc_hd__dfrtp_2 _26995_ (.CLK(B_in_serial_clk),
    .D(_00793_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26996_ (.CLK(B_in_serial_clk),
    .D(_00794_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26997_ (.CLK(B_in_serial_clk),
    .D(_00795_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26998_ (.CLK(B_in_serial_clk),
    .D(_00796_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26999_ (.CLK(B_in_serial_clk),
    .D(_00797_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27000_ (.CLK(B_in_serial_clk),
    .D(_00798_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27001_ (.CLK(B_in_serial_clk),
    .D(_00799_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27002_ (.CLK(B_in_serial_clk),
    .D(_00800_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27003_ (.CLK(B_in_serial_clk),
    .D(_00801_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27004_ (.CLK(B_in_serial_clk),
    .D(_00802_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27005_ (.CLK(B_in_serial_clk),
    .D(_00803_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27006_ (.CLK(B_in_serial_clk),
    .D(_00804_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27007_ (.CLK(B_in_serial_clk),
    .D(_00805_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27008_ (.CLK(B_in_serial_clk),
    .D(_00806_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27009_ (.CLK(B_in_serial_clk),
    .D(_00807_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27010_ (.CLK(B_in_serial_clk),
    .D(_00808_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[16] ));
 sky130_fd_sc_hd__dfrtp_2 _27011_ (.CLK(B_in_serial_clk),
    .D(_00809_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[17] ));
 sky130_fd_sc_hd__dfrtp_2 _27012_ (.CLK(B_in_serial_clk),
    .D(_00810_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[18] ));
 sky130_fd_sc_hd__dfrtp_2 _27013_ (.CLK(B_in_serial_clk),
    .D(_00811_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[19] ));
 sky130_fd_sc_hd__dfrtp_2 _27014_ (.CLK(B_in_serial_clk),
    .D(_00812_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[20] ));
 sky130_fd_sc_hd__dfrtp_2 _27015_ (.CLK(B_in_serial_clk),
    .D(_00813_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[21] ));
 sky130_fd_sc_hd__dfrtp_2 _27016_ (.CLK(B_in_serial_clk),
    .D(_00814_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[22] ));
 sky130_fd_sc_hd__dfrtp_2 _27017_ (.CLK(B_in_serial_clk),
    .D(_00815_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[23] ));
 sky130_fd_sc_hd__dfrtp_2 _27018_ (.CLK(B_in_serial_clk),
    .D(_00816_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[24] ));
 sky130_fd_sc_hd__dfrtp_2 _27019_ (.CLK(B_in_serial_clk),
    .D(_00817_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[25] ));
 sky130_fd_sc_hd__dfrtp_2 _27020_ (.CLK(B_in_serial_clk),
    .D(_00818_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[26] ));
 sky130_fd_sc_hd__dfrtp_2 _27021_ (.CLK(B_in_serial_clk),
    .D(_00819_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[27] ));
 sky130_fd_sc_hd__dfrtp_2 _27022_ (.CLK(B_in_serial_clk),
    .D(_00820_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[28] ));
 sky130_fd_sc_hd__dfrtp_2 _27023_ (.CLK(B_in_serial_clk),
    .D(_00821_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[29] ));
 sky130_fd_sc_hd__dfrtp_2 _27024_ (.CLK(B_in_serial_clk),
    .D(_00822_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[30] ));
 sky130_fd_sc_hd__dfrtp_2 _27025_ (.CLK(B_in_serial_clk),
    .D(_00823_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[31] ));
 sky130_fd_sc_hd__dfrtp_2 _27026_ (.CLK(B_in_serial_clk),
    .D(_00824_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[32] ));
 sky130_fd_sc_hd__dfrtp_2 _27027_ (.CLK(B_in_serial_clk),
    .D(_00825_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[33] ));
 sky130_fd_sc_hd__dfrtp_2 _27028_ (.CLK(B_in_serial_clk),
    .D(_00826_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[34] ));
 sky130_fd_sc_hd__dfrtp_2 _27029_ (.CLK(B_in_serial_clk),
    .D(_00827_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[35] ));
 sky130_fd_sc_hd__dfrtp_2 _27030_ (.CLK(B_in_serial_clk),
    .D(_00828_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[36] ));
 sky130_fd_sc_hd__dfrtp_2 _27031_ (.CLK(B_in_serial_clk),
    .D(_00829_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[37] ));
 sky130_fd_sc_hd__dfrtp_2 _27032_ (.CLK(B_in_serial_clk),
    .D(_00830_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[38] ));
 sky130_fd_sc_hd__dfrtp_2 _27033_ (.CLK(B_in_serial_clk),
    .D(_00831_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[39] ));
 sky130_fd_sc_hd__dfrtp_2 _27034_ (.CLK(B_in_serial_clk),
    .D(_00832_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[40] ));
 sky130_fd_sc_hd__dfrtp_2 _27035_ (.CLK(B_in_serial_clk),
    .D(_00833_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[41] ));
 sky130_fd_sc_hd__dfrtp_2 _27036_ (.CLK(B_in_serial_clk),
    .D(_00834_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[42] ));
 sky130_fd_sc_hd__dfrtp_2 _27037_ (.CLK(B_in_serial_clk),
    .D(_00835_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[43] ));
 sky130_fd_sc_hd__dfrtp_2 _27038_ (.CLK(B_in_serial_clk),
    .D(_00836_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[44] ));
 sky130_fd_sc_hd__dfrtp_2 _27039_ (.CLK(B_in_serial_clk),
    .D(_00837_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[45] ));
 sky130_fd_sc_hd__dfrtp_2 _27040_ (.CLK(B_in_serial_clk),
    .D(_00838_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[46] ));
 sky130_fd_sc_hd__dfrtp_2 _27041_ (.CLK(B_in_serial_clk),
    .D(_00839_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[47] ));
 sky130_fd_sc_hd__dfrtp_2 _27042_ (.CLK(B_in_serial_clk),
    .D(_00840_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[48] ));
 sky130_fd_sc_hd__dfrtp_2 _27043_ (.CLK(B_in_serial_clk),
    .D(_00841_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[49] ));
 sky130_fd_sc_hd__dfrtp_2 _27044_ (.CLK(B_in_serial_clk),
    .D(_00842_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[50] ));
 sky130_fd_sc_hd__dfrtp_2 _27045_ (.CLK(B_in_serial_clk),
    .D(_00843_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[51] ));
 sky130_fd_sc_hd__dfrtp_2 _27046_ (.CLK(B_in_serial_clk),
    .D(_00844_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[52] ));
 sky130_fd_sc_hd__dfrtp_2 _27047_ (.CLK(B_in_serial_clk),
    .D(_00845_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[53] ));
 sky130_fd_sc_hd__dfrtp_2 _27048_ (.CLK(B_in_serial_clk),
    .D(_00846_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[54] ));
 sky130_fd_sc_hd__dfrtp_2 _27049_ (.CLK(B_in_serial_clk),
    .D(_00847_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[55] ));
 sky130_fd_sc_hd__dfrtp_2 _27050_ (.CLK(B_in_serial_clk),
    .D(_00848_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[56] ));
 sky130_fd_sc_hd__dfrtp_2 _27051_ (.CLK(B_in_serial_clk),
    .D(_00849_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[57] ));
 sky130_fd_sc_hd__dfrtp_2 _27052_ (.CLK(B_in_serial_clk),
    .D(_00850_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[58] ));
 sky130_fd_sc_hd__dfrtp_2 _27053_ (.CLK(B_in_serial_clk),
    .D(_00851_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[59] ));
 sky130_fd_sc_hd__dfrtp_2 _27054_ (.CLK(B_in_serial_clk),
    .D(_00852_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[60] ));
 sky130_fd_sc_hd__dfrtp_2 _27055_ (.CLK(B_in_serial_clk),
    .D(_00853_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[61] ));
 sky130_fd_sc_hd__dfrtp_2 _27056_ (.CLK(B_in_serial_clk),
    .D(_00854_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[62] ));
 sky130_fd_sc_hd__dfrtp_2 _27057_ (.CLK(B_in_serial_clk),
    .D(_00855_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[63] ));
 sky130_fd_sc_hd__dfrtp_2 _27058_ (.CLK(B_in_serial_clk),
    .D(_00856_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[64] ));
 sky130_fd_sc_hd__dfrtp_2 _27059_ (.CLK(B_in_serial_clk),
    .D(_00857_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[65] ));
 sky130_fd_sc_hd__dfrtp_2 _27060_ (.CLK(B_in_serial_clk),
    .D(_00858_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[66] ));
 sky130_fd_sc_hd__dfrtp_2 _27061_ (.CLK(B_in_serial_clk),
    .D(_00859_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[67] ));
 sky130_fd_sc_hd__dfrtp_2 _27062_ (.CLK(B_in_serial_clk),
    .D(_00860_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[68] ));
 sky130_fd_sc_hd__dfrtp_2 _27063_ (.CLK(B_in_serial_clk),
    .D(_00861_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[69] ));
 sky130_fd_sc_hd__dfrtp_2 _27064_ (.CLK(B_in_serial_clk),
    .D(_00862_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[70] ));
 sky130_fd_sc_hd__dfrtp_2 _27065_ (.CLK(B_in_serial_clk),
    .D(_00863_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[71] ));
 sky130_fd_sc_hd__dfrtp_2 _27066_ (.CLK(B_in_serial_clk),
    .D(_00864_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[72] ));
 sky130_fd_sc_hd__dfrtp_2 _27067_ (.CLK(B_in_serial_clk),
    .D(_00865_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[73] ));
 sky130_fd_sc_hd__dfrtp_2 _27068_ (.CLK(B_in_serial_clk),
    .D(_00866_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[74] ));
 sky130_fd_sc_hd__dfrtp_2 _27069_ (.CLK(B_in_serial_clk),
    .D(_00867_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[75] ));
 sky130_fd_sc_hd__dfrtp_2 _27070_ (.CLK(B_in_serial_clk),
    .D(_00868_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[76] ));
 sky130_fd_sc_hd__dfrtp_2 _27071_ (.CLK(B_in_serial_clk),
    .D(_00869_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[77] ));
 sky130_fd_sc_hd__dfrtp_2 _27072_ (.CLK(B_in_serial_clk),
    .D(_00870_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[78] ));
 sky130_fd_sc_hd__dfrtp_2 _27073_ (.CLK(B_in_serial_clk),
    .D(_00871_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[79] ));
 sky130_fd_sc_hd__dfrtp_2 _27074_ (.CLK(B_in_serial_clk),
    .D(_00872_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[80] ));
 sky130_fd_sc_hd__dfrtp_2 _27075_ (.CLK(B_in_serial_clk),
    .D(_00873_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[81] ));
 sky130_fd_sc_hd__dfrtp_2 _27076_ (.CLK(B_in_serial_clk),
    .D(_00874_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[82] ));
 sky130_fd_sc_hd__dfrtp_2 _27077_ (.CLK(B_in_serial_clk),
    .D(_00875_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[83] ));
 sky130_fd_sc_hd__dfrtp_2 _27078_ (.CLK(B_in_serial_clk),
    .D(_00876_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[84] ));
 sky130_fd_sc_hd__dfrtp_2 _27079_ (.CLK(B_in_serial_clk),
    .D(_00877_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[85] ));
 sky130_fd_sc_hd__dfrtp_2 _27080_ (.CLK(B_in_serial_clk),
    .D(_00878_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[86] ));
 sky130_fd_sc_hd__dfrtp_2 _27081_ (.CLK(B_in_serial_clk),
    .D(_00879_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[87] ));
 sky130_fd_sc_hd__dfrtp_2 _27082_ (.CLK(B_in_serial_clk),
    .D(_00880_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[88] ));
 sky130_fd_sc_hd__dfrtp_2 _27083_ (.CLK(B_in_serial_clk),
    .D(_00881_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[89] ));
 sky130_fd_sc_hd__dfrtp_2 _27084_ (.CLK(B_in_serial_clk),
    .D(_00882_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[90] ));
 sky130_fd_sc_hd__dfrtp_2 _27085_ (.CLK(B_in_serial_clk),
    .D(_00883_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[91] ));
 sky130_fd_sc_hd__dfrtp_2 _27086_ (.CLK(B_in_serial_clk),
    .D(_00884_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[92] ));
 sky130_fd_sc_hd__dfrtp_2 _27087_ (.CLK(B_in_serial_clk),
    .D(_00885_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[93] ));
 sky130_fd_sc_hd__dfrtp_2 _27088_ (.CLK(B_in_serial_clk),
    .D(_00886_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[94] ));
 sky130_fd_sc_hd__dfrtp_2 _27089_ (.CLK(B_in_serial_clk),
    .D(_00887_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[95] ));
 sky130_fd_sc_hd__dfrtp_2 _27090_ (.CLK(B_in_serial_clk),
    .D(_00888_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[96] ));
 sky130_fd_sc_hd__dfrtp_2 _27091_ (.CLK(B_in_serial_clk),
    .D(_00889_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[97] ));
 sky130_fd_sc_hd__dfrtp_2 _27092_ (.CLK(B_in_serial_clk),
    .D(_00890_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[98] ));
 sky130_fd_sc_hd__dfrtp_2 _27093_ (.CLK(B_in_serial_clk),
    .D(_00891_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[99] ));
 sky130_fd_sc_hd__dfrtp_2 _27094_ (.CLK(B_in_serial_clk),
    .D(_00892_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[100] ));
 sky130_fd_sc_hd__dfrtp_2 _27095_ (.CLK(B_in_serial_clk),
    .D(_00893_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[101] ));
 sky130_fd_sc_hd__dfrtp_2 _27096_ (.CLK(B_in_serial_clk),
    .D(_00894_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[102] ));
 sky130_fd_sc_hd__dfrtp_2 _27097_ (.CLK(B_in_serial_clk),
    .D(_00895_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[103] ));
 sky130_fd_sc_hd__dfrtp_2 _27098_ (.CLK(B_in_serial_clk),
    .D(_00896_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[104] ));
 sky130_fd_sc_hd__dfrtp_2 _27099_ (.CLK(B_in_serial_clk),
    .D(_00897_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[105] ));
 sky130_fd_sc_hd__dfrtp_2 _27100_ (.CLK(B_in_serial_clk),
    .D(_00898_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[106] ));
 sky130_fd_sc_hd__dfrtp_2 _27101_ (.CLK(B_in_serial_clk),
    .D(_00899_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[107] ));
 sky130_fd_sc_hd__dfrtp_2 _27102_ (.CLK(B_in_serial_clk),
    .D(_00900_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[108] ));
 sky130_fd_sc_hd__dfrtp_2 _27103_ (.CLK(B_in_serial_clk),
    .D(_00901_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[109] ));
 sky130_fd_sc_hd__dfrtp_2 _27104_ (.CLK(B_in_serial_clk),
    .D(_00902_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[110] ));
 sky130_fd_sc_hd__dfrtp_2 _27105_ (.CLK(B_in_serial_clk),
    .D(_00903_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[111] ));
 sky130_fd_sc_hd__dfrtp_2 _27106_ (.CLK(B_in_serial_clk),
    .D(_00904_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[112] ));
 sky130_fd_sc_hd__dfrtp_2 _27107_ (.CLK(B_in_serial_clk),
    .D(_00905_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[113] ));
 sky130_fd_sc_hd__dfrtp_2 _27108_ (.CLK(B_in_serial_clk),
    .D(_00906_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[114] ));
 sky130_fd_sc_hd__dfrtp_2 _27109_ (.CLK(B_in_serial_clk),
    .D(_00907_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[115] ));
 sky130_fd_sc_hd__dfrtp_2 _27110_ (.CLK(B_in_serial_clk),
    .D(_00908_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[116] ));
 sky130_fd_sc_hd__dfrtp_2 _27111_ (.CLK(B_in_serial_clk),
    .D(_00909_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[117] ));
 sky130_fd_sc_hd__dfrtp_2 _27112_ (.CLK(B_in_serial_clk),
    .D(_00910_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[118] ));
 sky130_fd_sc_hd__dfrtp_2 _27113_ (.CLK(B_in_serial_clk),
    .D(_00911_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[119] ));
 sky130_fd_sc_hd__dfrtp_2 _27114_ (.CLK(B_in_serial_clk),
    .D(_00912_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[120] ));
 sky130_fd_sc_hd__dfrtp_2 _27115_ (.CLK(B_in_serial_clk),
    .D(_00913_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[121] ));
 sky130_fd_sc_hd__dfrtp_2 _27116_ (.CLK(B_in_serial_clk),
    .D(_00914_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[122] ));
 sky130_fd_sc_hd__dfrtp_2 _27117_ (.CLK(B_in_serial_clk),
    .D(_00915_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[123] ));
 sky130_fd_sc_hd__dfrtp_2 _27118_ (.CLK(B_in_serial_clk),
    .D(_00916_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[124] ));
 sky130_fd_sc_hd__dfrtp_2 _27119_ (.CLK(B_in_serial_clk),
    .D(_00917_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[125] ));
 sky130_fd_sc_hd__dfrtp_2 _27120_ (.CLK(B_in_serial_clk),
    .D(_00918_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[126] ));
 sky130_fd_sc_hd__dfrtp_2 _27121_ (.CLK(B_in_serial_clk),
    .D(_00919_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[127] ));
 sky130_fd_sc_hd__dfrtp_2 _27122_ (.CLK(A_in_serial_clk),
    .D(_00920_),
    .RESET_B(rst_n),
    .Q(\deser_A.shift_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27123_ (.CLK(B_in_serial_clk),
    .D(_00921_),
    .RESET_B(rst_n),
    .Q(\deser_B.shift_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27124_ (.CLK(clk),
    .D(_00922_),
    .Q(\systolic_inst.A_shift[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27125_ (.CLK(clk),
    .D(_00923_),
    .Q(\systolic_inst.A_shift[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27126_ (.CLK(clk),
    .D(_00924_),
    .Q(\systolic_inst.A_shift[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27127_ (.CLK(clk),
    .D(_00925_),
    .Q(\systolic_inst.A_shift[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27128_ (.CLK(clk),
    .D(_00926_),
    .Q(\systolic_inst.A_shift[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27129_ (.CLK(clk),
    .D(_00927_),
    .Q(\systolic_inst.A_shift[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27130_ (.CLK(clk),
    .D(_00928_),
    .Q(\systolic_inst.A_shift[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27131_ (.CLK(clk),
    .D(_00929_),
    .Q(\systolic_inst.A_shift[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27132_ (.CLK(clk),
    .D(_00930_),
    .Q(\systolic_inst.B_shift[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27133_ (.CLK(clk),
    .D(_00931_),
    .Q(\systolic_inst.B_shift[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27134_ (.CLK(clk),
    .D(_00932_),
    .Q(\systolic_inst.B_shift[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27135_ (.CLK(clk),
    .D(_00933_),
    .Q(\systolic_inst.B_shift[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27136_ (.CLK(clk),
    .D(_00934_),
    .Q(\systolic_inst.B_shift[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27137_ (.CLK(clk),
    .D(_00935_),
    .Q(\systolic_inst.B_shift[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27138_ (.CLK(clk),
    .D(_00936_),
    .Q(\systolic_inst.B_shift[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27139_ (.CLK(clk),
    .D(_00937_),
    .Q(\systolic_inst.B_shift[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27140_ (.CLK(clk),
    .D(_00938_),
    .Q(\systolic_inst.A_shift[21][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27141_ (.CLK(clk),
    .D(_00939_),
    .Q(\systolic_inst.A_shift[21][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27142_ (.CLK(clk),
    .D(_00940_),
    .Q(\systolic_inst.A_shift[21][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27143_ (.CLK(clk),
    .D(_00941_),
    .Q(\systolic_inst.A_shift[21][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27144_ (.CLK(clk),
    .D(_00942_),
    .Q(\systolic_inst.A_shift[21][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27145_ (.CLK(clk),
    .D(_00943_),
    .Q(\systolic_inst.A_shift[21][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27146_ (.CLK(clk),
    .D(_00944_),
    .Q(\systolic_inst.A_shift[21][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27147_ (.CLK(clk),
    .D(_00945_),
    .Q(\systolic_inst.A_shift[21][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27148_ (.CLK(clk),
    .D(_00946_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[15][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27149_ (.CLK(clk),
    .D(_00947_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[15][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27150_ (.CLK(clk),
    .D(_00948_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[15][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27151_ (.CLK(clk),
    .D(_00949_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[15][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27152_ (.CLK(clk),
    .D(_00950_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[15][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27153_ (.CLK(clk),
    .D(_00951_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[15][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27154_ (.CLK(clk),
    .D(_00952_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[15][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27155_ (.CLK(clk),
    .D(_00953_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[15][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27156_ (.CLK(clk),
    .D(_00954_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[14][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27157_ (.CLK(clk),
    .D(_00955_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[14][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27158_ (.CLK(clk),
    .D(_00956_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[14][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27159_ (.CLK(clk),
    .D(_00957_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[14][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27160_ (.CLK(clk),
    .D(_00958_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[14][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27161_ (.CLK(clk),
    .D(_00959_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[14][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27162_ (.CLK(clk),
    .D(_00960_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[14][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27163_ (.CLK(clk),
    .D(_00961_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[14][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27164_ (.CLK(clk),
    .D(_00962_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27165_ (.CLK(clk),
    .D(_00963_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27166_ (.CLK(clk),
    .D(_00964_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27167_ (.CLK(clk),
    .D(_00965_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27168_ (.CLK(clk),
    .D(_00966_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27169_ (.CLK(clk),
    .D(_00967_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27170_ (.CLK(clk),
    .D(_00968_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27171_ (.CLK(clk),
    .D(_00969_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27172_ (.CLK(clk),
    .D(_00970_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27173_ (.CLK(clk),
    .D(_00971_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27174_ (.CLK(clk),
    .D(_00972_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27175_ (.CLK(clk),
    .D(_00973_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27176_ (.CLK(clk),
    .D(_00974_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27177_ (.CLK(clk),
    .D(_00975_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27178_ (.CLK(clk),
    .D(_00976_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27179_ (.CLK(clk),
    .D(_00977_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[3].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27180_ (.CLK(clk),
    .D(_00978_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27181_ (.CLK(clk),
    .D(_00979_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27182_ (.CLK(clk),
    .D(_00980_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27183_ (.CLK(clk),
    .D(_00981_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27184_ (.CLK(clk),
    .D(_00982_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27185_ (.CLK(clk),
    .D(_00983_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27186_ (.CLK(clk),
    .D(_00984_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27187_ (.CLK(clk),
    .D(_00985_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27188_ (.CLK(clk),
    .D(_00986_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27189_ (.CLK(clk),
    .D(_00987_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27190_ (.CLK(clk),
    .D(_00988_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27191_ (.CLK(clk),
    .D(_00989_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27192_ (.CLK(clk),
    .D(_00990_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27193_ (.CLK(clk),
    .D(_00991_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27194_ (.CLK(clk),
    .D(_00992_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27195_ (.CLK(clk),
    .D(_00993_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27196_ (.CLK(clk),
    .D(_00994_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27197_ (.CLK(clk),
    .D(_00995_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27198_ (.CLK(clk),
    .D(_00996_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27199_ (.CLK(clk),
    .D(_00997_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27200_ (.CLK(clk),
    .D(_00998_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27201_ (.CLK(clk),
    .D(_00999_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27202_ (.CLK(clk),
    .D(_01000_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27203_ (.CLK(clk),
    .D(_01001_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27204_ (.CLK(clk),
    .D(_01002_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27205_ (.CLK(clk),
    .D(_01003_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27206_ (.CLK(clk),
    .D(_01004_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27207_ (.CLK(clk),
    .D(_01005_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27208_ (.CLK(clk),
    .D(_01006_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27209_ (.CLK(clk),
    .D(_01007_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27210_ (.CLK(clk),
    .D(_01008_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27211_ (.CLK(clk),
    .D(_01009_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[15][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27212_ (.CLK(clk),
    .D(_01010_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[14][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27213_ (.CLK(clk),
    .D(_01011_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[14][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27214_ (.CLK(clk),
    .D(_01012_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[14][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27215_ (.CLK(clk),
    .D(_01013_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[14][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27216_ (.CLK(clk),
    .D(_01014_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[14][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27217_ (.CLK(clk),
    .D(_01015_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[14][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27218_ (.CLK(clk),
    .D(_01016_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[14][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27219_ (.CLK(clk),
    .D(_01017_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[14][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27220_ (.CLK(clk),
    .D(_01018_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[13][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27221_ (.CLK(clk),
    .D(_01019_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[13][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27222_ (.CLK(clk),
    .D(_01020_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[13][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27223_ (.CLK(clk),
    .D(_01021_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[13][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27224_ (.CLK(clk),
    .D(_01022_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[13][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27225_ (.CLK(clk),
    .D(_01023_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[13][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27226_ (.CLK(clk),
    .D(_01024_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[13][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27227_ (.CLK(clk),
    .D(_01025_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[13][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27228_ (.CLK(clk),
    .D(_01026_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27229_ (.CLK(clk),
    .D(_01027_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27230_ (.CLK(clk),
    .D(_01028_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27231_ (.CLK(clk),
    .D(_01029_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27232_ (.CLK(clk),
    .D(_01030_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27233_ (.CLK(clk),
    .D(_01031_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27234_ (.CLK(clk),
    .D(_01032_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27235_ (.CLK(clk),
    .D(_01033_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27236_ (.CLK(clk),
    .D(_01034_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27237_ (.CLK(clk),
    .D(_01035_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27238_ (.CLK(clk),
    .D(_01036_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27239_ (.CLK(clk),
    .D(_01037_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27240_ (.CLK(clk),
    .D(_01038_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27241_ (.CLK(clk),
    .D(_01039_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27242_ (.CLK(clk),
    .D(_01040_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27243_ (.CLK(clk),
    .D(_01041_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[2].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27244_ (.CLK(clk),
    .D(_01042_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27245_ (.CLK(clk),
    .D(_01043_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27246_ (.CLK(clk),
    .D(_01044_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27247_ (.CLK(clk),
    .D(_01045_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27248_ (.CLK(clk),
    .D(_01046_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27249_ (.CLK(clk),
    .D(_01047_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27250_ (.CLK(clk),
    .D(_01048_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27251_ (.CLK(clk),
    .D(_01049_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27252_ (.CLK(clk),
    .D(_01050_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27253_ (.CLK(clk),
    .D(_01051_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27254_ (.CLK(clk),
    .D(_01052_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27255_ (.CLK(clk),
    .D(_01053_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27256_ (.CLK(clk),
    .D(_01054_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27257_ (.CLK(clk),
    .D(_01055_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27258_ (.CLK(clk),
    .D(_01056_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27259_ (.CLK(clk),
    .D(_01057_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27260_ (.CLK(clk),
    .D(_01058_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27261_ (.CLK(clk),
    .D(_01059_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27262_ (.CLK(clk),
    .D(_01060_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27263_ (.CLK(clk),
    .D(_01061_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27264_ (.CLK(clk),
    .D(_01062_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27265_ (.CLK(clk),
    .D(_01063_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27266_ (.CLK(clk),
    .D(_01064_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27267_ (.CLK(clk),
    .D(_01065_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27268_ (.CLK(clk),
    .D(_01066_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27269_ (.CLK(clk),
    .D(_01067_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27270_ (.CLK(clk),
    .D(_01068_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27271_ (.CLK(clk),
    .D(_01069_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27272_ (.CLK(clk),
    .D(_01070_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27273_ (.CLK(clk),
    .D(_01071_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27274_ (.CLK(clk),
    .D(_01072_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27275_ (.CLK(clk),
    .D(_01073_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[14][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27276_ (.CLK(clk),
    .D(_01074_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[13][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27277_ (.CLK(clk),
    .D(_01075_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[13][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27278_ (.CLK(clk),
    .D(_01076_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[13][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27279_ (.CLK(clk),
    .D(_01077_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[13][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27280_ (.CLK(clk),
    .D(_01078_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[13][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27281_ (.CLK(clk),
    .D(_01079_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[13][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27282_ (.CLK(clk),
    .D(_01080_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[13][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27283_ (.CLK(clk),
    .D(_01081_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[13][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27284_ (.CLK(clk),
    .D(_01082_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[12][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27285_ (.CLK(clk),
    .D(_01083_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[12][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27286_ (.CLK(clk),
    .D(_01084_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[12][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27287_ (.CLK(clk),
    .D(_01085_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[12][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27288_ (.CLK(clk),
    .D(_01086_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[12][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27289_ (.CLK(clk),
    .D(_01087_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[12][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27290_ (.CLK(clk),
    .D(_01088_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[12][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27291_ (.CLK(clk),
    .D(_01089_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[12][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27292_ (.CLK(clk),
    .D(_01090_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27293_ (.CLK(clk),
    .D(_01091_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27294_ (.CLK(clk),
    .D(_01092_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27295_ (.CLK(clk),
    .D(_01093_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27296_ (.CLK(clk),
    .D(_01094_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27297_ (.CLK(clk),
    .D(_01095_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27298_ (.CLK(clk),
    .D(_01096_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27299_ (.CLK(clk),
    .D(_01097_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27300_ (.CLK(clk),
    .D(_01098_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27301_ (.CLK(clk),
    .D(_01099_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27302_ (.CLK(clk),
    .D(_01100_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27303_ (.CLK(clk),
    .D(_01101_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27304_ (.CLK(clk),
    .D(_01102_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27305_ (.CLK(clk),
    .D(_01103_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27306_ (.CLK(clk),
    .D(_01104_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27307_ (.CLK(clk),
    .D(_01105_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[1].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27308_ (.CLK(clk),
    .D(_01106_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27309_ (.CLK(clk),
    .D(_01107_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27310_ (.CLK(clk),
    .D(_01108_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27311_ (.CLK(clk),
    .D(_01109_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27312_ (.CLK(clk),
    .D(_01110_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27313_ (.CLK(clk),
    .D(_01111_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27314_ (.CLK(clk),
    .D(_01112_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27315_ (.CLK(clk),
    .D(_01113_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27316_ (.CLK(clk),
    .D(_01114_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27317_ (.CLK(clk),
    .D(_01115_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27318_ (.CLK(clk),
    .D(_01116_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27319_ (.CLK(clk),
    .D(_01117_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27320_ (.CLK(clk),
    .D(_01118_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27321_ (.CLK(clk),
    .D(_01119_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27322_ (.CLK(clk),
    .D(_01120_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27323_ (.CLK(clk),
    .D(_01121_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27324_ (.CLK(clk),
    .D(_01122_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27325_ (.CLK(clk),
    .D(_01123_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27326_ (.CLK(clk),
    .D(_01124_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27327_ (.CLK(clk),
    .D(_01125_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27328_ (.CLK(clk),
    .D(_01126_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27329_ (.CLK(clk),
    .D(_01127_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27330_ (.CLK(clk),
    .D(_01128_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27331_ (.CLK(clk),
    .D(_01129_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27332_ (.CLK(clk),
    .D(_01130_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27333_ (.CLK(clk),
    .D(_01131_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27334_ (.CLK(clk),
    .D(_01132_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27335_ (.CLK(clk),
    .D(_01133_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27336_ (.CLK(clk),
    .D(_01134_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27337_ (.CLK(clk),
    .D(_01135_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27338_ (.CLK(clk),
    .D(_01136_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27339_ (.CLK(clk),
    .D(_01137_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[13][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27340_ (.CLK(clk),
    .D(_01138_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[12][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27341_ (.CLK(clk),
    .D(_01139_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[12][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27342_ (.CLK(clk),
    .D(_01140_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[12][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27343_ (.CLK(clk),
    .D(_01141_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[12][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27344_ (.CLK(clk),
    .D(_01142_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[12][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27345_ (.CLK(clk),
    .D(_01143_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[12][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27346_ (.CLK(clk),
    .D(_01144_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[12][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27347_ (.CLK(clk),
    .D(_01145_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[12][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27348_ (.CLK(clk),
    .D(_01146_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[11][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27349_ (.CLK(clk),
    .D(_01147_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[11][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27350_ (.CLK(clk),
    .D(_01148_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[11][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27351_ (.CLK(clk),
    .D(_01149_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[11][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27352_ (.CLK(clk),
    .D(_01150_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[11][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27353_ (.CLK(clk),
    .D(_01151_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[11][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27354_ (.CLK(clk),
    .D(_01152_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[11][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27355_ (.CLK(clk),
    .D(_01153_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[11][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27356_ (.CLK(clk),
    .D(_01154_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27357_ (.CLK(clk),
    .D(_01155_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27358_ (.CLK(clk),
    .D(_01156_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27359_ (.CLK(clk),
    .D(_01157_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27360_ (.CLK(clk),
    .D(_01158_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27361_ (.CLK(clk),
    .D(_01159_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27362_ (.CLK(clk),
    .D(_01160_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27363_ (.CLK(clk),
    .D(_01161_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27364_ (.CLK(clk),
    .D(_01162_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27365_ (.CLK(clk),
    .D(_01163_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27366_ (.CLK(clk),
    .D(_01164_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27367_ (.CLK(clk),
    .D(_01165_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27368_ (.CLK(clk),
    .D(_01166_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27369_ (.CLK(clk),
    .D(_01167_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27370_ (.CLK(clk),
    .D(_01168_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27371_ (.CLK(clk),
    .D(_01169_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[3].col_loop[0].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27372_ (.CLK(clk),
    .D(_01170_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27373_ (.CLK(clk),
    .D(_01171_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27374_ (.CLK(clk),
    .D(_01172_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27375_ (.CLK(clk),
    .D(_01173_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27376_ (.CLK(clk),
    .D(_01174_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27377_ (.CLK(clk),
    .D(_01175_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27378_ (.CLK(clk),
    .D(_01176_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27379_ (.CLK(clk),
    .D(_01177_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27380_ (.CLK(clk),
    .D(_01178_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27381_ (.CLK(clk),
    .D(_01179_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27382_ (.CLK(clk),
    .D(_01180_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27383_ (.CLK(clk),
    .D(_01181_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27384_ (.CLK(clk),
    .D(_01182_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27385_ (.CLK(clk),
    .D(_01183_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27386_ (.CLK(clk),
    .D(_01184_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27387_ (.CLK(clk),
    .D(_01185_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27388_ (.CLK(clk),
    .D(_01186_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27389_ (.CLK(clk),
    .D(_01187_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27390_ (.CLK(clk),
    .D(_01188_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27391_ (.CLK(clk),
    .D(_01189_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27392_ (.CLK(clk),
    .D(_01190_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27393_ (.CLK(clk),
    .D(_01191_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27394_ (.CLK(clk),
    .D(_01192_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27395_ (.CLK(clk),
    .D(_01193_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27396_ (.CLK(clk),
    .D(_01194_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27397_ (.CLK(clk),
    .D(_01195_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27398_ (.CLK(clk),
    .D(_01196_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27399_ (.CLK(clk),
    .D(_01197_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27400_ (.CLK(clk),
    .D(_01198_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27401_ (.CLK(clk),
    .D(_01199_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27402_ (.CLK(clk),
    .D(_01200_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27403_ (.CLK(clk),
    .D(_01201_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[12][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27404_ (.CLK(clk),
    .D(_01202_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[11][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27405_ (.CLK(clk),
    .D(_01203_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[11][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27406_ (.CLK(clk),
    .D(_01204_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[11][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27407_ (.CLK(clk),
    .D(_01205_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[11][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27408_ (.CLK(clk),
    .D(_01206_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[11][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27409_ (.CLK(clk),
    .D(_01207_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[11][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27410_ (.CLK(clk),
    .D(_01208_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[11][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27411_ (.CLK(clk),
    .D(_01209_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[11][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27412_ (.CLK(clk),
    .D(_01210_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[10][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27413_ (.CLK(clk),
    .D(_01211_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[10][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27414_ (.CLK(clk),
    .D(_01212_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[10][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27415_ (.CLK(clk),
    .D(_01213_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[10][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27416_ (.CLK(clk),
    .D(_01214_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[10][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27417_ (.CLK(clk),
    .D(_01215_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[10][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27418_ (.CLK(clk),
    .D(_01216_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[10][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27419_ (.CLK(clk),
    .D(_01217_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[10][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27420_ (.CLK(clk),
    .D(_01218_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27421_ (.CLK(clk),
    .D(_01219_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27422_ (.CLK(clk),
    .D(_01220_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27423_ (.CLK(clk),
    .D(_01221_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27424_ (.CLK(clk),
    .D(_01222_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27425_ (.CLK(clk),
    .D(_01223_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27426_ (.CLK(clk),
    .D(_01224_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27427_ (.CLK(clk),
    .D(_01225_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27428_ (.CLK(clk),
    .D(_01226_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27429_ (.CLK(clk),
    .D(_01227_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27430_ (.CLK(clk),
    .D(_01228_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27431_ (.CLK(clk),
    .D(_01229_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27432_ (.CLK(clk),
    .D(_01230_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27433_ (.CLK(clk),
    .D(_01231_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27434_ (.CLK(clk),
    .D(_01232_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27435_ (.CLK(clk),
    .D(_01233_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[3].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27436_ (.CLK(clk),
    .D(_01234_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27437_ (.CLK(clk),
    .D(_01235_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27438_ (.CLK(clk),
    .D(_01236_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27439_ (.CLK(clk),
    .D(_01237_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27440_ (.CLK(clk),
    .D(_01238_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27441_ (.CLK(clk),
    .D(_01239_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27442_ (.CLK(clk),
    .D(_01240_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27443_ (.CLK(clk),
    .D(_01241_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27444_ (.CLK(clk),
    .D(_01242_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27445_ (.CLK(clk),
    .D(_01243_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27446_ (.CLK(clk),
    .D(_01244_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27447_ (.CLK(clk),
    .D(_01245_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27448_ (.CLK(clk),
    .D(_01246_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27449_ (.CLK(clk),
    .D(_01247_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27450_ (.CLK(clk),
    .D(_01248_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27451_ (.CLK(clk),
    .D(_01249_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27452_ (.CLK(clk),
    .D(_01250_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27453_ (.CLK(clk),
    .D(_01251_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27454_ (.CLK(clk),
    .D(_01252_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27455_ (.CLK(clk),
    .D(_01253_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27456_ (.CLK(clk),
    .D(_01254_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27457_ (.CLK(clk),
    .D(_01255_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27458_ (.CLK(clk),
    .D(_01256_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27459_ (.CLK(clk),
    .D(_01257_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27460_ (.CLK(clk),
    .D(_01258_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27461_ (.CLK(clk),
    .D(_01259_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27462_ (.CLK(clk),
    .D(_01260_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27463_ (.CLK(clk),
    .D(_01261_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27464_ (.CLK(clk),
    .D(_01262_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27465_ (.CLK(clk),
    .D(_01263_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27466_ (.CLK(clk),
    .D(_01264_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27467_ (.CLK(clk),
    .D(_01265_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[11][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27468_ (.CLK(clk),
    .D(_01266_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[10][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27469_ (.CLK(clk),
    .D(_01267_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[10][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27470_ (.CLK(clk),
    .D(_01268_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[10][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27471_ (.CLK(clk),
    .D(_01269_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[10][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27472_ (.CLK(clk),
    .D(_01270_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[10][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27473_ (.CLK(clk),
    .D(_01271_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[10][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27474_ (.CLK(clk),
    .D(_01272_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[10][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27475_ (.CLK(clk),
    .D(_01273_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[10][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27476_ (.CLK(clk),
    .D(_01274_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[9][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27477_ (.CLK(clk),
    .D(_01275_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[9][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27478_ (.CLK(clk),
    .D(_01276_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[9][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27479_ (.CLK(clk),
    .D(_01277_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[9][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27480_ (.CLK(clk),
    .D(_01278_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[9][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27481_ (.CLK(clk),
    .D(_01279_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[9][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27482_ (.CLK(clk),
    .D(_01280_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[9][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27483_ (.CLK(clk),
    .D(_01281_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[9][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27484_ (.CLK(clk),
    .D(_01282_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27485_ (.CLK(clk),
    .D(_01283_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27486_ (.CLK(clk),
    .D(_01284_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27487_ (.CLK(clk),
    .D(_01285_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27488_ (.CLK(clk),
    .D(_01286_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27489_ (.CLK(clk),
    .D(_01287_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27490_ (.CLK(clk),
    .D(_01288_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27491_ (.CLK(clk),
    .D(_01289_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27492_ (.CLK(clk),
    .D(_01290_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27493_ (.CLK(clk),
    .D(_01291_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27494_ (.CLK(clk),
    .D(_01292_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27495_ (.CLK(clk),
    .D(_01293_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27496_ (.CLK(clk),
    .D(_01294_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27497_ (.CLK(clk),
    .D(_01295_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27498_ (.CLK(clk),
    .D(_01296_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27499_ (.CLK(clk),
    .D(_01297_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[2].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27500_ (.CLK(clk),
    .D(_01298_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27501_ (.CLK(clk),
    .D(_01299_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27502_ (.CLK(clk),
    .D(_01300_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27503_ (.CLK(clk),
    .D(_01301_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27504_ (.CLK(clk),
    .D(_01302_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27505_ (.CLK(clk),
    .D(_01303_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27506_ (.CLK(clk),
    .D(_01304_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27507_ (.CLK(clk),
    .D(_01305_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27508_ (.CLK(clk),
    .D(_01306_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27509_ (.CLK(clk),
    .D(_01307_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27510_ (.CLK(clk),
    .D(_01308_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27511_ (.CLK(clk),
    .D(_01309_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27512_ (.CLK(clk),
    .D(_01310_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27513_ (.CLK(clk),
    .D(_01311_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27514_ (.CLK(clk),
    .D(_01312_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27515_ (.CLK(clk),
    .D(_01313_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27516_ (.CLK(clk),
    .D(_01314_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27517_ (.CLK(clk),
    .D(_01315_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27518_ (.CLK(clk),
    .D(_01316_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27519_ (.CLK(clk),
    .D(_01317_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27520_ (.CLK(clk),
    .D(_01318_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27521_ (.CLK(clk),
    .D(_01319_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27522_ (.CLK(clk),
    .D(_01320_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27523_ (.CLK(clk),
    .D(_01321_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27524_ (.CLK(clk),
    .D(_01322_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27525_ (.CLK(clk),
    .D(_01323_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27526_ (.CLK(clk),
    .D(_01324_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27527_ (.CLK(clk),
    .D(_01325_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27528_ (.CLK(clk),
    .D(_01326_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27529_ (.CLK(clk),
    .D(_01327_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27530_ (.CLK(clk),
    .D(_01328_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27531_ (.CLK(clk),
    .D(_01329_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[10][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27532_ (.CLK(clk),
    .D(_01330_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[9][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27533_ (.CLK(clk),
    .D(_01331_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[9][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27534_ (.CLK(clk),
    .D(_01332_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[9][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27535_ (.CLK(clk),
    .D(_01333_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[9][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27536_ (.CLK(clk),
    .D(_01334_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[9][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27537_ (.CLK(clk),
    .D(_01335_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[9][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27538_ (.CLK(clk),
    .D(_01336_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[9][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27539_ (.CLK(clk),
    .D(_01337_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[9][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27540_ (.CLK(clk),
    .D(_01338_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[8][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27541_ (.CLK(clk),
    .D(_01339_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[8][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27542_ (.CLK(clk),
    .D(_01340_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[8][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27543_ (.CLK(clk),
    .D(_01341_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[8][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27544_ (.CLK(clk),
    .D(_01342_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[8][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27545_ (.CLK(clk),
    .D(_01343_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[8][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27546_ (.CLK(clk),
    .D(_01344_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[8][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27547_ (.CLK(clk),
    .D(_01345_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[8][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27548_ (.CLK(clk),
    .D(_01346_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27549_ (.CLK(clk),
    .D(_01347_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27550_ (.CLK(clk),
    .D(_01348_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27551_ (.CLK(clk),
    .D(_01349_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27552_ (.CLK(clk),
    .D(_01350_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27553_ (.CLK(clk),
    .D(_01351_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27554_ (.CLK(clk),
    .D(_01352_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27555_ (.CLK(clk),
    .D(_01353_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27556_ (.CLK(clk),
    .D(_01354_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27557_ (.CLK(clk),
    .D(_01355_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27558_ (.CLK(clk),
    .D(_01356_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27559_ (.CLK(clk),
    .D(_01357_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27560_ (.CLK(clk),
    .D(_01358_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27561_ (.CLK(clk),
    .D(_01359_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27562_ (.CLK(clk),
    .D(_01360_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27563_ (.CLK(clk),
    .D(_01361_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[1].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27564_ (.CLK(clk),
    .D(_01362_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27565_ (.CLK(clk),
    .D(_01363_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27566_ (.CLK(clk),
    .D(_01364_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27567_ (.CLK(clk),
    .D(_01365_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27568_ (.CLK(clk),
    .D(_01366_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27569_ (.CLK(clk),
    .D(_01367_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27570_ (.CLK(clk),
    .D(_01368_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27571_ (.CLK(clk),
    .D(_01369_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27572_ (.CLK(clk),
    .D(_01370_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27573_ (.CLK(clk),
    .D(_01371_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27574_ (.CLK(clk),
    .D(_01372_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27575_ (.CLK(clk),
    .D(_01373_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27576_ (.CLK(clk),
    .D(_01374_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27577_ (.CLK(clk),
    .D(_01375_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27578_ (.CLK(clk),
    .D(_01376_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27579_ (.CLK(clk),
    .D(_01377_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27580_ (.CLK(clk),
    .D(_01378_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27581_ (.CLK(clk),
    .D(_01379_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27582_ (.CLK(clk),
    .D(_01380_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27583_ (.CLK(clk),
    .D(_01381_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27584_ (.CLK(clk),
    .D(_01382_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27585_ (.CLK(clk),
    .D(_01383_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27586_ (.CLK(clk),
    .D(_01384_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27587_ (.CLK(clk),
    .D(_01385_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27588_ (.CLK(clk),
    .D(_01386_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27589_ (.CLK(clk),
    .D(_01387_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27590_ (.CLK(clk),
    .D(_01388_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27591_ (.CLK(clk),
    .D(_01389_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27592_ (.CLK(clk),
    .D(_01390_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27593_ (.CLK(clk),
    .D(_01391_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27594_ (.CLK(clk),
    .D(_01392_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27595_ (.CLK(clk),
    .D(_01393_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[9][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27596_ (.CLK(clk),
    .D(_01394_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[8][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27597_ (.CLK(clk),
    .D(_01395_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[8][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27598_ (.CLK(clk),
    .D(_01396_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[8][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27599_ (.CLK(clk),
    .D(_01397_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[8][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27600_ (.CLK(clk),
    .D(_01398_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[8][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27601_ (.CLK(clk),
    .D(_01399_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[8][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27602_ (.CLK(clk),
    .D(_01400_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[8][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27603_ (.CLK(clk),
    .D(_01401_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[8][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27604_ (.CLK(clk),
    .D(_01402_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[7][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27605_ (.CLK(clk),
    .D(_01403_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[7][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27606_ (.CLK(clk),
    .D(_01404_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[7][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27607_ (.CLK(clk),
    .D(_01405_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[7][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27608_ (.CLK(clk),
    .D(_01406_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[7][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27609_ (.CLK(clk),
    .D(_01407_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[7][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27610_ (.CLK(clk),
    .D(_01408_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[7][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27611_ (.CLK(clk),
    .D(_01409_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[7][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27612_ (.CLK(clk),
    .D(_01410_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27613_ (.CLK(clk),
    .D(_01411_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27614_ (.CLK(clk),
    .D(_01412_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27615_ (.CLK(clk),
    .D(_01413_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27616_ (.CLK(clk),
    .D(_01414_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27617_ (.CLK(clk),
    .D(_01415_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27618_ (.CLK(clk),
    .D(_01416_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27619_ (.CLK(clk),
    .D(_01417_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27620_ (.CLK(clk),
    .D(_01418_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27621_ (.CLK(clk),
    .D(_01419_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27622_ (.CLK(clk),
    .D(_01420_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27623_ (.CLK(clk),
    .D(_01421_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27624_ (.CLK(clk),
    .D(_01422_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27625_ (.CLK(clk),
    .D(_01423_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27626_ (.CLK(clk),
    .D(_01424_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27627_ (.CLK(clk),
    .D(_01425_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[2].col_loop[0].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27628_ (.CLK(clk),
    .D(_01426_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27629_ (.CLK(clk),
    .D(_01427_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27630_ (.CLK(clk),
    .D(_01428_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27631_ (.CLK(clk),
    .D(_01429_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27632_ (.CLK(clk),
    .D(_01430_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27633_ (.CLK(clk),
    .D(_01431_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27634_ (.CLK(clk),
    .D(_01432_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27635_ (.CLK(clk),
    .D(_01433_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27636_ (.CLK(clk),
    .D(_01434_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27637_ (.CLK(clk),
    .D(_01435_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27638_ (.CLK(clk),
    .D(_01436_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27639_ (.CLK(clk),
    .D(_01437_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27640_ (.CLK(clk),
    .D(_01438_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27641_ (.CLK(clk),
    .D(_01439_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27642_ (.CLK(clk),
    .D(_01440_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27643_ (.CLK(clk),
    .D(_01441_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27644_ (.CLK(clk),
    .D(_01442_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27645_ (.CLK(clk),
    .D(_01443_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27646_ (.CLK(clk),
    .D(_01444_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27647_ (.CLK(clk),
    .D(_01445_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27648_ (.CLK(clk),
    .D(_01446_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27649_ (.CLK(clk),
    .D(_01447_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27650_ (.CLK(clk),
    .D(_01448_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27651_ (.CLK(clk),
    .D(_01449_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27652_ (.CLK(clk),
    .D(_01450_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27653_ (.CLK(clk),
    .D(_01451_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27654_ (.CLK(clk),
    .D(_01452_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27655_ (.CLK(clk),
    .D(_01453_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27656_ (.CLK(clk),
    .D(_01454_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27657_ (.CLK(clk),
    .D(_01455_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27658_ (.CLK(clk),
    .D(_01456_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27659_ (.CLK(clk),
    .D(_01457_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[8][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27660_ (.CLK(clk),
    .D(_01458_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[7][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27661_ (.CLK(clk),
    .D(_01459_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[7][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27662_ (.CLK(clk),
    .D(_01460_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[7][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27663_ (.CLK(clk),
    .D(_01461_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[7][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27664_ (.CLK(clk),
    .D(_01462_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[7][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27665_ (.CLK(clk),
    .D(_01463_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[7][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27666_ (.CLK(clk),
    .D(_01464_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[7][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27667_ (.CLK(clk),
    .D(_01465_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[7][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27668_ (.CLK(clk),
    .D(_01466_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[6][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27669_ (.CLK(clk),
    .D(_01467_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[6][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27670_ (.CLK(clk),
    .D(_01468_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[6][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27671_ (.CLK(clk),
    .D(_01469_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[6][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27672_ (.CLK(clk),
    .D(_01470_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[6][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27673_ (.CLK(clk),
    .D(_01471_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[6][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27674_ (.CLK(clk),
    .D(_01472_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[6][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27675_ (.CLK(clk),
    .D(_01473_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[6][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27676_ (.CLK(clk),
    .D(_01474_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27677_ (.CLK(clk),
    .D(_01475_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27678_ (.CLK(clk),
    .D(_01476_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27679_ (.CLK(clk),
    .D(_01477_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27680_ (.CLK(clk),
    .D(_01478_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27681_ (.CLK(clk),
    .D(_01479_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27682_ (.CLK(clk),
    .D(_01480_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27683_ (.CLK(clk),
    .D(_01481_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27684_ (.CLK(clk),
    .D(_01482_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27685_ (.CLK(clk),
    .D(_01483_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27686_ (.CLK(clk),
    .D(_01484_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27687_ (.CLK(clk),
    .D(_01485_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27688_ (.CLK(clk),
    .D(_01486_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27689_ (.CLK(clk),
    .D(_01487_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27690_ (.CLK(clk),
    .D(_01488_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27691_ (.CLK(clk),
    .D(_01489_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[3].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27692_ (.CLK(clk),
    .D(_01490_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27693_ (.CLK(clk),
    .D(_01491_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27694_ (.CLK(clk),
    .D(_01492_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27695_ (.CLK(clk),
    .D(_01493_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27696_ (.CLK(clk),
    .D(_01494_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27697_ (.CLK(clk),
    .D(_01495_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27698_ (.CLK(clk),
    .D(_01496_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27699_ (.CLK(clk),
    .D(_01497_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27700_ (.CLK(clk),
    .D(_01498_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27701_ (.CLK(clk),
    .D(_01499_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27702_ (.CLK(clk),
    .D(_01500_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27703_ (.CLK(clk),
    .D(_01501_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27704_ (.CLK(clk),
    .D(_01502_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27705_ (.CLK(clk),
    .D(_01503_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27706_ (.CLK(clk),
    .D(_01504_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27707_ (.CLK(clk),
    .D(_01505_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27708_ (.CLK(clk),
    .D(_01506_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27709_ (.CLK(clk),
    .D(_01507_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27710_ (.CLK(clk),
    .D(_01508_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27711_ (.CLK(clk),
    .D(_01509_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27712_ (.CLK(clk),
    .D(_01510_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27713_ (.CLK(clk),
    .D(_01511_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27714_ (.CLK(clk),
    .D(_01512_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27715_ (.CLK(clk),
    .D(_01513_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27716_ (.CLK(clk),
    .D(_01514_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27717_ (.CLK(clk),
    .D(_01515_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27718_ (.CLK(clk),
    .D(_01516_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27719_ (.CLK(clk),
    .D(_01517_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27720_ (.CLK(clk),
    .D(_01518_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27721_ (.CLK(clk),
    .D(_01519_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27722_ (.CLK(clk),
    .D(_01520_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27723_ (.CLK(clk),
    .D(_01521_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[7][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27724_ (.CLK(clk),
    .D(_01522_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[6][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27725_ (.CLK(clk),
    .D(_01523_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[6][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27726_ (.CLK(clk),
    .D(_01524_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[6][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27727_ (.CLK(clk),
    .D(_01525_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[6][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27728_ (.CLK(clk),
    .D(_01526_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[6][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27729_ (.CLK(clk),
    .D(_01527_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[6][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27730_ (.CLK(clk),
    .D(_01528_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[6][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27731_ (.CLK(clk),
    .D(_01529_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[6][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27732_ (.CLK(clk),
    .D(_01530_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[5][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27733_ (.CLK(clk),
    .D(_01531_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[5][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27734_ (.CLK(clk),
    .D(_01532_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[5][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27735_ (.CLK(clk),
    .D(_01533_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[5][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27736_ (.CLK(clk),
    .D(_01534_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[5][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27737_ (.CLK(clk),
    .D(_01535_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[5][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27738_ (.CLK(clk),
    .D(_01536_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[5][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27739_ (.CLK(clk),
    .D(_01537_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[5][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27740_ (.CLK(clk),
    .D(_01538_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27741_ (.CLK(clk),
    .D(_01539_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27742_ (.CLK(clk),
    .D(_01540_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27743_ (.CLK(clk),
    .D(_01541_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27744_ (.CLK(clk),
    .D(_01542_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27745_ (.CLK(clk),
    .D(_01543_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27746_ (.CLK(clk),
    .D(_01544_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27747_ (.CLK(clk),
    .D(_01545_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27748_ (.CLK(clk),
    .D(_01546_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27749_ (.CLK(clk),
    .D(_01547_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27750_ (.CLK(clk),
    .D(_01548_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27751_ (.CLK(clk),
    .D(_01549_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27752_ (.CLK(clk),
    .D(_01550_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27753_ (.CLK(clk),
    .D(_01551_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27754_ (.CLK(clk),
    .D(_01552_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27755_ (.CLK(clk),
    .D(_01553_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[2].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27756_ (.CLK(clk),
    .D(_01554_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27757_ (.CLK(clk),
    .D(_01555_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27758_ (.CLK(clk),
    .D(_01556_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27759_ (.CLK(clk),
    .D(_01557_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27760_ (.CLK(clk),
    .D(_01558_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27761_ (.CLK(clk),
    .D(_01559_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27762_ (.CLK(clk),
    .D(_01560_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27763_ (.CLK(clk),
    .D(_01561_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27764_ (.CLK(clk),
    .D(_01562_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27765_ (.CLK(clk),
    .D(_01563_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27766_ (.CLK(clk),
    .D(_01564_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27767_ (.CLK(clk),
    .D(_01565_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27768_ (.CLK(clk),
    .D(_01566_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27769_ (.CLK(clk),
    .D(_01567_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27770_ (.CLK(clk),
    .D(_01568_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27771_ (.CLK(clk),
    .D(_01569_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27772_ (.CLK(clk),
    .D(_01570_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27773_ (.CLK(clk),
    .D(_01571_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27774_ (.CLK(clk),
    .D(_01572_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27775_ (.CLK(clk),
    .D(_01573_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27776_ (.CLK(clk),
    .D(_01574_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27777_ (.CLK(clk),
    .D(_01575_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27778_ (.CLK(clk),
    .D(_01576_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27779_ (.CLK(clk),
    .D(_01577_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27780_ (.CLK(clk),
    .D(_01578_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27781_ (.CLK(clk),
    .D(_01579_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27782_ (.CLK(clk),
    .D(_01580_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27783_ (.CLK(clk),
    .D(_01581_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27784_ (.CLK(clk),
    .D(_01582_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27785_ (.CLK(clk),
    .D(_01583_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27786_ (.CLK(clk),
    .D(_01584_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27787_ (.CLK(clk),
    .D(_01585_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[6][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27788_ (.CLK(clk),
    .D(_01586_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[5][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27789_ (.CLK(clk),
    .D(_01587_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[5][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27790_ (.CLK(clk),
    .D(_01588_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[5][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27791_ (.CLK(clk),
    .D(_01589_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[5][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27792_ (.CLK(clk),
    .D(_01590_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[5][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27793_ (.CLK(clk),
    .D(_01591_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[5][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27794_ (.CLK(clk),
    .D(_01592_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[5][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27795_ (.CLK(clk),
    .D(_01593_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[5][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27796_ (.CLK(clk),
    .D(_01594_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[4][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27797_ (.CLK(clk),
    .D(_01595_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[4][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27798_ (.CLK(clk),
    .D(_01596_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[4][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27799_ (.CLK(clk),
    .D(_01597_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[4][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27800_ (.CLK(clk),
    .D(_01598_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[4][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27801_ (.CLK(clk),
    .D(_01599_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[4][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27802_ (.CLK(clk),
    .D(_01600_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[4][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27803_ (.CLK(clk),
    .D(_01601_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[4][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27804_ (.CLK(clk),
    .D(_01602_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27805_ (.CLK(clk),
    .D(_01603_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27806_ (.CLK(clk),
    .D(_01604_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27807_ (.CLK(clk),
    .D(_01605_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27808_ (.CLK(clk),
    .D(_01606_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27809_ (.CLK(clk),
    .D(_01607_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27810_ (.CLK(clk),
    .D(_01608_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27811_ (.CLK(clk),
    .D(_01609_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27812_ (.CLK(clk),
    .D(_01610_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27813_ (.CLK(clk),
    .D(_01611_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27814_ (.CLK(clk),
    .D(_01612_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27815_ (.CLK(clk),
    .D(_01613_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27816_ (.CLK(clk),
    .D(_01614_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27817_ (.CLK(clk),
    .D(_01615_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27818_ (.CLK(clk),
    .D(_01616_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27819_ (.CLK(clk),
    .D(_01617_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[1].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27820_ (.CLK(clk),
    .D(_01618_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27821_ (.CLK(clk),
    .D(_01619_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27822_ (.CLK(clk),
    .D(_01620_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27823_ (.CLK(clk),
    .D(_01621_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27824_ (.CLK(clk),
    .D(_01622_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27825_ (.CLK(clk),
    .D(_01623_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27826_ (.CLK(clk),
    .D(_01624_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27827_ (.CLK(clk),
    .D(_01625_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27828_ (.CLK(clk),
    .D(_01626_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27829_ (.CLK(clk),
    .D(_01627_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27830_ (.CLK(clk),
    .D(_01628_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27831_ (.CLK(clk),
    .D(_01629_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27832_ (.CLK(clk),
    .D(_01630_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27833_ (.CLK(clk),
    .D(_01631_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27834_ (.CLK(clk),
    .D(_01632_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27835_ (.CLK(clk),
    .D(_01633_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27836_ (.CLK(clk),
    .D(_01634_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27837_ (.CLK(clk),
    .D(_01635_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27838_ (.CLK(clk),
    .D(_01636_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27839_ (.CLK(clk),
    .D(_01637_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27840_ (.CLK(clk),
    .D(_01638_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27841_ (.CLK(clk),
    .D(_01639_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27842_ (.CLK(clk),
    .D(_01640_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27843_ (.CLK(clk),
    .D(_01641_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27844_ (.CLK(clk),
    .D(_01642_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27845_ (.CLK(clk),
    .D(_01643_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27846_ (.CLK(clk),
    .D(_01644_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27847_ (.CLK(clk),
    .D(_01645_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27848_ (.CLK(clk),
    .D(_01646_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27849_ (.CLK(clk),
    .D(_01647_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27850_ (.CLK(clk),
    .D(_01648_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27851_ (.CLK(clk),
    .D(_01649_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[5][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27852_ (.CLK(clk),
    .D(_01650_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[4][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27853_ (.CLK(clk),
    .D(_01651_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[4][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27854_ (.CLK(clk),
    .D(_01652_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[4][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27855_ (.CLK(clk),
    .D(_01653_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[4][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27856_ (.CLK(clk),
    .D(_01654_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[4][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27857_ (.CLK(clk),
    .D(_01655_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[4][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27858_ (.CLK(clk),
    .D(_01656_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[4][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27859_ (.CLK(clk),
    .D(_01657_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[4][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27860_ (.CLK(clk),
    .D(_01658_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[3][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27861_ (.CLK(clk),
    .D(_01659_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[3][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27862_ (.CLK(clk),
    .D(_01660_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[3][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27863_ (.CLK(clk),
    .D(_01661_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[3][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27864_ (.CLK(clk),
    .D(_01662_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[3][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27865_ (.CLK(clk),
    .D(_01663_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[3][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27866_ (.CLK(clk),
    .D(_01664_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[3][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27867_ (.CLK(clk),
    .D(_01665_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[3][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27868_ (.CLK(clk),
    .D(_01666_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27869_ (.CLK(clk),
    .D(_01667_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27870_ (.CLK(clk),
    .D(_01668_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27871_ (.CLK(clk),
    .D(_01669_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27872_ (.CLK(clk),
    .D(_01670_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27873_ (.CLK(clk),
    .D(_01671_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27874_ (.CLK(clk),
    .D(_01672_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27875_ (.CLK(clk),
    .D(_01673_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27876_ (.CLK(clk),
    .D(_01674_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27877_ (.CLK(clk),
    .D(_01675_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27878_ (.CLK(clk),
    .D(_01676_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27879_ (.CLK(clk),
    .D(_01677_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27880_ (.CLK(clk),
    .D(_01678_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27881_ (.CLK(clk),
    .D(_01679_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27882_ (.CLK(clk),
    .D(_01680_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27883_ (.CLK(clk),
    .D(_01681_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[1].col_loop[0].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27884_ (.CLK(clk),
    .D(_01682_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27885_ (.CLK(clk),
    .D(_01683_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27886_ (.CLK(clk),
    .D(_01684_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27887_ (.CLK(clk),
    .D(_01685_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27888_ (.CLK(clk),
    .D(_01686_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27889_ (.CLK(clk),
    .D(_01687_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27890_ (.CLK(clk),
    .D(_01688_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27891_ (.CLK(clk),
    .D(_01689_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27892_ (.CLK(clk),
    .D(_01690_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27893_ (.CLK(clk),
    .D(_01691_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27894_ (.CLK(clk),
    .D(_01692_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27895_ (.CLK(clk),
    .D(_01693_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27896_ (.CLK(clk),
    .D(_01694_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27897_ (.CLK(clk),
    .D(_01695_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27898_ (.CLK(clk),
    .D(_01696_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27899_ (.CLK(clk),
    .D(_01697_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27900_ (.CLK(clk),
    .D(_01698_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27901_ (.CLK(clk),
    .D(_01699_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27902_ (.CLK(clk),
    .D(_01700_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27903_ (.CLK(clk),
    .D(_01701_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27904_ (.CLK(clk),
    .D(_01702_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27905_ (.CLK(clk),
    .D(_01703_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27906_ (.CLK(clk),
    .D(_01704_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27907_ (.CLK(clk),
    .D(_01705_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27908_ (.CLK(clk),
    .D(_01706_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27909_ (.CLK(clk),
    .D(_01707_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27910_ (.CLK(clk),
    .D(_01708_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27911_ (.CLK(clk),
    .D(_01709_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27912_ (.CLK(clk),
    .D(_01710_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27913_ (.CLK(clk),
    .D(_01711_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27914_ (.CLK(clk),
    .D(_01712_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27915_ (.CLK(clk),
    .D(_01713_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[4][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27916_ (.CLK(clk),
    .D(_01714_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[3][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27917_ (.CLK(clk),
    .D(_01715_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[3][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27918_ (.CLK(clk),
    .D(_01716_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[3][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27919_ (.CLK(clk),
    .D(_01717_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[3][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27920_ (.CLK(clk),
    .D(_01718_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[3][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27921_ (.CLK(clk),
    .D(_01719_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[3][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27922_ (.CLK(clk),
    .D(_01720_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[3][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27923_ (.CLK(clk),
    .D(_01721_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[3][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27924_ (.CLK(clk),
    .D(_01722_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[2][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27925_ (.CLK(clk),
    .D(_01723_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[2][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27926_ (.CLK(clk),
    .D(_01724_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[2][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27927_ (.CLK(clk),
    .D(_01725_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[2][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27928_ (.CLK(clk),
    .D(_01726_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[2][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27929_ (.CLK(clk),
    .D(_01727_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[2][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27930_ (.CLK(clk),
    .D(_01728_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[2][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27931_ (.CLK(clk),
    .D(_01729_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[2][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27932_ (.CLK(clk),
    .D(_01730_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27933_ (.CLK(clk),
    .D(_01731_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27934_ (.CLK(clk),
    .D(_01732_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27935_ (.CLK(clk),
    .D(_01733_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27936_ (.CLK(clk),
    .D(_01734_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27937_ (.CLK(clk),
    .D(_01735_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27938_ (.CLK(clk),
    .D(_01736_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27939_ (.CLK(clk),
    .D(_01737_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27940_ (.CLK(clk),
    .D(_01738_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27941_ (.CLK(clk),
    .D(_01739_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27942_ (.CLK(clk),
    .D(_01740_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _27943_ (.CLK(clk),
    .D(_01741_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _27944_ (.CLK(clk),
    .D(_01742_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _27945_ (.CLK(clk),
    .D(_01743_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _27946_ (.CLK(clk),
    .D(_01744_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _27947_ (.CLK(clk),
    .D(_01745_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[3].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27948_ (.CLK(clk),
    .D(_01746_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27949_ (.CLK(clk),
    .D(_01747_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27950_ (.CLK(clk),
    .D(_01748_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27951_ (.CLK(clk),
    .D(_01749_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27952_ (.CLK(clk),
    .D(_01750_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27953_ (.CLK(clk),
    .D(_01751_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27954_ (.CLK(clk),
    .D(_01752_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27955_ (.CLK(clk),
    .D(_01753_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27956_ (.CLK(clk),
    .D(_01754_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][8] ));
 sky130_fd_sc_hd__dfrtp_2 _27957_ (.CLK(clk),
    .D(_01755_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][9] ));
 sky130_fd_sc_hd__dfrtp_2 _27958_ (.CLK(clk),
    .D(_01756_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][10] ));
 sky130_fd_sc_hd__dfrtp_2 _27959_ (.CLK(clk),
    .D(_01757_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][11] ));
 sky130_fd_sc_hd__dfrtp_2 _27960_ (.CLK(clk),
    .D(_01758_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][12] ));
 sky130_fd_sc_hd__dfrtp_2 _27961_ (.CLK(clk),
    .D(_01759_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][13] ));
 sky130_fd_sc_hd__dfrtp_2 _27962_ (.CLK(clk),
    .D(_01760_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][14] ));
 sky130_fd_sc_hd__dfrtp_2 _27963_ (.CLK(clk),
    .D(_01761_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][15] ));
 sky130_fd_sc_hd__dfrtp_2 _27964_ (.CLK(clk),
    .D(_01762_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][16] ));
 sky130_fd_sc_hd__dfrtp_2 _27965_ (.CLK(clk),
    .D(_01763_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][17] ));
 sky130_fd_sc_hd__dfrtp_2 _27966_ (.CLK(clk),
    .D(_01764_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][18] ));
 sky130_fd_sc_hd__dfrtp_2 _27967_ (.CLK(clk),
    .D(_01765_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][19] ));
 sky130_fd_sc_hd__dfrtp_2 _27968_ (.CLK(clk),
    .D(_01766_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][20] ));
 sky130_fd_sc_hd__dfrtp_2 _27969_ (.CLK(clk),
    .D(_01767_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][21] ));
 sky130_fd_sc_hd__dfrtp_2 _27970_ (.CLK(clk),
    .D(_01768_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][22] ));
 sky130_fd_sc_hd__dfrtp_2 _27971_ (.CLK(clk),
    .D(_01769_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][23] ));
 sky130_fd_sc_hd__dfrtp_2 _27972_ (.CLK(clk),
    .D(_01770_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][24] ));
 sky130_fd_sc_hd__dfrtp_2 _27973_ (.CLK(clk),
    .D(_01771_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][25] ));
 sky130_fd_sc_hd__dfrtp_2 _27974_ (.CLK(clk),
    .D(_01772_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][26] ));
 sky130_fd_sc_hd__dfrtp_2 _27975_ (.CLK(clk),
    .D(_01773_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][27] ));
 sky130_fd_sc_hd__dfrtp_2 _27976_ (.CLK(clk),
    .D(_01774_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][28] ));
 sky130_fd_sc_hd__dfrtp_2 _27977_ (.CLK(clk),
    .D(_01775_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][29] ));
 sky130_fd_sc_hd__dfrtp_2 _27978_ (.CLK(clk),
    .D(_01776_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][30] ));
 sky130_fd_sc_hd__dfrtp_2 _27979_ (.CLK(clk),
    .D(_01777_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[3][31] ));
 sky130_fd_sc_hd__dfrtp_2 _27980_ (.CLK(clk),
    .D(_01778_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[2][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27981_ (.CLK(clk),
    .D(_01779_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[2][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27982_ (.CLK(clk),
    .D(_01780_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[2][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27983_ (.CLK(clk),
    .D(_01781_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[2][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27984_ (.CLK(clk),
    .D(_01782_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[2][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27985_ (.CLK(clk),
    .D(_01783_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[2][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27986_ (.CLK(clk),
    .D(_01784_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[2][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27987_ (.CLK(clk),
    .D(_01785_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[2][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27988_ (.CLK(clk),
    .D(_01786_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[1][0] ));
 sky130_fd_sc_hd__dfrtp_2 _27989_ (.CLK(clk),
    .D(_01787_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[1][1] ));
 sky130_fd_sc_hd__dfrtp_2 _27990_ (.CLK(clk),
    .D(_01788_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[1][2] ));
 sky130_fd_sc_hd__dfrtp_2 _27991_ (.CLK(clk),
    .D(_01789_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[1][3] ));
 sky130_fd_sc_hd__dfrtp_2 _27992_ (.CLK(clk),
    .D(_01790_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[1][4] ));
 sky130_fd_sc_hd__dfrtp_2 _27993_ (.CLK(clk),
    .D(_01791_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[1][5] ));
 sky130_fd_sc_hd__dfrtp_2 _27994_ (.CLK(clk),
    .D(_01792_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[1][6] ));
 sky130_fd_sc_hd__dfrtp_2 _27995_ (.CLK(clk),
    .D(_01793_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[1][7] ));
 sky130_fd_sc_hd__dfrtp_2 _27996_ (.CLK(clk),
    .D(_01794_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27997_ (.CLK(clk),
    .D(_01795_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27998_ (.CLK(clk),
    .D(_01796_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27999_ (.CLK(clk),
    .D(_01797_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _28000_ (.CLK(clk),
    .D(_01798_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _28001_ (.CLK(clk),
    .D(_01799_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _28002_ (.CLK(clk),
    .D(_01800_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _28003_ (.CLK(clk),
    .D(_01801_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _28004_ (.CLK(clk),
    .D(_01802_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _28005_ (.CLK(clk),
    .D(_01803_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _28006_ (.CLK(clk),
    .D(_01804_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _28007_ (.CLK(clk),
    .D(_01805_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _28008_ (.CLK(clk),
    .D(_01806_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _28009_ (.CLK(clk),
    .D(_01807_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _28010_ (.CLK(clk),
    .D(_01808_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _28011_ (.CLK(clk),
    .D(_01809_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[2].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _28012_ (.CLK(clk),
    .D(_01810_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][0] ));
 sky130_fd_sc_hd__dfrtp_2 _28013_ (.CLK(clk),
    .D(_01811_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][1] ));
 sky130_fd_sc_hd__dfrtp_2 _28014_ (.CLK(clk),
    .D(_01812_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][2] ));
 sky130_fd_sc_hd__dfrtp_2 _28015_ (.CLK(clk),
    .D(_01813_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][3] ));
 sky130_fd_sc_hd__dfrtp_2 _28016_ (.CLK(clk),
    .D(_01814_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][4] ));
 sky130_fd_sc_hd__dfrtp_2 _28017_ (.CLK(clk),
    .D(_01815_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][5] ));
 sky130_fd_sc_hd__dfrtp_2 _28018_ (.CLK(clk),
    .D(_01816_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][6] ));
 sky130_fd_sc_hd__dfrtp_2 _28019_ (.CLK(clk),
    .D(_01817_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28020_ (.CLK(clk),
    .D(_01818_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][8] ));
 sky130_fd_sc_hd__dfrtp_2 _28021_ (.CLK(clk),
    .D(_01819_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][9] ));
 sky130_fd_sc_hd__dfrtp_2 _28022_ (.CLK(clk),
    .D(_01820_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][10] ));
 sky130_fd_sc_hd__dfrtp_2 _28023_ (.CLK(clk),
    .D(_01821_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][11] ));
 sky130_fd_sc_hd__dfrtp_2 _28024_ (.CLK(clk),
    .D(_01822_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][12] ));
 sky130_fd_sc_hd__dfrtp_2 _28025_ (.CLK(clk),
    .D(_01823_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][13] ));
 sky130_fd_sc_hd__dfrtp_2 _28026_ (.CLK(clk),
    .D(_01824_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][14] ));
 sky130_fd_sc_hd__dfrtp_2 _28027_ (.CLK(clk),
    .D(_01825_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][15] ));
 sky130_fd_sc_hd__dfrtp_2 _28028_ (.CLK(clk),
    .D(_01826_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][16] ));
 sky130_fd_sc_hd__dfrtp_2 _28029_ (.CLK(clk),
    .D(_01827_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][17] ));
 sky130_fd_sc_hd__dfrtp_2 _28030_ (.CLK(clk),
    .D(_01828_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][18] ));
 sky130_fd_sc_hd__dfrtp_2 _28031_ (.CLK(clk),
    .D(_01829_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][19] ));
 sky130_fd_sc_hd__dfrtp_2 _28032_ (.CLK(clk),
    .D(_01830_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][20] ));
 sky130_fd_sc_hd__dfrtp_2 _28033_ (.CLK(clk),
    .D(_01831_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][21] ));
 sky130_fd_sc_hd__dfrtp_2 _28034_ (.CLK(clk),
    .D(_01832_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][22] ));
 sky130_fd_sc_hd__dfrtp_2 _28035_ (.CLK(clk),
    .D(_01833_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][23] ));
 sky130_fd_sc_hd__dfrtp_2 _28036_ (.CLK(clk),
    .D(_01834_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][24] ));
 sky130_fd_sc_hd__dfrtp_2 _28037_ (.CLK(clk),
    .D(_01835_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][25] ));
 sky130_fd_sc_hd__dfrtp_2 _28038_ (.CLK(clk),
    .D(_01836_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][26] ));
 sky130_fd_sc_hd__dfrtp_2 _28039_ (.CLK(clk),
    .D(_01837_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][27] ));
 sky130_fd_sc_hd__dfrtp_2 _28040_ (.CLK(clk),
    .D(_01838_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][28] ));
 sky130_fd_sc_hd__dfrtp_2 _28041_ (.CLK(clk),
    .D(_01839_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][29] ));
 sky130_fd_sc_hd__dfrtp_2 _28042_ (.CLK(clk),
    .D(_01840_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][30] ));
 sky130_fd_sc_hd__dfrtp_2 _28043_ (.CLK(clk),
    .D(_01841_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[2][31] ));
 sky130_fd_sc_hd__dfrtp_2 _28044_ (.CLK(clk),
    .D(_01842_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[1][0] ));
 sky130_fd_sc_hd__dfrtp_2 _28045_ (.CLK(clk),
    .D(_01843_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[1][1] ));
 sky130_fd_sc_hd__dfrtp_2 _28046_ (.CLK(clk),
    .D(_01844_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[1][2] ));
 sky130_fd_sc_hd__dfrtp_2 _28047_ (.CLK(clk),
    .D(_01845_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[1][3] ));
 sky130_fd_sc_hd__dfrtp_2 _28048_ (.CLK(clk),
    .D(_01846_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[1][4] ));
 sky130_fd_sc_hd__dfrtp_2 _28049_ (.CLK(clk),
    .D(_01847_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[1][5] ));
 sky130_fd_sc_hd__dfrtp_2 _28050_ (.CLK(clk),
    .D(_01848_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[1][6] ));
 sky130_fd_sc_hd__dfrtp_2 _28051_ (.CLK(clk),
    .D(_01849_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[1][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28052_ (.CLK(clk),
    .D(_01850_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _28053_ (.CLK(clk),
    .D(_01851_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _28054_ (.CLK(clk),
    .D(_01852_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _28055_ (.CLK(clk),
    .D(_01853_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _28056_ (.CLK(clk),
    .D(_01854_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _28057_ (.CLK(clk),
    .D(_01855_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _28058_ (.CLK(clk),
    .D(_01856_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _28059_ (.CLK(clk),
    .D(_01857_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28060_ (.CLK(clk),
    .D(_01858_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _28061_ (.CLK(clk),
    .D(_01859_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _28062_ (.CLK(clk),
    .D(_01860_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _28063_ (.CLK(clk),
    .D(_01861_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _28064_ (.CLK(clk),
    .D(_01862_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _28065_ (.CLK(clk),
    .D(_01863_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _28066_ (.CLK(clk),
    .D(_01864_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _28067_ (.CLK(clk),
    .D(_01865_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _28068_ (.CLK(clk),
    .D(_01866_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _28069_ (.CLK(clk),
    .D(_01867_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _28070_ (.CLK(clk),
    .D(_01868_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _28071_ (.CLK(clk),
    .D(_01869_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _28072_ (.CLK(clk),
    .D(_01870_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _28073_ (.CLK(clk),
    .D(_01871_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _28074_ (.CLK(clk),
    .D(_01872_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _28075_ (.CLK(clk),
    .D(_01873_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[1].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _28076_ (.CLK(clk),
    .D(_01874_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][0] ));
 sky130_fd_sc_hd__dfrtp_2 _28077_ (.CLK(clk),
    .D(_01875_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][1] ));
 sky130_fd_sc_hd__dfrtp_2 _28078_ (.CLK(clk),
    .D(_01876_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][2] ));
 sky130_fd_sc_hd__dfrtp_2 _28079_ (.CLK(clk),
    .D(_01877_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][3] ));
 sky130_fd_sc_hd__dfrtp_2 _28080_ (.CLK(clk),
    .D(_01878_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][4] ));
 sky130_fd_sc_hd__dfrtp_2 _28081_ (.CLK(clk),
    .D(_01879_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][5] ));
 sky130_fd_sc_hd__dfrtp_2 _28082_ (.CLK(clk),
    .D(_01880_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][6] ));
 sky130_fd_sc_hd__dfrtp_2 _28083_ (.CLK(clk),
    .D(_01881_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28084_ (.CLK(clk),
    .D(_01882_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][8] ));
 sky130_fd_sc_hd__dfrtp_2 _28085_ (.CLK(clk),
    .D(_01883_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][9] ));
 sky130_fd_sc_hd__dfrtp_2 _28086_ (.CLK(clk),
    .D(_01884_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][10] ));
 sky130_fd_sc_hd__dfrtp_2 _28087_ (.CLK(clk),
    .D(_01885_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][11] ));
 sky130_fd_sc_hd__dfrtp_2 _28088_ (.CLK(clk),
    .D(_01886_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][12] ));
 sky130_fd_sc_hd__dfrtp_2 _28089_ (.CLK(clk),
    .D(_01887_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][13] ));
 sky130_fd_sc_hd__dfrtp_2 _28090_ (.CLK(clk),
    .D(_01888_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][14] ));
 sky130_fd_sc_hd__dfrtp_2 _28091_ (.CLK(clk),
    .D(_01889_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][15] ));
 sky130_fd_sc_hd__dfrtp_2 _28092_ (.CLK(clk),
    .D(_01890_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][16] ));
 sky130_fd_sc_hd__dfrtp_2 _28093_ (.CLK(clk),
    .D(_01891_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][17] ));
 sky130_fd_sc_hd__dfrtp_2 _28094_ (.CLK(clk),
    .D(_01892_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][18] ));
 sky130_fd_sc_hd__dfrtp_2 _28095_ (.CLK(clk),
    .D(_01893_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][19] ));
 sky130_fd_sc_hd__dfrtp_2 _28096_ (.CLK(clk),
    .D(_01894_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][20] ));
 sky130_fd_sc_hd__dfrtp_2 _28097_ (.CLK(clk),
    .D(_01895_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][21] ));
 sky130_fd_sc_hd__dfrtp_2 _28098_ (.CLK(clk),
    .D(_01896_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][22] ));
 sky130_fd_sc_hd__dfrtp_2 _28099_ (.CLK(clk),
    .D(_01897_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][23] ));
 sky130_fd_sc_hd__dfrtp_2 _28100_ (.CLK(clk),
    .D(_01898_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][24] ));
 sky130_fd_sc_hd__dfrtp_2 _28101_ (.CLK(clk),
    .D(_01899_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][25] ));
 sky130_fd_sc_hd__dfrtp_2 _28102_ (.CLK(clk),
    .D(_01900_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][26] ));
 sky130_fd_sc_hd__dfrtp_2 _28103_ (.CLK(clk),
    .D(_01901_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][27] ));
 sky130_fd_sc_hd__dfrtp_2 _28104_ (.CLK(clk),
    .D(_01902_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][28] ));
 sky130_fd_sc_hd__dfrtp_2 _28105_ (.CLK(clk),
    .D(_01903_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][29] ));
 sky130_fd_sc_hd__dfrtp_2 _28106_ (.CLK(clk),
    .D(_01904_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][30] ));
 sky130_fd_sc_hd__dfrtp_2 _28107_ (.CLK(clk),
    .D(_01905_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[1][31] ));
 sky130_fd_sc_hd__dfrtp_2 _28108_ (.CLK(clk),
    .D(_01906_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _28109_ (.CLK(clk),
    .D(_01907_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _28110_ (.CLK(clk),
    .D(_01908_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _28111_ (.CLK(clk),
    .D(_01909_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _28112_ (.CLK(clk),
    .D(_01910_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _28113_ (.CLK(clk),
    .D(_01911_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _28114_ (.CLK(clk),
    .D(_01912_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _28115_ (.CLK(clk),
    .D(_01913_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.A_outs[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28116_ (.CLK(clk),
    .D(_01914_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _28117_ (.CLK(clk),
    .D(_01915_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _28118_ (.CLK(clk),
    .D(_01916_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _28119_ (.CLK(clk),
    .D(_01917_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _28120_ (.CLK(clk),
    .D(_01918_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _28121_ (.CLK(clk),
    .D(_01919_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _28122_ (.CLK(clk),
    .D(_01920_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _28123_ (.CLK(clk),
    .D(_01921_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _28124_ (.CLK(clk),
    .D(_01922_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _28125_ (.CLK(clk),
    .D(_01923_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _28126_ (.CLK(clk),
    .D(_01924_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _28127_ (.CLK(clk),
    .D(_01925_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _28128_ (.CLK(clk),
    .D(_01926_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _28129_ (.CLK(clk),
    .D(_01927_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _28130_ (.CLK(clk),
    .D(_01928_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _28131_ (.CLK(clk),
    .D(_01929_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.row_loop[0].col_loop[0].pe_i.prod_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _28132_ (.CLK(clk),
    .D(_01930_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _28133_ (.CLK(clk),
    .D(_01931_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _28134_ (.CLK(clk),
    .D(_01932_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _28135_ (.CLK(clk),
    .D(_01933_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _28136_ (.CLK(clk),
    .D(_01934_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _28137_ (.CLK(clk),
    .D(_01935_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _28138_ (.CLK(clk),
    .D(_01936_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _28139_ (.CLK(clk),
    .D(_01937_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28140_ (.CLK(clk),
    .D(_01938_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][8] ));
 sky130_fd_sc_hd__dfrtp_2 _28141_ (.CLK(clk),
    .D(_01939_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][9] ));
 sky130_fd_sc_hd__dfrtp_2 _28142_ (.CLK(clk),
    .D(_01940_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][10] ));
 sky130_fd_sc_hd__dfrtp_2 _28143_ (.CLK(clk),
    .D(_01941_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][11] ));
 sky130_fd_sc_hd__dfrtp_2 _28144_ (.CLK(clk),
    .D(_01942_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][12] ));
 sky130_fd_sc_hd__dfrtp_2 _28145_ (.CLK(clk),
    .D(_01943_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][13] ));
 sky130_fd_sc_hd__dfrtp_2 _28146_ (.CLK(clk),
    .D(_01944_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][14] ));
 sky130_fd_sc_hd__dfrtp_2 _28147_ (.CLK(clk),
    .D(_01945_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][15] ));
 sky130_fd_sc_hd__dfrtp_2 _28148_ (.CLK(clk),
    .D(_01946_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][16] ));
 sky130_fd_sc_hd__dfrtp_2 _28149_ (.CLK(clk),
    .D(_01947_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][17] ));
 sky130_fd_sc_hd__dfrtp_2 _28150_ (.CLK(clk),
    .D(_01948_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][18] ));
 sky130_fd_sc_hd__dfrtp_2 _28151_ (.CLK(clk),
    .D(_01949_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][19] ));
 sky130_fd_sc_hd__dfrtp_2 _28152_ (.CLK(clk),
    .D(_01950_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][20] ));
 sky130_fd_sc_hd__dfrtp_2 _28153_ (.CLK(clk),
    .D(_01951_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][21] ));
 sky130_fd_sc_hd__dfrtp_2 _28154_ (.CLK(clk),
    .D(_01952_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][22] ));
 sky130_fd_sc_hd__dfrtp_2 _28155_ (.CLK(clk),
    .D(_01953_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][23] ));
 sky130_fd_sc_hd__dfrtp_2 _28156_ (.CLK(clk),
    .D(_01954_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][24] ));
 sky130_fd_sc_hd__dfrtp_2 _28157_ (.CLK(clk),
    .D(_01955_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][25] ));
 sky130_fd_sc_hd__dfrtp_2 _28158_ (.CLK(clk),
    .D(_01956_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][26] ));
 sky130_fd_sc_hd__dfrtp_2 _28159_ (.CLK(clk),
    .D(_01957_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][27] ));
 sky130_fd_sc_hd__dfrtp_2 _28160_ (.CLK(clk),
    .D(_01958_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][28] ));
 sky130_fd_sc_hd__dfrtp_2 _28161_ (.CLK(clk),
    .D(_01959_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][29] ));
 sky130_fd_sc_hd__dfrtp_2 _28162_ (.CLK(clk),
    .D(_01960_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][30] ));
 sky130_fd_sc_hd__dfrtp_2 _28163_ (.CLK(clk),
    .D(_01961_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.acc_wires[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28164_ (.CLK(clk),
    .D(_01962_),
    .Q(\systolic_inst.B_shift[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28165_ (.CLK(clk),
    .D(_01963_),
    .Q(\systolic_inst.B_shift[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28166_ (.CLK(clk),
    .D(_01964_),
    .Q(\systolic_inst.B_shift[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28167_ (.CLK(clk),
    .D(_01965_),
    .Q(\systolic_inst.B_shift[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28168_ (.CLK(clk),
    .D(_01966_),
    .Q(\systolic_inst.B_shift[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28169_ (.CLK(clk),
    .D(_01967_),
    .Q(\systolic_inst.B_shift[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28170_ (.CLK(clk),
    .D(_01968_),
    .Q(\systolic_inst.B_shift[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28171_ (.CLK(clk),
    .D(_01969_),
    .Q(\systolic_inst.B_shift[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28172_ (.CLK(clk),
    .D(_01970_),
    .Q(\systolic_inst.B_shift[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28173_ (.CLK(clk),
    .D(_01971_),
    .Q(\systolic_inst.B_shift[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28174_ (.CLK(clk),
    .D(_01972_),
    .Q(\systolic_inst.B_shift[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28175_ (.CLK(clk),
    .D(_01973_),
    .Q(\systolic_inst.B_shift[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28176_ (.CLK(clk),
    .D(_01974_),
    .Q(\systolic_inst.B_shift[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28177_ (.CLK(clk),
    .D(_01975_),
    .Q(\systolic_inst.B_shift[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28178_ (.CLK(clk),
    .D(_01976_),
    .Q(\systolic_inst.B_shift[18][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28179_ (.CLK(clk),
    .D(_01977_),
    .Q(\systolic_inst.B_shift[18][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28180_ (.CLK(clk),
    .D(_01978_),
    .Q(\systolic_inst.A_shift[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28181_ (.CLK(clk),
    .D(_01979_),
    .Q(\systolic_inst.A_shift[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28182_ (.CLK(clk),
    .D(_01980_),
    .Q(\systolic_inst.A_shift[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28183_ (.CLK(clk),
    .D(_01981_),
    .Q(\systolic_inst.A_shift[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28184_ (.CLK(clk),
    .D(_01982_),
    .Q(\systolic_inst.A_shift[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28185_ (.CLK(clk),
    .D(_01983_),
    .Q(\systolic_inst.A_shift[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28186_ (.CLK(clk),
    .D(_01984_),
    .Q(\systolic_inst.A_shift[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28187_ (.CLK(clk),
    .D(_01985_),
    .Q(\systolic_inst.A_shift[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28188_ (.CLK(clk),
    .D(_01986_),
    .Q(\systolic_inst.B_shift[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28189_ (.CLK(clk),
    .D(_01987_),
    .Q(\systolic_inst.B_shift[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28190_ (.CLK(clk),
    .D(_01988_),
    .Q(\systolic_inst.B_shift[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28191_ (.CLK(clk),
    .D(_01989_),
    .Q(\systolic_inst.B_shift[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28192_ (.CLK(clk),
    .D(_01990_),
    .Q(\systolic_inst.B_shift[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28193_ (.CLK(clk),
    .D(_01991_),
    .Q(\systolic_inst.B_shift[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28194_ (.CLK(clk),
    .D(_01992_),
    .Q(\systolic_inst.B_shift[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28195_ (.CLK(clk),
    .D(_01993_),
    .Q(\systolic_inst.B_shift[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28196_ (.CLK(clk),
    .D(_01994_),
    .Q(\systolic_inst.B_shift[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28197_ (.CLK(clk),
    .D(_01995_),
    .Q(\systolic_inst.B_shift[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28198_ (.CLK(clk),
    .D(_01996_),
    .Q(\systolic_inst.B_shift[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28199_ (.CLK(clk),
    .D(_01997_),
    .Q(\systolic_inst.B_shift[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28200_ (.CLK(clk),
    .D(_01998_),
    .Q(\systolic_inst.B_shift[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28201_ (.CLK(clk),
    .D(_01999_),
    .Q(\systolic_inst.B_shift[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28202_ (.CLK(clk),
    .D(_02000_),
    .Q(\systolic_inst.B_shift[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28203_ (.CLK(clk),
    .D(_02001_),
    .Q(\systolic_inst.B_shift[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28204_ (.CLK(clk),
    .D(_02002_),
    .Q(\systolic_inst.B_shift[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28205_ (.CLK(clk),
    .D(_02003_),
    .Q(\systolic_inst.B_shift[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28206_ (.CLK(clk),
    .D(_02004_),
    .Q(\systolic_inst.B_shift[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28207_ (.CLK(clk),
    .D(_02005_),
    .Q(\systolic_inst.B_shift[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28208_ (.CLK(clk),
    .D(_02006_),
    .Q(\systolic_inst.B_shift[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28209_ (.CLK(clk),
    .D(_02007_),
    .Q(\systolic_inst.B_shift[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28210_ (.CLK(clk),
    .D(_02008_),
    .Q(\systolic_inst.B_shift[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28211_ (.CLK(clk),
    .D(_02009_),
    .Q(\systolic_inst.B_shift[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28212_ (.CLK(clk),
    .D(_02010_),
    .Q(\systolic_inst.B_shift[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28213_ (.CLK(clk),
    .D(_02011_),
    .Q(\systolic_inst.B_shift[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28214_ (.CLK(clk),
    .D(_02012_),
    .Q(\systolic_inst.B_shift[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28215_ (.CLK(clk),
    .D(_02013_),
    .Q(\systolic_inst.B_shift[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28216_ (.CLK(clk),
    .D(_02014_),
    .Q(\systolic_inst.B_shift[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28217_ (.CLK(clk),
    .D(_02015_),
    .Q(\systolic_inst.B_shift[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28218_ (.CLK(clk),
    .D(_02016_),
    .Q(\systolic_inst.B_shift[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28219_ (.CLK(clk),
    .D(_02017_),
    .Q(\systolic_inst.B_shift[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28220_ (.CLK(clk),
    .D(_02018_),
    .Q(\systolic_inst.B_shift[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28221_ (.CLK(clk),
    .D(_02019_),
    .Q(\systolic_inst.B_shift[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28222_ (.CLK(clk),
    .D(_02020_),
    .Q(\systolic_inst.B_shift[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28223_ (.CLK(clk),
    .D(_02021_),
    .Q(\systolic_inst.B_shift[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28224_ (.CLK(clk),
    .D(_02022_),
    .Q(\systolic_inst.B_shift[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28225_ (.CLK(clk),
    .D(_02023_),
    .Q(\systolic_inst.B_shift[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28226_ (.CLK(clk),
    .D(_02024_),
    .Q(\systolic_inst.B_shift[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28227_ (.CLK(clk),
    .D(_02025_),
    .Q(\systolic_inst.B_shift[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28228_ (.CLK(clk),
    .D(_02026_),
    .Q(\systolic_inst.B_shift[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28229_ (.CLK(clk),
    .D(_02027_),
    .Q(\systolic_inst.B_shift[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28230_ (.CLK(clk),
    .D(_02028_),
    .Q(\systolic_inst.B_shift[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28231_ (.CLK(clk),
    .D(_02029_),
    .Q(\systolic_inst.B_shift[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28232_ (.CLK(clk),
    .D(_02030_),
    .Q(\systolic_inst.B_shift[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28233_ (.CLK(clk),
    .D(_02031_),
    .Q(\systolic_inst.B_shift[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28234_ (.CLK(clk),
    .D(_02032_),
    .Q(\systolic_inst.B_shift[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28235_ (.CLK(clk),
    .D(_02033_),
    .Q(\systolic_inst.B_shift[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28236_ (.CLK(clk),
    .D(_02034_),
    .Q(\systolic_inst.B_shift[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28237_ (.CLK(clk),
    .D(_02035_),
    .Q(\systolic_inst.B_shift[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28238_ (.CLK(clk),
    .D(_02036_),
    .Q(\systolic_inst.B_shift[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28239_ (.CLK(clk),
    .D(_02037_),
    .Q(\systolic_inst.B_shift[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28240_ (.CLK(clk),
    .D(_02038_),
    .Q(\systolic_inst.B_shift[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28241_ (.CLK(clk),
    .D(_02039_),
    .Q(\systolic_inst.B_shift[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28242_ (.CLK(clk),
    .D(_02040_),
    .Q(\systolic_inst.B_shift[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28243_ (.CLK(clk),
    .D(_02041_),
    .Q(\systolic_inst.B_shift[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28244_ (.CLK(clk),
    .D(_02042_),
    .Q(\systolic_inst.B_shift[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28245_ (.CLK(clk),
    .D(_02043_),
    .Q(\systolic_inst.B_shift[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28246_ (.CLK(clk),
    .D(_02044_),
    .Q(\systolic_inst.B_shift[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28247_ (.CLK(clk),
    .D(_02045_),
    .Q(\systolic_inst.B_shift[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28248_ (.CLK(clk),
    .D(_02046_),
    .Q(\systolic_inst.B_shift[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28249_ (.CLK(clk),
    .D(_02047_),
    .Q(\systolic_inst.B_shift[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28250_ (.CLK(clk),
    .D(_02048_),
    .Q(\systolic_inst.B_shift[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28251_ (.CLK(clk),
    .D(_02049_),
    .Q(\systolic_inst.B_shift[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28252_ (.CLK(clk),
    .D(_02050_),
    .Q(\systolic_inst.B_shift[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28253_ (.CLK(clk),
    .D(_02051_),
    .Q(\systolic_inst.B_shift[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28254_ (.CLK(clk),
    .D(_02052_),
    .Q(\systolic_inst.B_shift[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28255_ (.CLK(clk),
    .D(_02053_),
    .Q(\systolic_inst.B_shift[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28256_ (.CLK(clk),
    .D(_02054_),
    .Q(\systolic_inst.B_shift[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28257_ (.CLK(clk),
    .D(_02055_),
    .Q(\systolic_inst.B_shift[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28258_ (.CLK(clk),
    .D(_02056_),
    .Q(\systolic_inst.B_shift[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28259_ (.CLK(clk),
    .D(_02057_),
    .Q(\systolic_inst.B_shift[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28260_ (.CLK(clk),
    .D(_02058_),
    .Q(\systolic_inst.B_shift[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28261_ (.CLK(clk),
    .D(_02059_),
    .Q(\systolic_inst.B_shift[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28262_ (.CLK(clk),
    .D(_02060_),
    .Q(\systolic_inst.B_shift[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28263_ (.CLK(clk),
    .D(_02061_),
    .Q(\systolic_inst.B_shift[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28264_ (.CLK(clk),
    .D(_02062_),
    .Q(\systolic_inst.B_shift[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28265_ (.CLK(clk),
    .D(_02063_),
    .Q(\systolic_inst.B_shift[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28266_ (.CLK(clk),
    .D(_02064_),
    .Q(\systolic_inst.B_shift[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28267_ (.CLK(clk),
    .D(_02065_),
    .Q(\systolic_inst.B_shift[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28268_ (.CLK(clk),
    .D(_02066_),
    .Q(\systolic_inst.B_shift[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28269_ (.CLK(clk),
    .D(_02067_),
    .Q(\systolic_inst.B_shift[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28270_ (.CLK(clk),
    .D(_02068_),
    .Q(\systolic_inst.B_shift[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28271_ (.CLK(clk),
    .D(_02069_),
    .Q(\systolic_inst.B_shift[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28272_ (.CLK(clk),
    .D(_02070_),
    .Q(\systolic_inst.B_shift[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28273_ (.CLK(clk),
    .D(_02071_),
    .Q(\systolic_inst.B_shift[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28274_ (.CLK(clk),
    .D(_02072_),
    .Q(\systolic_inst.B_shift[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28275_ (.CLK(clk),
    .D(_02073_),
    .Q(\systolic_inst.B_shift[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28276_ (.CLK(clk),
    .D(_02074_),
    .Q(\systolic_inst.B_shift[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28277_ (.CLK(clk),
    .D(_02075_),
    .Q(\systolic_inst.B_shift[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28278_ (.CLK(clk),
    .D(_02076_),
    .Q(\systolic_inst.B_shift[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28279_ (.CLK(clk),
    .D(_02077_),
    .Q(\systolic_inst.B_shift[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28280_ (.CLK(clk),
    .D(_02078_),
    .Q(\systolic_inst.B_shift[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28281_ (.CLK(clk),
    .D(_02079_),
    .Q(\systolic_inst.B_shift[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28282_ (.CLK(clk),
    .D(_02080_),
    .Q(\systolic_inst.B_shift[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28283_ (.CLK(clk),
    .D(_02081_),
    .Q(\systolic_inst.B_shift[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28284_ (.CLK(clk),
    .D(_02082_),
    .Q(\systolic_inst.B_shift[19][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28285_ (.CLK(clk),
    .D(_02083_),
    .Q(\systolic_inst.B_shift[19][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28286_ (.CLK(clk),
    .D(_02084_),
    .Q(\systolic_inst.B_shift[19][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28287_ (.CLK(clk),
    .D(_02085_),
    .Q(\systolic_inst.B_shift[19][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28288_ (.CLK(clk),
    .D(_02086_),
    .Q(\systolic_inst.B_shift[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28289_ (.CLK(clk),
    .D(_02087_),
    .Q(\systolic_inst.B_shift[19][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28290_ (.CLK(clk),
    .D(_02088_),
    .Q(\systolic_inst.B_shift[19][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28291_ (.CLK(clk),
    .D(_02089_),
    .Q(\systolic_inst.B_shift[19][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28292_ (.CLK(clk),
    .D(_02090_),
    .Q(\systolic_inst.B_shift[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28293_ (.CLK(clk),
    .D(_02091_),
    .Q(\systolic_inst.B_shift[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28294_ (.CLK(clk),
    .D(_02092_),
    .Q(\systolic_inst.B_shift[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28295_ (.CLK(clk),
    .D(_02093_),
    .Q(\systolic_inst.B_shift[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28296_ (.CLK(clk),
    .D(_02094_),
    .Q(\systolic_inst.B_shift[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28297_ (.CLK(clk),
    .D(_02095_),
    .Q(\systolic_inst.B_shift[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28298_ (.CLK(clk),
    .D(_02096_),
    .Q(\systolic_inst.B_shift[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28299_ (.CLK(clk),
    .D(_02097_),
    .Q(\systolic_inst.B_shift[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28300_ (.CLK(clk),
    .D(_02098_),
    .Q(\systolic_inst.B_shift[27][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28301_ (.CLK(clk),
    .D(_02099_),
    .Q(\systolic_inst.B_shift[27][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28302_ (.CLK(clk),
    .D(_02100_),
    .Q(\systolic_inst.B_shift[27][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28303_ (.CLK(clk),
    .D(_02101_),
    .Q(\systolic_inst.B_shift[27][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28304_ (.CLK(clk),
    .D(_02102_),
    .Q(\systolic_inst.B_shift[27][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28305_ (.CLK(clk),
    .D(_02103_),
    .Q(\systolic_inst.B_shift[27][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28306_ (.CLK(clk),
    .D(_02104_),
    .Q(\systolic_inst.B_shift[27][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28307_ (.CLK(clk),
    .D(_02105_),
    .Q(\systolic_inst.B_shift[27][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28308_ (.CLK(clk),
    .D(_02106_),
    .Q(\systolic_inst.A_shift[29][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28309_ (.CLK(clk),
    .D(_02107_),
    .Q(\systolic_inst.A_shift[29][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28310_ (.CLK(clk),
    .D(_02108_),
    .Q(\systolic_inst.A_shift[29][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28311_ (.CLK(clk),
    .D(_02109_),
    .Q(\systolic_inst.A_shift[29][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28312_ (.CLK(clk),
    .D(_02110_),
    .Q(\systolic_inst.A_shift[29][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28313_ (.CLK(clk),
    .D(_02111_),
    .Q(\systolic_inst.A_shift[29][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28314_ (.CLK(clk),
    .D(_02112_),
    .Q(\systolic_inst.A_shift[29][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28315_ (.CLK(clk),
    .D(_02113_),
    .Q(\systolic_inst.A_shift[29][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28316_ (.CLK(clk),
    .D(_02114_),
    .Q(\systolic_inst.A_shift[28][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28317_ (.CLK(clk),
    .D(_02115_),
    .Q(\systolic_inst.A_shift[28][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28318_ (.CLK(clk),
    .D(_02116_),
    .Q(\systolic_inst.A_shift[28][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28319_ (.CLK(clk),
    .D(_02117_),
    .Q(\systolic_inst.A_shift[28][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28320_ (.CLK(clk),
    .D(_02118_),
    .Q(\systolic_inst.A_shift[28][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28321_ (.CLK(clk),
    .D(_02119_),
    .Q(\systolic_inst.A_shift[28][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28322_ (.CLK(clk),
    .D(_02120_),
    .Q(\systolic_inst.A_shift[28][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28323_ (.CLK(clk),
    .D(_02121_),
    .Q(\systolic_inst.A_shift[28][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28324_ (.CLK(clk),
    .D(_02122_),
    .Q(\systolic_inst.A_shift[27][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28325_ (.CLK(clk),
    .D(_02123_),
    .Q(\systolic_inst.A_shift[27][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28326_ (.CLK(clk),
    .D(_02124_),
    .Q(\systolic_inst.A_shift[27][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28327_ (.CLK(clk),
    .D(_02125_),
    .Q(\systolic_inst.A_shift[27][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28328_ (.CLK(clk),
    .D(_02126_),
    .Q(\systolic_inst.A_shift[27][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28329_ (.CLK(clk),
    .D(_02127_),
    .Q(\systolic_inst.A_shift[27][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28330_ (.CLK(clk),
    .D(_02128_),
    .Q(\systolic_inst.A_shift[27][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28331_ (.CLK(clk),
    .D(_02129_),
    .Q(\systolic_inst.A_shift[27][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28332_ (.CLK(clk),
    .D(_02130_),
    .Q(\systolic_inst.A_shift[26][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28333_ (.CLK(clk),
    .D(_02131_),
    .Q(\systolic_inst.A_shift[26][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28334_ (.CLK(clk),
    .D(_02132_),
    .Q(\systolic_inst.A_shift[26][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28335_ (.CLK(clk),
    .D(_02133_),
    .Q(\systolic_inst.A_shift[26][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28336_ (.CLK(clk),
    .D(_02134_),
    .Q(\systolic_inst.A_shift[26][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28337_ (.CLK(clk),
    .D(_02135_),
    .Q(\systolic_inst.A_shift[26][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28338_ (.CLK(clk),
    .D(_02136_),
    .Q(\systolic_inst.A_shift[26][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28339_ (.CLK(clk),
    .D(_02137_),
    .Q(\systolic_inst.A_shift[26][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28340_ (.CLK(clk),
    .D(_02138_),
    .Q(\systolic_inst.A_shift[25][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28341_ (.CLK(clk),
    .D(_02139_),
    .Q(\systolic_inst.A_shift[25][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28342_ (.CLK(clk),
    .D(_02140_),
    .Q(\systolic_inst.A_shift[25][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28343_ (.CLK(clk),
    .D(_02141_),
    .Q(\systolic_inst.A_shift[25][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28344_ (.CLK(clk),
    .D(_02142_),
    .Q(\systolic_inst.A_shift[25][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28345_ (.CLK(clk),
    .D(_02143_),
    .Q(\systolic_inst.A_shift[25][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28346_ (.CLK(clk),
    .D(_02144_),
    .Q(\systolic_inst.A_shift[25][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28347_ (.CLK(clk),
    .D(_02145_),
    .Q(\systolic_inst.A_shift[25][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28348_ (.CLK(clk),
    .D(_02146_),
    .Q(\systolic_inst.A_shift[24][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28349_ (.CLK(clk),
    .D(_02147_),
    .Q(\systolic_inst.A_shift[24][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28350_ (.CLK(clk),
    .D(_02148_),
    .Q(\systolic_inst.A_shift[24][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28351_ (.CLK(clk),
    .D(_02149_),
    .Q(\systolic_inst.A_shift[24][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28352_ (.CLK(clk),
    .D(_02150_),
    .Q(\systolic_inst.A_shift[24][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28353_ (.CLK(clk),
    .D(_02151_),
    .Q(\systolic_inst.A_shift[24][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28354_ (.CLK(clk),
    .D(_02152_),
    .Q(\systolic_inst.A_shift[24][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28355_ (.CLK(clk),
    .D(_02153_),
    .Q(\systolic_inst.A_shift[24][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28356_ (.CLK(clk),
    .D(_02154_),
    .Q(\systolic_inst.B_shift[22][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28357_ (.CLK(clk),
    .D(_02155_),
    .Q(\systolic_inst.B_shift[22][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28358_ (.CLK(clk),
    .D(_02156_),
    .Q(\systolic_inst.B_shift[22][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28359_ (.CLK(clk),
    .D(_02157_),
    .Q(\systolic_inst.B_shift[22][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28360_ (.CLK(clk),
    .D(_02158_),
    .Q(\systolic_inst.B_shift[22][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28361_ (.CLK(clk),
    .D(_02159_),
    .Q(\systolic_inst.B_shift[22][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28362_ (.CLK(clk),
    .D(_02160_),
    .Q(\systolic_inst.B_shift[22][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28363_ (.CLK(clk),
    .D(_02161_),
    .Q(\systolic_inst.B_shift[22][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28364_ (.CLK(clk),
    .D(_02162_),
    .Q(\systolic_inst.A_shift[20][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28365_ (.CLK(clk),
    .D(_02163_),
    .Q(\systolic_inst.A_shift[20][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28366_ (.CLK(clk),
    .D(_02164_),
    .Q(\systolic_inst.A_shift[20][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28367_ (.CLK(clk),
    .D(_02165_),
    .Q(\systolic_inst.A_shift[20][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28368_ (.CLK(clk),
    .D(_02166_),
    .Q(\systolic_inst.A_shift[20][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28369_ (.CLK(clk),
    .D(_02167_),
    .Q(\systolic_inst.A_shift[20][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28370_ (.CLK(clk),
    .D(_02168_),
    .Q(\systolic_inst.A_shift[20][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28371_ (.CLK(clk),
    .D(_02169_),
    .Q(\systolic_inst.A_shift[20][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28372_ (.CLK(clk),
    .D(_02170_),
    .Q(\systolic_inst.A_shift[19][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28373_ (.CLK(clk),
    .D(_02171_),
    .Q(\systolic_inst.A_shift[19][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28374_ (.CLK(clk),
    .D(_02172_),
    .Q(\systolic_inst.A_shift[19][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28375_ (.CLK(clk),
    .D(_02173_),
    .Q(\systolic_inst.A_shift[19][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28376_ (.CLK(clk),
    .D(_02174_),
    .Q(\systolic_inst.A_shift[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28377_ (.CLK(clk),
    .D(_02175_),
    .Q(\systolic_inst.A_shift[19][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28378_ (.CLK(clk),
    .D(_02176_),
    .Q(\systolic_inst.A_shift[19][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28379_ (.CLK(clk),
    .D(_02177_),
    .Q(\systolic_inst.A_shift[19][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28380_ (.CLK(clk),
    .D(_02178_),
    .Q(\systolic_inst.A_shift[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28381_ (.CLK(clk),
    .D(_02179_),
    .Q(\systolic_inst.A_shift[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28382_ (.CLK(clk),
    .D(_02180_),
    .Q(\systolic_inst.A_shift[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28383_ (.CLK(clk),
    .D(_02181_),
    .Q(\systolic_inst.A_shift[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28384_ (.CLK(clk),
    .D(_02182_),
    .Q(\systolic_inst.A_shift[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28385_ (.CLK(clk),
    .D(_02183_),
    .Q(\systolic_inst.A_shift[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28386_ (.CLK(clk),
    .D(_02184_),
    .Q(\systolic_inst.A_shift[18][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28387_ (.CLK(clk),
    .D(_02185_),
    .Q(\systolic_inst.A_shift[18][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28388_ (.CLK(clk),
    .D(_02186_),
    .Q(\systolic_inst.A_shift[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28389_ (.CLK(clk),
    .D(_02187_),
    .Q(\systolic_inst.A_shift[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28390_ (.CLK(clk),
    .D(_02188_),
    .Q(\systolic_inst.A_shift[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28391_ (.CLK(clk),
    .D(_02189_),
    .Q(\systolic_inst.A_shift[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28392_ (.CLK(clk),
    .D(_02190_),
    .Q(\systolic_inst.A_shift[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28393_ (.CLK(clk),
    .D(_02191_),
    .Q(\systolic_inst.A_shift[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28394_ (.CLK(clk),
    .D(_02192_),
    .Q(\systolic_inst.A_shift[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28395_ (.CLK(clk),
    .D(_02193_),
    .Q(\systolic_inst.A_shift[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28396_ (.CLK(clk),
    .D(_02194_),
    .Q(\systolic_inst.A_shift[16][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28397_ (.CLK(clk),
    .D(_02195_),
    .Q(\systolic_inst.A_shift[16][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28398_ (.CLK(clk),
    .D(_02196_),
    .Q(\systolic_inst.A_shift[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28399_ (.CLK(clk),
    .D(_02197_),
    .Q(\systolic_inst.A_shift[16][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28400_ (.CLK(clk),
    .D(_02198_),
    .Q(\systolic_inst.A_shift[16][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28401_ (.CLK(clk),
    .D(_02199_),
    .Q(\systolic_inst.A_shift[16][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28402_ (.CLK(clk),
    .D(_02200_),
    .Q(\systolic_inst.A_shift[16][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28403_ (.CLK(clk),
    .D(_02201_),
    .Q(\systolic_inst.A_shift[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28404_ (.CLK(clk),
    .D(_02202_),
    .Q(\systolic_inst.B_shift[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28405_ (.CLK(clk),
    .D(_02203_),
    .Q(\systolic_inst.B_shift[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28406_ (.CLK(clk),
    .D(_02204_),
    .Q(\systolic_inst.B_shift[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28407_ (.CLK(clk),
    .D(_02205_),
    .Q(\systolic_inst.B_shift[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28408_ (.CLK(clk),
    .D(_02206_),
    .Q(\systolic_inst.B_shift[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28409_ (.CLK(clk),
    .D(_02207_),
    .Q(\systolic_inst.B_shift[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28410_ (.CLK(clk),
    .D(_02208_),
    .Q(\systolic_inst.B_shift[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28411_ (.CLK(clk),
    .D(_02209_),
    .Q(\systolic_inst.B_shift[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28412_ (.CLK(clk),
    .D(_02210_),
    .Q(\systolic_inst.B_shift[23][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28413_ (.CLK(clk),
    .D(_02211_),
    .Q(\systolic_inst.B_shift[23][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28414_ (.CLK(clk),
    .D(_02212_),
    .Q(\systolic_inst.B_shift[23][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28415_ (.CLK(clk),
    .D(_02213_),
    .Q(\systolic_inst.B_shift[23][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28416_ (.CLK(clk),
    .D(_02214_),
    .Q(\systolic_inst.B_shift[23][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28417_ (.CLK(clk),
    .D(_02215_),
    .Q(\systolic_inst.B_shift[23][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28418_ (.CLK(clk),
    .D(_02216_),
    .Q(\systolic_inst.B_shift[23][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28419_ (.CLK(clk),
    .D(_02217_),
    .Q(\systolic_inst.B_shift[23][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28420_ (.CLK(clk),
    .D(_02218_),
    .Q(\systolic_inst.A_shift[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28421_ (.CLK(clk),
    .D(_02219_),
    .Q(\systolic_inst.A_shift[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28422_ (.CLK(clk),
    .D(_02220_),
    .Q(\systolic_inst.A_shift[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28423_ (.CLK(clk),
    .D(_02221_),
    .Q(\systolic_inst.A_shift[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28424_ (.CLK(clk),
    .D(_02222_),
    .Q(\systolic_inst.A_shift[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28425_ (.CLK(clk),
    .D(_02223_),
    .Q(\systolic_inst.A_shift[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28426_ (.CLK(clk),
    .D(_02224_),
    .Q(\systolic_inst.A_shift[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28427_ (.CLK(clk),
    .D(_02225_),
    .Q(\systolic_inst.A_shift[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28428_ (.CLK(clk),
    .D(_02226_),
    .Q(\systolic_inst.A_shift[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28429_ (.CLK(clk),
    .D(_02227_),
    .Q(\systolic_inst.A_shift[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28430_ (.CLK(clk),
    .D(_02228_),
    .Q(\systolic_inst.A_shift[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28431_ (.CLK(clk),
    .D(_02229_),
    .Q(\systolic_inst.A_shift[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28432_ (.CLK(clk),
    .D(_02230_),
    .Q(\systolic_inst.A_shift[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28433_ (.CLK(clk),
    .D(_02231_),
    .Q(\systolic_inst.A_shift[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28434_ (.CLK(clk),
    .D(_02232_),
    .Q(\systolic_inst.A_shift[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28435_ (.CLK(clk),
    .D(_02233_),
    .Q(\systolic_inst.A_shift[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28436_ (.CLK(clk),
    .D(_02234_),
    .Q(\systolic_inst.A_shift[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28437_ (.CLK(clk),
    .D(_02235_),
    .Q(\systolic_inst.A_shift[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28438_ (.CLK(clk),
    .D(_02236_),
    .Q(\systolic_inst.A_shift[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28439_ (.CLK(clk),
    .D(_02237_),
    .Q(\systolic_inst.A_shift[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28440_ (.CLK(clk),
    .D(_02238_),
    .Q(\systolic_inst.A_shift[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28441_ (.CLK(clk),
    .D(_02239_),
    .Q(\systolic_inst.A_shift[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28442_ (.CLK(clk),
    .D(_02240_),
    .Q(\systolic_inst.A_shift[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28443_ (.CLK(clk),
    .D(_02241_),
    .Q(\systolic_inst.A_shift[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28444_ (.CLK(clk),
    .D(_02242_),
    .Q(\systolic_inst.A_shift[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28445_ (.CLK(clk),
    .D(_02243_),
    .Q(\systolic_inst.A_shift[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28446_ (.CLK(clk),
    .D(_02244_),
    .Q(\systolic_inst.A_shift[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28447_ (.CLK(clk),
    .D(_02245_),
    .Q(\systolic_inst.A_shift[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28448_ (.CLK(clk),
    .D(_02246_),
    .Q(\systolic_inst.A_shift[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28449_ (.CLK(clk),
    .D(_02247_),
    .Q(\systolic_inst.A_shift[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28450_ (.CLK(clk),
    .D(_02248_),
    .Q(\systolic_inst.A_shift[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28451_ (.CLK(clk),
    .D(_02249_),
    .Q(\systolic_inst.A_shift[8][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28452_ (.CLK(clk),
    .D(_02250_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _28453_ (.CLK(clk),
    .D(_02251_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _28454_ (.CLK(clk),
    .D(_02252_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _28455_ (.CLK(clk),
    .D(_02253_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 _28456_ (.CLK(clk),
    .D(_02254_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_2 _28457_ (.CLK(clk),
    .D(_02255_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _28458_ (.CLK(clk),
    .D(_02256_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_2 _28459_ (.CLK(clk),
    .D(_02257_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[7] ));
 sky130_fd_sc_hd__dfrtp_2 _28460_ (.CLK(clk),
    .D(_02258_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[8] ));
 sky130_fd_sc_hd__dfrtp_2 _28461_ (.CLK(clk),
    .D(_02259_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[9] ));
 sky130_fd_sc_hd__dfrtp_2 _28462_ (.CLK(clk),
    .D(_02260_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[10] ));
 sky130_fd_sc_hd__dfrtp_2 _28463_ (.CLK(clk),
    .D(_02261_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[11] ));
 sky130_fd_sc_hd__dfrtp_2 _28464_ (.CLK(clk),
    .D(_02262_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[12] ));
 sky130_fd_sc_hd__dfrtp_2 _28465_ (.CLK(clk),
    .D(_02263_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[13] ));
 sky130_fd_sc_hd__dfrtp_2 _28466_ (.CLK(clk),
    .D(_02264_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[14] ));
 sky130_fd_sc_hd__dfrtp_2 _28467_ (.CLK(clk),
    .D(_02265_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[15] ));
 sky130_fd_sc_hd__dfrtp_2 _28468_ (.CLK(clk),
    .D(_02266_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[16] ));
 sky130_fd_sc_hd__dfrtp_2 _28469_ (.CLK(clk),
    .D(_02267_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[17] ));
 sky130_fd_sc_hd__dfrtp_2 _28470_ (.CLK(clk),
    .D(_02268_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[18] ));
 sky130_fd_sc_hd__dfrtp_2 _28471_ (.CLK(clk),
    .D(_02269_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[19] ));
 sky130_fd_sc_hd__dfrtp_2 _28472_ (.CLK(clk),
    .D(_02270_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[20] ));
 sky130_fd_sc_hd__dfrtp_2 _28473_ (.CLK(clk),
    .D(_02271_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[21] ));
 sky130_fd_sc_hd__dfrtp_2 _28474_ (.CLK(clk),
    .D(_02272_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[22] ));
 sky130_fd_sc_hd__dfrtp_2 _28475_ (.CLK(clk),
    .D(_02273_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[23] ));
 sky130_fd_sc_hd__dfrtp_2 _28476_ (.CLK(clk),
    .D(_02274_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[24] ));
 sky130_fd_sc_hd__dfrtp_2 _28477_ (.CLK(clk),
    .D(_02275_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[25] ));
 sky130_fd_sc_hd__dfrtp_2 _28478_ (.CLK(clk),
    .D(_02276_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[26] ));
 sky130_fd_sc_hd__dfrtp_2 _28479_ (.CLK(clk),
    .D(_02277_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[27] ));
 sky130_fd_sc_hd__dfrtp_2 _28480_ (.CLK(clk),
    .D(_02278_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[28] ));
 sky130_fd_sc_hd__dfrtp_2 _28481_ (.CLK(clk),
    .D(_02279_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[29] ));
 sky130_fd_sc_hd__dfrtp_2 _28482_ (.CLK(clk),
    .D(_02280_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[30] ));
 sky130_fd_sc_hd__dfrtp_2 _28483_ (.CLK(clk),
    .D(_02281_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[31] ));
 sky130_fd_sc_hd__dfrtp_2 _28484_ (.CLK(clk),
    .D(_02282_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[32] ));
 sky130_fd_sc_hd__dfrtp_2 _28485_ (.CLK(clk),
    .D(_02283_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[33] ));
 sky130_fd_sc_hd__dfrtp_2 _28486_ (.CLK(clk),
    .D(_02284_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[34] ));
 sky130_fd_sc_hd__dfrtp_2 _28487_ (.CLK(clk),
    .D(_02285_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[35] ));
 sky130_fd_sc_hd__dfrtp_2 _28488_ (.CLK(clk),
    .D(_02286_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[36] ));
 sky130_fd_sc_hd__dfrtp_2 _28489_ (.CLK(clk),
    .D(_02287_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[37] ));
 sky130_fd_sc_hd__dfrtp_2 _28490_ (.CLK(clk),
    .D(_02288_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[38] ));
 sky130_fd_sc_hd__dfrtp_2 _28491_ (.CLK(clk),
    .D(_02289_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[39] ));
 sky130_fd_sc_hd__dfrtp_2 _28492_ (.CLK(clk),
    .D(_02290_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[40] ));
 sky130_fd_sc_hd__dfrtp_2 _28493_ (.CLK(clk),
    .D(_02291_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[41] ));
 sky130_fd_sc_hd__dfrtp_2 _28494_ (.CLK(clk),
    .D(_02292_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[42] ));
 sky130_fd_sc_hd__dfrtp_2 _28495_ (.CLK(clk),
    .D(_02293_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[43] ));
 sky130_fd_sc_hd__dfrtp_2 _28496_ (.CLK(clk),
    .D(_02294_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[44] ));
 sky130_fd_sc_hd__dfrtp_2 _28497_ (.CLK(clk),
    .D(_02295_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[45] ));
 sky130_fd_sc_hd__dfrtp_2 _28498_ (.CLK(clk),
    .D(_02296_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[46] ));
 sky130_fd_sc_hd__dfrtp_2 _28499_ (.CLK(clk),
    .D(_02297_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[47] ));
 sky130_fd_sc_hd__dfrtp_2 _28500_ (.CLK(clk),
    .D(_02298_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[48] ));
 sky130_fd_sc_hd__dfrtp_2 _28501_ (.CLK(clk),
    .D(_02299_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[49] ));
 sky130_fd_sc_hd__dfrtp_2 _28502_ (.CLK(clk),
    .D(_02300_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[50] ));
 sky130_fd_sc_hd__dfrtp_2 _28503_ (.CLK(clk),
    .D(_02301_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[51] ));
 sky130_fd_sc_hd__dfrtp_2 _28504_ (.CLK(clk),
    .D(_02302_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[52] ));
 sky130_fd_sc_hd__dfrtp_2 _28505_ (.CLK(clk),
    .D(_02303_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[53] ));
 sky130_fd_sc_hd__dfrtp_2 _28506_ (.CLK(clk),
    .D(_02304_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[54] ));
 sky130_fd_sc_hd__dfrtp_2 _28507_ (.CLK(clk),
    .D(_02305_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[55] ));
 sky130_fd_sc_hd__dfrtp_2 _28508_ (.CLK(clk),
    .D(_02306_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[56] ));
 sky130_fd_sc_hd__dfrtp_2 _28509_ (.CLK(clk),
    .D(_02307_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[57] ));
 sky130_fd_sc_hd__dfrtp_2 _28510_ (.CLK(clk),
    .D(_02308_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[58] ));
 sky130_fd_sc_hd__dfrtp_2 _28511_ (.CLK(clk),
    .D(_02309_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[59] ));
 sky130_fd_sc_hd__dfrtp_2 _28512_ (.CLK(clk),
    .D(_02310_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[60] ));
 sky130_fd_sc_hd__dfrtp_2 _28513_ (.CLK(clk),
    .D(_02311_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[61] ));
 sky130_fd_sc_hd__dfrtp_2 _28514_ (.CLK(clk),
    .D(_02312_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[62] ));
 sky130_fd_sc_hd__dfrtp_2 _28515_ (.CLK(clk),
    .D(_02313_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[63] ));
 sky130_fd_sc_hd__dfrtp_2 _28516_ (.CLK(clk),
    .D(_02314_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[64] ));
 sky130_fd_sc_hd__dfrtp_2 _28517_ (.CLK(clk),
    .D(_02315_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[65] ));
 sky130_fd_sc_hd__dfrtp_2 _28518_ (.CLK(clk),
    .D(_02316_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[66] ));
 sky130_fd_sc_hd__dfrtp_2 _28519_ (.CLK(clk),
    .D(_02317_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[67] ));
 sky130_fd_sc_hd__dfrtp_2 _28520_ (.CLK(clk),
    .D(_02318_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[68] ));
 sky130_fd_sc_hd__dfrtp_2 _28521_ (.CLK(clk),
    .D(_02319_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[69] ));
 sky130_fd_sc_hd__dfrtp_2 _28522_ (.CLK(clk),
    .D(_02320_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[70] ));
 sky130_fd_sc_hd__dfrtp_2 _28523_ (.CLK(clk),
    .D(_02321_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[71] ));
 sky130_fd_sc_hd__dfrtp_2 _28524_ (.CLK(clk),
    .D(_02322_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[72] ));
 sky130_fd_sc_hd__dfrtp_2 _28525_ (.CLK(clk),
    .D(_02323_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[73] ));
 sky130_fd_sc_hd__dfrtp_2 _28526_ (.CLK(clk),
    .D(_02324_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[74] ));
 sky130_fd_sc_hd__dfrtp_2 _28527_ (.CLK(clk),
    .D(_02325_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[75] ));
 sky130_fd_sc_hd__dfrtp_2 _28528_ (.CLK(clk),
    .D(_02326_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[76] ));
 sky130_fd_sc_hd__dfrtp_2 _28529_ (.CLK(clk),
    .D(_02327_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[77] ));
 sky130_fd_sc_hd__dfrtp_2 _28530_ (.CLK(clk),
    .D(_02328_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[78] ));
 sky130_fd_sc_hd__dfrtp_2 _28531_ (.CLK(clk),
    .D(_02329_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[79] ));
 sky130_fd_sc_hd__dfrtp_2 _28532_ (.CLK(clk),
    .D(_02330_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[80] ));
 sky130_fd_sc_hd__dfrtp_2 _28533_ (.CLK(clk),
    .D(_02331_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[81] ));
 sky130_fd_sc_hd__dfrtp_2 _28534_ (.CLK(clk),
    .D(_02332_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[82] ));
 sky130_fd_sc_hd__dfrtp_2 _28535_ (.CLK(clk),
    .D(_02333_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[83] ));
 sky130_fd_sc_hd__dfrtp_2 _28536_ (.CLK(clk),
    .D(_02334_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[84] ));
 sky130_fd_sc_hd__dfrtp_2 _28537_ (.CLK(clk),
    .D(_02335_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[85] ));
 sky130_fd_sc_hd__dfrtp_2 _28538_ (.CLK(clk),
    .D(_02336_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[86] ));
 sky130_fd_sc_hd__dfrtp_2 _28539_ (.CLK(clk),
    .D(_02337_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[87] ));
 sky130_fd_sc_hd__dfrtp_2 _28540_ (.CLK(clk),
    .D(_02338_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[88] ));
 sky130_fd_sc_hd__dfrtp_2 _28541_ (.CLK(clk),
    .D(_02339_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[89] ));
 sky130_fd_sc_hd__dfrtp_2 _28542_ (.CLK(clk),
    .D(_02340_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[90] ));
 sky130_fd_sc_hd__dfrtp_2 _28543_ (.CLK(clk),
    .D(_02341_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[91] ));
 sky130_fd_sc_hd__dfrtp_2 _28544_ (.CLK(clk),
    .D(_02342_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[92] ));
 sky130_fd_sc_hd__dfrtp_2 _28545_ (.CLK(clk),
    .D(_02343_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[93] ));
 sky130_fd_sc_hd__dfrtp_2 _28546_ (.CLK(clk),
    .D(_02344_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[94] ));
 sky130_fd_sc_hd__dfrtp_2 _28547_ (.CLK(clk),
    .D(_02345_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[95] ));
 sky130_fd_sc_hd__dfrtp_2 _28548_ (.CLK(clk),
    .D(_02346_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[96] ));
 sky130_fd_sc_hd__dfrtp_2 _28549_ (.CLK(clk),
    .D(_02347_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[97] ));
 sky130_fd_sc_hd__dfrtp_2 _28550_ (.CLK(clk),
    .D(_02348_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[98] ));
 sky130_fd_sc_hd__dfrtp_2 _28551_ (.CLK(clk),
    .D(_02349_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[99] ));
 sky130_fd_sc_hd__dfrtp_2 _28552_ (.CLK(clk),
    .D(_02350_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[100] ));
 sky130_fd_sc_hd__dfrtp_2 _28553_ (.CLK(clk),
    .D(_02351_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[101] ));
 sky130_fd_sc_hd__dfrtp_2 _28554_ (.CLK(clk),
    .D(_02352_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[102] ));
 sky130_fd_sc_hd__dfrtp_2 _28555_ (.CLK(clk),
    .D(_02353_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[103] ));
 sky130_fd_sc_hd__dfrtp_2 _28556_ (.CLK(clk),
    .D(_02354_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[104] ));
 sky130_fd_sc_hd__dfrtp_2 _28557_ (.CLK(clk),
    .D(_02355_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[105] ));
 sky130_fd_sc_hd__dfrtp_2 _28558_ (.CLK(clk),
    .D(_02356_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[106] ));
 sky130_fd_sc_hd__dfrtp_2 _28559_ (.CLK(clk),
    .D(_02357_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[107] ));
 sky130_fd_sc_hd__dfrtp_2 _28560_ (.CLK(clk),
    .D(_02358_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[108] ));
 sky130_fd_sc_hd__dfrtp_2 _28561_ (.CLK(clk),
    .D(_02359_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[109] ));
 sky130_fd_sc_hd__dfrtp_2 _28562_ (.CLK(clk),
    .D(_02360_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[110] ));
 sky130_fd_sc_hd__dfrtp_2 _28563_ (.CLK(clk),
    .D(_02361_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[111] ));
 sky130_fd_sc_hd__dfrtp_2 _28564_ (.CLK(clk),
    .D(_02362_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[112] ));
 sky130_fd_sc_hd__dfrtp_2 _28565_ (.CLK(clk),
    .D(_02363_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[113] ));
 sky130_fd_sc_hd__dfrtp_2 _28566_ (.CLK(clk),
    .D(_02364_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[114] ));
 sky130_fd_sc_hd__dfrtp_2 _28567_ (.CLK(clk),
    .D(_02365_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[115] ));
 sky130_fd_sc_hd__dfrtp_2 _28568_ (.CLK(clk),
    .D(_02366_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[116] ));
 sky130_fd_sc_hd__dfrtp_2 _28569_ (.CLK(clk),
    .D(_02367_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[117] ));
 sky130_fd_sc_hd__dfrtp_2 _28570_ (.CLK(clk),
    .D(_02368_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[118] ));
 sky130_fd_sc_hd__dfrtp_2 _28571_ (.CLK(clk),
    .D(_02369_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[119] ));
 sky130_fd_sc_hd__dfrtp_2 _28572_ (.CLK(clk),
    .D(_02370_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[120] ));
 sky130_fd_sc_hd__dfrtp_2 _28573_ (.CLK(clk),
    .D(_02371_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[121] ));
 sky130_fd_sc_hd__dfrtp_2 _28574_ (.CLK(clk),
    .D(_02372_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[122] ));
 sky130_fd_sc_hd__dfrtp_2 _28575_ (.CLK(clk),
    .D(_02373_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[123] ));
 sky130_fd_sc_hd__dfrtp_2 _28576_ (.CLK(clk),
    .D(_02374_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[124] ));
 sky130_fd_sc_hd__dfrtp_2 _28577_ (.CLK(clk),
    .D(_02375_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[125] ));
 sky130_fd_sc_hd__dfrtp_2 _28578_ (.CLK(clk),
    .D(_02376_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[126] ));
 sky130_fd_sc_hd__dfrtp_2 _28579_ (.CLK(clk),
    .D(_02377_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[127] ));
 sky130_fd_sc_hd__dfrtp_2 _28580_ (.CLK(clk),
    .D(_02378_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[128] ));
 sky130_fd_sc_hd__dfrtp_2 _28581_ (.CLK(clk),
    .D(_02379_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[129] ));
 sky130_fd_sc_hd__dfrtp_2 _28582_ (.CLK(clk),
    .D(_02380_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[130] ));
 sky130_fd_sc_hd__dfrtp_2 _28583_ (.CLK(clk),
    .D(_02381_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[131] ));
 sky130_fd_sc_hd__dfrtp_2 _28584_ (.CLK(clk),
    .D(_02382_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[132] ));
 sky130_fd_sc_hd__dfrtp_2 _28585_ (.CLK(clk),
    .D(_02383_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[133] ));
 sky130_fd_sc_hd__dfrtp_2 _28586_ (.CLK(clk),
    .D(_02384_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[134] ));
 sky130_fd_sc_hd__dfrtp_2 _28587_ (.CLK(clk),
    .D(_02385_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[135] ));
 sky130_fd_sc_hd__dfrtp_2 _28588_ (.CLK(clk),
    .D(_02386_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[136] ));
 sky130_fd_sc_hd__dfrtp_2 _28589_ (.CLK(clk),
    .D(_02387_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[137] ));
 sky130_fd_sc_hd__dfrtp_2 _28590_ (.CLK(clk),
    .D(_02388_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[138] ));
 sky130_fd_sc_hd__dfrtp_2 _28591_ (.CLK(clk),
    .D(_02389_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[139] ));
 sky130_fd_sc_hd__dfrtp_2 _28592_ (.CLK(clk),
    .D(_02390_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[140] ));
 sky130_fd_sc_hd__dfrtp_2 _28593_ (.CLK(clk),
    .D(_02391_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[141] ));
 sky130_fd_sc_hd__dfrtp_2 _28594_ (.CLK(clk),
    .D(_02392_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[142] ));
 sky130_fd_sc_hd__dfrtp_2 _28595_ (.CLK(clk),
    .D(_02393_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[143] ));
 sky130_fd_sc_hd__dfrtp_2 _28596_ (.CLK(clk),
    .D(_02394_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[144] ));
 sky130_fd_sc_hd__dfrtp_2 _28597_ (.CLK(clk),
    .D(_02395_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[145] ));
 sky130_fd_sc_hd__dfrtp_2 _28598_ (.CLK(clk),
    .D(_02396_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[146] ));
 sky130_fd_sc_hd__dfrtp_2 _28599_ (.CLK(clk),
    .D(_02397_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[147] ));
 sky130_fd_sc_hd__dfrtp_2 _28600_ (.CLK(clk),
    .D(_02398_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[148] ));
 sky130_fd_sc_hd__dfrtp_2 _28601_ (.CLK(clk),
    .D(_02399_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[149] ));
 sky130_fd_sc_hd__dfrtp_2 _28602_ (.CLK(clk),
    .D(_02400_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[150] ));
 sky130_fd_sc_hd__dfrtp_2 _28603_ (.CLK(clk),
    .D(_02401_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[151] ));
 sky130_fd_sc_hd__dfrtp_2 _28604_ (.CLK(clk),
    .D(_02402_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[152] ));
 sky130_fd_sc_hd__dfrtp_2 _28605_ (.CLK(clk),
    .D(_02403_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[153] ));
 sky130_fd_sc_hd__dfrtp_2 _28606_ (.CLK(clk),
    .D(_02404_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[154] ));
 sky130_fd_sc_hd__dfrtp_2 _28607_ (.CLK(clk),
    .D(_02405_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[155] ));
 sky130_fd_sc_hd__dfrtp_2 _28608_ (.CLK(clk),
    .D(_02406_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[156] ));
 sky130_fd_sc_hd__dfrtp_2 _28609_ (.CLK(clk),
    .D(_02407_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[157] ));
 sky130_fd_sc_hd__dfrtp_2 _28610_ (.CLK(clk),
    .D(_02408_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[158] ));
 sky130_fd_sc_hd__dfrtp_2 _28611_ (.CLK(clk),
    .D(_02409_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[159] ));
 sky130_fd_sc_hd__dfrtp_2 _28612_ (.CLK(clk),
    .D(_02410_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[160] ));
 sky130_fd_sc_hd__dfrtp_2 _28613_ (.CLK(clk),
    .D(_02411_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[161] ));
 sky130_fd_sc_hd__dfrtp_2 _28614_ (.CLK(clk),
    .D(_02412_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[162] ));
 sky130_fd_sc_hd__dfrtp_2 _28615_ (.CLK(clk),
    .D(_02413_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[163] ));
 sky130_fd_sc_hd__dfrtp_2 _28616_ (.CLK(clk),
    .D(_02414_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[164] ));
 sky130_fd_sc_hd__dfrtp_2 _28617_ (.CLK(clk),
    .D(_02415_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[165] ));
 sky130_fd_sc_hd__dfrtp_2 _28618_ (.CLK(clk),
    .D(_02416_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[166] ));
 sky130_fd_sc_hd__dfrtp_2 _28619_ (.CLK(clk),
    .D(_02417_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[167] ));
 sky130_fd_sc_hd__dfrtp_2 _28620_ (.CLK(clk),
    .D(_02418_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[168] ));
 sky130_fd_sc_hd__dfrtp_2 _28621_ (.CLK(clk),
    .D(_02419_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[169] ));
 sky130_fd_sc_hd__dfrtp_2 _28622_ (.CLK(clk),
    .D(_02420_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[170] ));
 sky130_fd_sc_hd__dfrtp_2 _28623_ (.CLK(clk),
    .D(_02421_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[171] ));
 sky130_fd_sc_hd__dfrtp_2 _28624_ (.CLK(clk),
    .D(_02422_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[172] ));
 sky130_fd_sc_hd__dfrtp_2 _28625_ (.CLK(clk),
    .D(_02423_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[173] ));
 sky130_fd_sc_hd__dfrtp_2 _28626_ (.CLK(clk),
    .D(_02424_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[174] ));
 sky130_fd_sc_hd__dfrtp_2 _28627_ (.CLK(clk),
    .D(_02425_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[175] ));
 sky130_fd_sc_hd__dfrtp_2 _28628_ (.CLK(clk),
    .D(_02426_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[176] ));
 sky130_fd_sc_hd__dfrtp_2 _28629_ (.CLK(clk),
    .D(_02427_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[177] ));
 sky130_fd_sc_hd__dfrtp_2 _28630_ (.CLK(clk),
    .D(_02428_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[178] ));
 sky130_fd_sc_hd__dfrtp_2 _28631_ (.CLK(clk),
    .D(_02429_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[179] ));
 sky130_fd_sc_hd__dfrtp_2 _28632_ (.CLK(clk),
    .D(_02430_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[180] ));
 sky130_fd_sc_hd__dfrtp_2 _28633_ (.CLK(clk),
    .D(_02431_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[181] ));
 sky130_fd_sc_hd__dfrtp_2 _28634_ (.CLK(clk),
    .D(_02432_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[182] ));
 sky130_fd_sc_hd__dfrtp_2 _28635_ (.CLK(clk),
    .D(_02433_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[183] ));
 sky130_fd_sc_hd__dfrtp_2 _28636_ (.CLK(clk),
    .D(_02434_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[184] ));
 sky130_fd_sc_hd__dfrtp_2 _28637_ (.CLK(clk),
    .D(_02435_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[185] ));
 sky130_fd_sc_hd__dfrtp_2 _28638_ (.CLK(clk),
    .D(_02436_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[186] ));
 sky130_fd_sc_hd__dfrtp_2 _28639_ (.CLK(clk),
    .D(_02437_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[187] ));
 sky130_fd_sc_hd__dfrtp_2 _28640_ (.CLK(clk),
    .D(_02438_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[188] ));
 sky130_fd_sc_hd__dfrtp_2 _28641_ (.CLK(clk),
    .D(_02439_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[189] ));
 sky130_fd_sc_hd__dfrtp_2 _28642_ (.CLK(clk),
    .D(_02440_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[190] ));
 sky130_fd_sc_hd__dfrtp_2 _28643_ (.CLK(clk),
    .D(_02441_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[191] ));
 sky130_fd_sc_hd__dfrtp_2 _28644_ (.CLK(clk),
    .D(_02442_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[192] ));
 sky130_fd_sc_hd__dfrtp_2 _28645_ (.CLK(clk),
    .D(_02443_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[193] ));
 sky130_fd_sc_hd__dfrtp_2 _28646_ (.CLK(clk),
    .D(_02444_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[194] ));
 sky130_fd_sc_hd__dfrtp_2 _28647_ (.CLK(clk),
    .D(_02445_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[195] ));
 sky130_fd_sc_hd__dfrtp_2 _28648_ (.CLK(clk),
    .D(_02446_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[196] ));
 sky130_fd_sc_hd__dfrtp_2 _28649_ (.CLK(clk),
    .D(_02447_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[197] ));
 sky130_fd_sc_hd__dfrtp_2 _28650_ (.CLK(clk),
    .D(_02448_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[198] ));
 sky130_fd_sc_hd__dfrtp_2 _28651_ (.CLK(clk),
    .D(_02449_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[199] ));
 sky130_fd_sc_hd__dfrtp_2 _28652_ (.CLK(clk),
    .D(_02450_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[200] ));
 sky130_fd_sc_hd__dfrtp_2 _28653_ (.CLK(clk),
    .D(_02451_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[201] ));
 sky130_fd_sc_hd__dfrtp_2 _28654_ (.CLK(clk),
    .D(_02452_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[202] ));
 sky130_fd_sc_hd__dfrtp_2 _28655_ (.CLK(clk),
    .D(_02453_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[203] ));
 sky130_fd_sc_hd__dfrtp_2 _28656_ (.CLK(clk),
    .D(_02454_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[204] ));
 sky130_fd_sc_hd__dfrtp_2 _28657_ (.CLK(clk),
    .D(_02455_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[205] ));
 sky130_fd_sc_hd__dfrtp_2 _28658_ (.CLK(clk),
    .D(_02456_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[206] ));
 sky130_fd_sc_hd__dfrtp_2 _28659_ (.CLK(clk),
    .D(_02457_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[207] ));
 sky130_fd_sc_hd__dfrtp_2 _28660_ (.CLK(clk),
    .D(_02458_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[208] ));
 sky130_fd_sc_hd__dfrtp_2 _28661_ (.CLK(clk),
    .D(_02459_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[209] ));
 sky130_fd_sc_hd__dfrtp_2 _28662_ (.CLK(clk),
    .D(_02460_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[210] ));
 sky130_fd_sc_hd__dfrtp_2 _28663_ (.CLK(clk),
    .D(_02461_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[211] ));
 sky130_fd_sc_hd__dfrtp_2 _28664_ (.CLK(clk),
    .D(_02462_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[212] ));
 sky130_fd_sc_hd__dfrtp_2 _28665_ (.CLK(clk),
    .D(_02463_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[213] ));
 sky130_fd_sc_hd__dfrtp_2 _28666_ (.CLK(clk),
    .D(_02464_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[214] ));
 sky130_fd_sc_hd__dfrtp_2 _28667_ (.CLK(clk),
    .D(_02465_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[215] ));
 sky130_fd_sc_hd__dfrtp_2 _28668_ (.CLK(clk),
    .D(_02466_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[216] ));
 sky130_fd_sc_hd__dfrtp_2 _28669_ (.CLK(clk),
    .D(_02467_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[217] ));
 sky130_fd_sc_hd__dfrtp_2 _28670_ (.CLK(clk),
    .D(_02468_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[218] ));
 sky130_fd_sc_hd__dfrtp_2 _28671_ (.CLK(clk),
    .D(_02469_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[219] ));
 sky130_fd_sc_hd__dfrtp_2 _28672_ (.CLK(clk),
    .D(_02470_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[220] ));
 sky130_fd_sc_hd__dfrtp_2 _28673_ (.CLK(clk),
    .D(_02471_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[221] ));
 sky130_fd_sc_hd__dfrtp_2 _28674_ (.CLK(clk),
    .D(_02472_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[222] ));
 sky130_fd_sc_hd__dfrtp_2 _28675_ (.CLK(clk),
    .D(_02473_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[223] ));
 sky130_fd_sc_hd__dfrtp_2 _28676_ (.CLK(clk),
    .D(_02474_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[224] ));
 sky130_fd_sc_hd__dfrtp_2 _28677_ (.CLK(clk),
    .D(_02475_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[225] ));
 sky130_fd_sc_hd__dfrtp_2 _28678_ (.CLK(clk),
    .D(_02476_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[226] ));
 sky130_fd_sc_hd__dfrtp_2 _28679_ (.CLK(clk),
    .D(_02477_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[227] ));
 sky130_fd_sc_hd__dfrtp_2 _28680_ (.CLK(clk),
    .D(_02478_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[228] ));
 sky130_fd_sc_hd__dfrtp_2 _28681_ (.CLK(clk),
    .D(_02479_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[229] ));
 sky130_fd_sc_hd__dfrtp_2 _28682_ (.CLK(clk),
    .D(_02480_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[230] ));
 sky130_fd_sc_hd__dfrtp_2 _28683_ (.CLK(clk),
    .D(_02481_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[231] ));
 sky130_fd_sc_hd__dfrtp_2 _28684_ (.CLK(clk),
    .D(_02482_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[232] ));
 sky130_fd_sc_hd__dfrtp_2 _28685_ (.CLK(clk),
    .D(_02483_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[233] ));
 sky130_fd_sc_hd__dfrtp_2 _28686_ (.CLK(clk),
    .D(_02484_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[234] ));
 sky130_fd_sc_hd__dfrtp_2 _28687_ (.CLK(clk),
    .D(_02485_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[235] ));
 sky130_fd_sc_hd__dfrtp_2 _28688_ (.CLK(clk),
    .D(_02486_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[236] ));
 sky130_fd_sc_hd__dfrtp_2 _28689_ (.CLK(clk),
    .D(_02487_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[237] ));
 sky130_fd_sc_hd__dfrtp_2 _28690_ (.CLK(clk),
    .D(_02488_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[238] ));
 sky130_fd_sc_hd__dfrtp_2 _28691_ (.CLK(clk),
    .D(_02489_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[239] ));
 sky130_fd_sc_hd__dfrtp_2 _28692_ (.CLK(clk),
    .D(_02490_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[240] ));
 sky130_fd_sc_hd__dfrtp_2 _28693_ (.CLK(clk),
    .D(_02491_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[241] ));
 sky130_fd_sc_hd__dfrtp_2 _28694_ (.CLK(clk),
    .D(_02492_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[242] ));
 sky130_fd_sc_hd__dfrtp_2 _28695_ (.CLK(clk),
    .D(_02493_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[243] ));
 sky130_fd_sc_hd__dfrtp_2 _28696_ (.CLK(clk),
    .D(_02494_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[244] ));
 sky130_fd_sc_hd__dfrtp_2 _28697_ (.CLK(clk),
    .D(_02495_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[245] ));
 sky130_fd_sc_hd__dfrtp_2 _28698_ (.CLK(clk),
    .D(_02496_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[246] ));
 sky130_fd_sc_hd__dfrtp_2 _28699_ (.CLK(clk),
    .D(_02497_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[247] ));
 sky130_fd_sc_hd__dfrtp_2 _28700_ (.CLK(clk),
    .D(_02498_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[248] ));
 sky130_fd_sc_hd__dfrtp_2 _28701_ (.CLK(clk),
    .D(_02499_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[249] ));
 sky130_fd_sc_hd__dfrtp_2 _28702_ (.CLK(clk),
    .D(_02500_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[250] ));
 sky130_fd_sc_hd__dfrtp_2 _28703_ (.CLK(clk),
    .D(_02501_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[251] ));
 sky130_fd_sc_hd__dfrtp_2 _28704_ (.CLK(clk),
    .D(_02502_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[252] ));
 sky130_fd_sc_hd__dfrtp_2 _28705_ (.CLK(clk),
    .D(_02503_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[253] ));
 sky130_fd_sc_hd__dfrtp_2 _28706_ (.CLK(clk),
    .D(_02504_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[254] ));
 sky130_fd_sc_hd__dfrtp_2 _28707_ (.CLK(clk),
    .D(_02505_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[255] ));
 sky130_fd_sc_hd__dfrtp_2 _28708_ (.CLK(clk),
    .D(_02506_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[256] ));
 sky130_fd_sc_hd__dfrtp_2 _28709_ (.CLK(clk),
    .D(_02507_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[257] ));
 sky130_fd_sc_hd__dfrtp_2 _28710_ (.CLK(clk),
    .D(_02508_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[258] ));
 sky130_fd_sc_hd__dfrtp_2 _28711_ (.CLK(clk),
    .D(_02509_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[259] ));
 sky130_fd_sc_hd__dfrtp_2 _28712_ (.CLK(clk),
    .D(_02510_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[260] ));
 sky130_fd_sc_hd__dfrtp_2 _28713_ (.CLK(clk),
    .D(_02511_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[261] ));
 sky130_fd_sc_hd__dfrtp_2 _28714_ (.CLK(clk),
    .D(_02512_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[262] ));
 sky130_fd_sc_hd__dfrtp_2 _28715_ (.CLK(clk),
    .D(_02513_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[263] ));
 sky130_fd_sc_hd__dfrtp_2 _28716_ (.CLK(clk),
    .D(_02514_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[264] ));
 sky130_fd_sc_hd__dfrtp_2 _28717_ (.CLK(clk),
    .D(_02515_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[265] ));
 sky130_fd_sc_hd__dfrtp_2 _28718_ (.CLK(clk),
    .D(_02516_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[266] ));
 sky130_fd_sc_hd__dfrtp_2 _28719_ (.CLK(clk),
    .D(_02517_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[267] ));
 sky130_fd_sc_hd__dfrtp_2 _28720_ (.CLK(clk),
    .D(_02518_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[268] ));
 sky130_fd_sc_hd__dfrtp_2 _28721_ (.CLK(clk),
    .D(_02519_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[269] ));
 sky130_fd_sc_hd__dfrtp_2 _28722_ (.CLK(clk),
    .D(_02520_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[270] ));
 sky130_fd_sc_hd__dfrtp_2 _28723_ (.CLK(clk),
    .D(_02521_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[271] ));
 sky130_fd_sc_hd__dfrtp_2 _28724_ (.CLK(clk),
    .D(_02522_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[272] ));
 sky130_fd_sc_hd__dfrtp_2 _28725_ (.CLK(clk),
    .D(_02523_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[273] ));
 sky130_fd_sc_hd__dfrtp_2 _28726_ (.CLK(clk),
    .D(_02524_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[274] ));
 sky130_fd_sc_hd__dfrtp_2 _28727_ (.CLK(clk),
    .D(_02525_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[275] ));
 sky130_fd_sc_hd__dfrtp_2 _28728_ (.CLK(clk),
    .D(_02526_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[276] ));
 sky130_fd_sc_hd__dfrtp_2 _28729_ (.CLK(clk),
    .D(_02527_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[277] ));
 sky130_fd_sc_hd__dfrtp_2 _28730_ (.CLK(clk),
    .D(_02528_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[278] ));
 sky130_fd_sc_hd__dfrtp_2 _28731_ (.CLK(clk),
    .D(_02529_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[279] ));
 sky130_fd_sc_hd__dfrtp_2 _28732_ (.CLK(clk),
    .D(_02530_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[280] ));
 sky130_fd_sc_hd__dfrtp_2 _28733_ (.CLK(clk),
    .D(_02531_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[281] ));
 sky130_fd_sc_hd__dfrtp_2 _28734_ (.CLK(clk),
    .D(_02532_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[282] ));
 sky130_fd_sc_hd__dfrtp_2 _28735_ (.CLK(clk),
    .D(_02533_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[283] ));
 sky130_fd_sc_hd__dfrtp_2 _28736_ (.CLK(clk),
    .D(_02534_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[284] ));
 sky130_fd_sc_hd__dfrtp_2 _28737_ (.CLK(clk),
    .D(_02535_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[285] ));
 sky130_fd_sc_hd__dfrtp_2 _28738_ (.CLK(clk),
    .D(_02536_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[286] ));
 sky130_fd_sc_hd__dfrtp_2 _28739_ (.CLK(clk),
    .D(_02537_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[287] ));
 sky130_fd_sc_hd__dfrtp_2 _28740_ (.CLK(clk),
    .D(_02538_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[288] ));
 sky130_fd_sc_hd__dfrtp_2 _28741_ (.CLK(clk),
    .D(_02539_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[289] ));
 sky130_fd_sc_hd__dfrtp_2 _28742_ (.CLK(clk),
    .D(_02540_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[290] ));
 sky130_fd_sc_hd__dfrtp_2 _28743_ (.CLK(clk),
    .D(_02541_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[291] ));
 sky130_fd_sc_hd__dfrtp_2 _28744_ (.CLK(clk),
    .D(_02542_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[292] ));
 sky130_fd_sc_hd__dfrtp_2 _28745_ (.CLK(clk),
    .D(_02543_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[293] ));
 sky130_fd_sc_hd__dfrtp_2 _28746_ (.CLK(clk),
    .D(_02544_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[294] ));
 sky130_fd_sc_hd__dfrtp_2 _28747_ (.CLK(clk),
    .D(_02545_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[295] ));
 sky130_fd_sc_hd__dfrtp_2 _28748_ (.CLK(clk),
    .D(_02546_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[296] ));
 sky130_fd_sc_hd__dfrtp_2 _28749_ (.CLK(clk),
    .D(_02547_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[297] ));
 sky130_fd_sc_hd__dfrtp_2 _28750_ (.CLK(clk),
    .D(_02548_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[298] ));
 sky130_fd_sc_hd__dfrtp_2 _28751_ (.CLK(clk),
    .D(_02549_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[299] ));
 sky130_fd_sc_hd__dfrtp_2 _28752_ (.CLK(clk),
    .D(_02550_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[300] ));
 sky130_fd_sc_hd__dfrtp_2 _28753_ (.CLK(clk),
    .D(_02551_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[301] ));
 sky130_fd_sc_hd__dfrtp_2 _28754_ (.CLK(clk),
    .D(_02552_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[302] ));
 sky130_fd_sc_hd__dfrtp_2 _28755_ (.CLK(clk),
    .D(_02553_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[303] ));
 sky130_fd_sc_hd__dfrtp_2 _28756_ (.CLK(clk),
    .D(_02554_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[304] ));
 sky130_fd_sc_hd__dfrtp_2 _28757_ (.CLK(clk),
    .D(_02555_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[305] ));
 sky130_fd_sc_hd__dfrtp_2 _28758_ (.CLK(clk),
    .D(_02556_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[306] ));
 sky130_fd_sc_hd__dfrtp_2 _28759_ (.CLK(clk),
    .D(_02557_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[307] ));
 sky130_fd_sc_hd__dfrtp_2 _28760_ (.CLK(clk),
    .D(_02558_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[308] ));
 sky130_fd_sc_hd__dfrtp_2 _28761_ (.CLK(clk),
    .D(_02559_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[309] ));
 sky130_fd_sc_hd__dfrtp_2 _28762_ (.CLK(clk),
    .D(_02560_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[310] ));
 sky130_fd_sc_hd__dfrtp_2 _28763_ (.CLK(clk),
    .D(_02561_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[311] ));
 sky130_fd_sc_hd__dfrtp_2 _28764_ (.CLK(clk),
    .D(_02562_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[312] ));
 sky130_fd_sc_hd__dfrtp_2 _28765_ (.CLK(clk),
    .D(_02563_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[313] ));
 sky130_fd_sc_hd__dfrtp_2 _28766_ (.CLK(clk),
    .D(_02564_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[314] ));
 sky130_fd_sc_hd__dfrtp_2 _28767_ (.CLK(clk),
    .D(_02565_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[315] ));
 sky130_fd_sc_hd__dfrtp_2 _28768_ (.CLK(clk),
    .D(_02566_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[316] ));
 sky130_fd_sc_hd__dfrtp_2 _28769_ (.CLK(clk),
    .D(_02567_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[317] ));
 sky130_fd_sc_hd__dfrtp_2 _28770_ (.CLK(clk),
    .D(_02568_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[318] ));
 sky130_fd_sc_hd__dfrtp_2 _28771_ (.CLK(clk),
    .D(_02569_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[319] ));
 sky130_fd_sc_hd__dfrtp_2 _28772_ (.CLK(clk),
    .D(_02570_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[320] ));
 sky130_fd_sc_hd__dfrtp_2 _28773_ (.CLK(clk),
    .D(_02571_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[321] ));
 sky130_fd_sc_hd__dfrtp_2 _28774_ (.CLK(clk),
    .D(_02572_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[322] ));
 sky130_fd_sc_hd__dfrtp_2 _28775_ (.CLK(clk),
    .D(_02573_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[323] ));
 sky130_fd_sc_hd__dfrtp_2 _28776_ (.CLK(clk),
    .D(_02574_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[324] ));
 sky130_fd_sc_hd__dfrtp_2 _28777_ (.CLK(clk),
    .D(_02575_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[325] ));
 sky130_fd_sc_hd__dfrtp_2 _28778_ (.CLK(clk),
    .D(_02576_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[326] ));
 sky130_fd_sc_hd__dfrtp_2 _28779_ (.CLK(clk),
    .D(_02577_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[327] ));
 sky130_fd_sc_hd__dfrtp_2 _28780_ (.CLK(clk),
    .D(_02578_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[328] ));
 sky130_fd_sc_hd__dfrtp_2 _28781_ (.CLK(clk),
    .D(_02579_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[329] ));
 sky130_fd_sc_hd__dfrtp_2 _28782_ (.CLK(clk),
    .D(_02580_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[330] ));
 sky130_fd_sc_hd__dfrtp_2 _28783_ (.CLK(clk),
    .D(_02581_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[331] ));
 sky130_fd_sc_hd__dfrtp_2 _28784_ (.CLK(clk),
    .D(_02582_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[332] ));
 sky130_fd_sc_hd__dfrtp_2 _28785_ (.CLK(clk),
    .D(_02583_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[333] ));
 sky130_fd_sc_hd__dfrtp_2 _28786_ (.CLK(clk),
    .D(_02584_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[334] ));
 sky130_fd_sc_hd__dfrtp_2 _28787_ (.CLK(clk),
    .D(_02585_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[335] ));
 sky130_fd_sc_hd__dfrtp_2 _28788_ (.CLK(clk),
    .D(_02586_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[336] ));
 sky130_fd_sc_hd__dfrtp_2 _28789_ (.CLK(clk),
    .D(_02587_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[337] ));
 sky130_fd_sc_hd__dfrtp_2 _28790_ (.CLK(clk),
    .D(_02588_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[338] ));
 sky130_fd_sc_hd__dfrtp_2 _28791_ (.CLK(clk),
    .D(_02589_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[339] ));
 sky130_fd_sc_hd__dfrtp_2 _28792_ (.CLK(clk),
    .D(_02590_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[340] ));
 sky130_fd_sc_hd__dfrtp_2 _28793_ (.CLK(clk),
    .D(_02591_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[341] ));
 sky130_fd_sc_hd__dfrtp_2 _28794_ (.CLK(clk),
    .D(_02592_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[342] ));
 sky130_fd_sc_hd__dfrtp_2 _28795_ (.CLK(clk),
    .D(_02593_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[343] ));
 sky130_fd_sc_hd__dfrtp_2 _28796_ (.CLK(clk),
    .D(_02594_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[344] ));
 sky130_fd_sc_hd__dfrtp_2 _28797_ (.CLK(clk),
    .D(_02595_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[345] ));
 sky130_fd_sc_hd__dfrtp_2 _28798_ (.CLK(clk),
    .D(_02596_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[346] ));
 sky130_fd_sc_hd__dfrtp_2 _28799_ (.CLK(clk),
    .D(_02597_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[347] ));
 sky130_fd_sc_hd__dfrtp_2 _28800_ (.CLK(clk),
    .D(_02598_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[348] ));
 sky130_fd_sc_hd__dfrtp_2 _28801_ (.CLK(clk),
    .D(_02599_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[349] ));
 sky130_fd_sc_hd__dfrtp_2 _28802_ (.CLK(clk),
    .D(_02600_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[350] ));
 sky130_fd_sc_hd__dfrtp_2 _28803_ (.CLK(clk),
    .D(_02601_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[351] ));
 sky130_fd_sc_hd__dfrtp_2 _28804_ (.CLK(clk),
    .D(_02602_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[352] ));
 sky130_fd_sc_hd__dfrtp_2 _28805_ (.CLK(clk),
    .D(_02603_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[353] ));
 sky130_fd_sc_hd__dfrtp_2 _28806_ (.CLK(clk),
    .D(_02604_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[354] ));
 sky130_fd_sc_hd__dfrtp_2 _28807_ (.CLK(clk),
    .D(_02605_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[355] ));
 sky130_fd_sc_hd__dfrtp_2 _28808_ (.CLK(clk),
    .D(_02606_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[356] ));
 sky130_fd_sc_hd__dfrtp_2 _28809_ (.CLK(clk),
    .D(_02607_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[357] ));
 sky130_fd_sc_hd__dfrtp_2 _28810_ (.CLK(clk),
    .D(_02608_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[358] ));
 sky130_fd_sc_hd__dfrtp_2 _28811_ (.CLK(clk),
    .D(_02609_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[359] ));
 sky130_fd_sc_hd__dfrtp_2 _28812_ (.CLK(clk),
    .D(_02610_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[360] ));
 sky130_fd_sc_hd__dfrtp_2 _28813_ (.CLK(clk),
    .D(_02611_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[361] ));
 sky130_fd_sc_hd__dfrtp_2 _28814_ (.CLK(clk),
    .D(_02612_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[362] ));
 sky130_fd_sc_hd__dfrtp_2 _28815_ (.CLK(clk),
    .D(_02613_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[363] ));
 sky130_fd_sc_hd__dfrtp_2 _28816_ (.CLK(clk),
    .D(_02614_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[364] ));
 sky130_fd_sc_hd__dfrtp_2 _28817_ (.CLK(clk),
    .D(_02615_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[365] ));
 sky130_fd_sc_hd__dfrtp_2 _28818_ (.CLK(clk),
    .D(_02616_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[366] ));
 sky130_fd_sc_hd__dfrtp_2 _28819_ (.CLK(clk),
    .D(_02617_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[367] ));
 sky130_fd_sc_hd__dfrtp_2 _28820_ (.CLK(clk),
    .D(_02618_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[368] ));
 sky130_fd_sc_hd__dfrtp_2 _28821_ (.CLK(clk),
    .D(_02619_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[369] ));
 sky130_fd_sc_hd__dfrtp_2 _28822_ (.CLK(clk),
    .D(_02620_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[370] ));
 sky130_fd_sc_hd__dfrtp_2 _28823_ (.CLK(clk),
    .D(_02621_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[371] ));
 sky130_fd_sc_hd__dfrtp_2 _28824_ (.CLK(clk),
    .D(_02622_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[372] ));
 sky130_fd_sc_hd__dfrtp_2 _28825_ (.CLK(clk),
    .D(_02623_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[373] ));
 sky130_fd_sc_hd__dfrtp_2 _28826_ (.CLK(clk),
    .D(_02624_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[374] ));
 sky130_fd_sc_hd__dfrtp_2 _28827_ (.CLK(clk),
    .D(_02625_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[375] ));
 sky130_fd_sc_hd__dfrtp_2 _28828_ (.CLK(clk),
    .D(_02626_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[376] ));
 sky130_fd_sc_hd__dfrtp_2 _28829_ (.CLK(clk),
    .D(_02627_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[377] ));
 sky130_fd_sc_hd__dfrtp_2 _28830_ (.CLK(clk),
    .D(_02628_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[378] ));
 sky130_fd_sc_hd__dfrtp_2 _28831_ (.CLK(clk),
    .D(_02629_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[379] ));
 sky130_fd_sc_hd__dfrtp_2 _28832_ (.CLK(clk),
    .D(_02630_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[380] ));
 sky130_fd_sc_hd__dfrtp_2 _28833_ (.CLK(clk),
    .D(_02631_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[381] ));
 sky130_fd_sc_hd__dfrtp_2 _28834_ (.CLK(clk),
    .D(_02632_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[382] ));
 sky130_fd_sc_hd__dfrtp_2 _28835_ (.CLK(clk),
    .D(_02633_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[383] ));
 sky130_fd_sc_hd__dfrtp_2 _28836_ (.CLK(clk),
    .D(_02634_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[384] ));
 sky130_fd_sc_hd__dfrtp_2 _28837_ (.CLK(clk),
    .D(_02635_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[385] ));
 sky130_fd_sc_hd__dfrtp_2 _28838_ (.CLK(clk),
    .D(_02636_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[386] ));
 sky130_fd_sc_hd__dfrtp_2 _28839_ (.CLK(clk),
    .D(_02637_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[387] ));
 sky130_fd_sc_hd__dfrtp_2 _28840_ (.CLK(clk),
    .D(_02638_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[388] ));
 sky130_fd_sc_hd__dfrtp_2 _28841_ (.CLK(clk),
    .D(_02639_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[389] ));
 sky130_fd_sc_hd__dfrtp_2 _28842_ (.CLK(clk),
    .D(_02640_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[390] ));
 sky130_fd_sc_hd__dfrtp_2 _28843_ (.CLK(clk),
    .D(_02641_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[391] ));
 sky130_fd_sc_hd__dfrtp_2 _28844_ (.CLK(clk),
    .D(_02642_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[392] ));
 sky130_fd_sc_hd__dfrtp_2 _28845_ (.CLK(clk),
    .D(_02643_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[393] ));
 sky130_fd_sc_hd__dfrtp_2 _28846_ (.CLK(clk),
    .D(_02644_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[394] ));
 sky130_fd_sc_hd__dfrtp_2 _28847_ (.CLK(clk),
    .D(_02645_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[395] ));
 sky130_fd_sc_hd__dfrtp_2 _28848_ (.CLK(clk),
    .D(_02646_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[396] ));
 sky130_fd_sc_hd__dfrtp_2 _28849_ (.CLK(clk),
    .D(_02647_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[397] ));
 sky130_fd_sc_hd__dfrtp_2 _28850_ (.CLK(clk),
    .D(_02648_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[398] ));
 sky130_fd_sc_hd__dfrtp_2 _28851_ (.CLK(clk),
    .D(_02649_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[399] ));
 sky130_fd_sc_hd__dfrtp_2 _28852_ (.CLK(clk),
    .D(_02650_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[400] ));
 sky130_fd_sc_hd__dfrtp_2 _28853_ (.CLK(clk),
    .D(_02651_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[401] ));
 sky130_fd_sc_hd__dfrtp_2 _28854_ (.CLK(clk),
    .D(_02652_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[402] ));
 sky130_fd_sc_hd__dfrtp_2 _28855_ (.CLK(clk),
    .D(_02653_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[403] ));
 sky130_fd_sc_hd__dfrtp_2 _28856_ (.CLK(clk),
    .D(_02654_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[404] ));
 sky130_fd_sc_hd__dfrtp_2 _28857_ (.CLK(clk),
    .D(_02655_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[405] ));
 sky130_fd_sc_hd__dfrtp_2 _28858_ (.CLK(clk),
    .D(_02656_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[406] ));
 sky130_fd_sc_hd__dfrtp_2 _28859_ (.CLK(clk),
    .D(_02657_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[407] ));
 sky130_fd_sc_hd__dfrtp_2 _28860_ (.CLK(clk),
    .D(_02658_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[408] ));
 sky130_fd_sc_hd__dfrtp_2 _28861_ (.CLK(clk),
    .D(_02659_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[409] ));
 sky130_fd_sc_hd__dfrtp_2 _28862_ (.CLK(clk),
    .D(_02660_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[410] ));
 sky130_fd_sc_hd__dfrtp_2 _28863_ (.CLK(clk),
    .D(_02661_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[411] ));
 sky130_fd_sc_hd__dfrtp_2 _28864_ (.CLK(clk),
    .D(_02662_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[412] ));
 sky130_fd_sc_hd__dfrtp_2 _28865_ (.CLK(clk),
    .D(_02663_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[413] ));
 sky130_fd_sc_hd__dfrtp_2 _28866_ (.CLK(clk),
    .D(_02664_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[414] ));
 sky130_fd_sc_hd__dfrtp_2 _28867_ (.CLK(clk),
    .D(_02665_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[415] ));
 sky130_fd_sc_hd__dfrtp_2 _28868_ (.CLK(clk),
    .D(_02666_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[416] ));
 sky130_fd_sc_hd__dfrtp_2 _28869_ (.CLK(clk),
    .D(_02667_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[417] ));
 sky130_fd_sc_hd__dfrtp_2 _28870_ (.CLK(clk),
    .D(_02668_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[418] ));
 sky130_fd_sc_hd__dfrtp_2 _28871_ (.CLK(clk),
    .D(_02669_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[419] ));
 sky130_fd_sc_hd__dfrtp_2 _28872_ (.CLK(clk),
    .D(_02670_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[420] ));
 sky130_fd_sc_hd__dfrtp_2 _28873_ (.CLK(clk),
    .D(_02671_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[421] ));
 sky130_fd_sc_hd__dfrtp_2 _28874_ (.CLK(clk),
    .D(_02672_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[422] ));
 sky130_fd_sc_hd__dfrtp_2 _28875_ (.CLK(clk),
    .D(_02673_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[423] ));
 sky130_fd_sc_hd__dfrtp_2 _28876_ (.CLK(clk),
    .D(_02674_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[424] ));
 sky130_fd_sc_hd__dfrtp_2 _28877_ (.CLK(clk),
    .D(_02675_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[425] ));
 sky130_fd_sc_hd__dfrtp_2 _28878_ (.CLK(clk),
    .D(_02676_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[426] ));
 sky130_fd_sc_hd__dfrtp_2 _28879_ (.CLK(clk),
    .D(_02677_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[427] ));
 sky130_fd_sc_hd__dfrtp_2 _28880_ (.CLK(clk),
    .D(_02678_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[428] ));
 sky130_fd_sc_hd__dfrtp_2 _28881_ (.CLK(clk),
    .D(_02679_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[429] ));
 sky130_fd_sc_hd__dfrtp_2 _28882_ (.CLK(clk),
    .D(_02680_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[430] ));
 sky130_fd_sc_hd__dfrtp_2 _28883_ (.CLK(clk),
    .D(_02681_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[431] ));
 sky130_fd_sc_hd__dfrtp_2 _28884_ (.CLK(clk),
    .D(_02682_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[432] ));
 sky130_fd_sc_hd__dfrtp_2 _28885_ (.CLK(clk),
    .D(_02683_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[433] ));
 sky130_fd_sc_hd__dfrtp_2 _28886_ (.CLK(clk),
    .D(_02684_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[434] ));
 sky130_fd_sc_hd__dfrtp_2 _28887_ (.CLK(clk),
    .D(_02685_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[435] ));
 sky130_fd_sc_hd__dfrtp_2 _28888_ (.CLK(clk),
    .D(_02686_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[436] ));
 sky130_fd_sc_hd__dfrtp_2 _28889_ (.CLK(clk),
    .D(_02687_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[437] ));
 sky130_fd_sc_hd__dfrtp_2 _28890_ (.CLK(clk),
    .D(_02688_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[438] ));
 sky130_fd_sc_hd__dfrtp_2 _28891_ (.CLK(clk),
    .D(_02689_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[439] ));
 sky130_fd_sc_hd__dfrtp_2 _28892_ (.CLK(clk),
    .D(_02690_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[440] ));
 sky130_fd_sc_hd__dfrtp_2 _28893_ (.CLK(clk),
    .D(_02691_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[441] ));
 sky130_fd_sc_hd__dfrtp_2 _28894_ (.CLK(clk),
    .D(_02692_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[442] ));
 sky130_fd_sc_hd__dfrtp_2 _28895_ (.CLK(clk),
    .D(_02693_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[443] ));
 sky130_fd_sc_hd__dfrtp_2 _28896_ (.CLK(clk),
    .D(_02694_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[444] ));
 sky130_fd_sc_hd__dfrtp_2 _28897_ (.CLK(clk),
    .D(_02695_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[445] ));
 sky130_fd_sc_hd__dfrtp_2 _28898_ (.CLK(clk),
    .D(_02696_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[446] ));
 sky130_fd_sc_hd__dfrtp_2 _28899_ (.CLK(clk),
    .D(_02697_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[447] ));
 sky130_fd_sc_hd__dfrtp_2 _28900_ (.CLK(clk),
    .D(_02698_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[448] ));
 sky130_fd_sc_hd__dfrtp_2 _28901_ (.CLK(clk),
    .D(_02699_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[449] ));
 sky130_fd_sc_hd__dfrtp_2 _28902_ (.CLK(clk),
    .D(_02700_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[450] ));
 sky130_fd_sc_hd__dfrtp_2 _28903_ (.CLK(clk),
    .D(_02701_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[451] ));
 sky130_fd_sc_hd__dfrtp_2 _28904_ (.CLK(clk),
    .D(_02702_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[452] ));
 sky130_fd_sc_hd__dfrtp_2 _28905_ (.CLK(clk),
    .D(_02703_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[453] ));
 sky130_fd_sc_hd__dfrtp_2 _28906_ (.CLK(clk),
    .D(_02704_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[454] ));
 sky130_fd_sc_hd__dfrtp_2 _28907_ (.CLK(clk),
    .D(_02705_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[455] ));
 sky130_fd_sc_hd__dfrtp_2 _28908_ (.CLK(clk),
    .D(_02706_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[456] ));
 sky130_fd_sc_hd__dfrtp_2 _28909_ (.CLK(clk),
    .D(_02707_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[457] ));
 sky130_fd_sc_hd__dfrtp_2 _28910_ (.CLK(clk),
    .D(_02708_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[458] ));
 sky130_fd_sc_hd__dfrtp_2 _28911_ (.CLK(clk),
    .D(_02709_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[459] ));
 sky130_fd_sc_hd__dfrtp_2 _28912_ (.CLK(clk),
    .D(_02710_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[460] ));
 sky130_fd_sc_hd__dfrtp_2 _28913_ (.CLK(clk),
    .D(_02711_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[461] ));
 sky130_fd_sc_hd__dfrtp_2 _28914_ (.CLK(clk),
    .D(_02712_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[462] ));
 sky130_fd_sc_hd__dfrtp_2 _28915_ (.CLK(clk),
    .D(_02713_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[463] ));
 sky130_fd_sc_hd__dfrtp_2 _28916_ (.CLK(clk),
    .D(_02714_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[464] ));
 sky130_fd_sc_hd__dfrtp_2 _28917_ (.CLK(clk),
    .D(_02715_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[465] ));
 sky130_fd_sc_hd__dfrtp_2 _28918_ (.CLK(clk),
    .D(_02716_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[466] ));
 sky130_fd_sc_hd__dfrtp_2 _28919_ (.CLK(clk),
    .D(_02717_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[467] ));
 sky130_fd_sc_hd__dfrtp_2 _28920_ (.CLK(clk),
    .D(_02718_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[468] ));
 sky130_fd_sc_hd__dfrtp_2 _28921_ (.CLK(clk),
    .D(_02719_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[469] ));
 sky130_fd_sc_hd__dfrtp_2 _28922_ (.CLK(clk),
    .D(_02720_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[470] ));
 sky130_fd_sc_hd__dfrtp_2 _28923_ (.CLK(clk),
    .D(_02721_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[471] ));
 sky130_fd_sc_hd__dfrtp_2 _28924_ (.CLK(clk),
    .D(_02722_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[472] ));
 sky130_fd_sc_hd__dfrtp_2 _28925_ (.CLK(clk),
    .D(_02723_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[473] ));
 sky130_fd_sc_hd__dfrtp_2 _28926_ (.CLK(clk),
    .D(_02724_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[474] ));
 sky130_fd_sc_hd__dfrtp_2 _28927_ (.CLK(clk),
    .D(_02725_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[475] ));
 sky130_fd_sc_hd__dfrtp_2 _28928_ (.CLK(clk),
    .D(_02726_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[476] ));
 sky130_fd_sc_hd__dfrtp_2 _28929_ (.CLK(clk),
    .D(_02727_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[477] ));
 sky130_fd_sc_hd__dfrtp_2 _28930_ (.CLK(clk),
    .D(_02728_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[478] ));
 sky130_fd_sc_hd__dfrtp_2 _28931_ (.CLK(clk),
    .D(_02729_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[479] ));
 sky130_fd_sc_hd__dfrtp_2 _28932_ (.CLK(clk),
    .D(_02730_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[480] ));
 sky130_fd_sc_hd__dfrtp_2 _28933_ (.CLK(clk),
    .D(_02731_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[481] ));
 sky130_fd_sc_hd__dfrtp_2 _28934_ (.CLK(clk),
    .D(_02732_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[482] ));
 sky130_fd_sc_hd__dfrtp_2 _28935_ (.CLK(clk),
    .D(_02733_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[483] ));
 sky130_fd_sc_hd__dfrtp_2 _28936_ (.CLK(clk),
    .D(_02734_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[484] ));
 sky130_fd_sc_hd__dfrtp_2 _28937_ (.CLK(clk),
    .D(_02735_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[485] ));
 sky130_fd_sc_hd__dfrtp_2 _28938_ (.CLK(clk),
    .D(_02736_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[486] ));
 sky130_fd_sc_hd__dfrtp_2 _28939_ (.CLK(clk),
    .D(_02737_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[487] ));
 sky130_fd_sc_hd__dfrtp_2 _28940_ (.CLK(clk),
    .D(_02738_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[488] ));
 sky130_fd_sc_hd__dfrtp_2 _28941_ (.CLK(clk),
    .D(_02739_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[489] ));
 sky130_fd_sc_hd__dfrtp_2 _28942_ (.CLK(clk),
    .D(_02740_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[490] ));
 sky130_fd_sc_hd__dfrtp_2 _28943_ (.CLK(clk),
    .D(_02741_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[491] ));
 sky130_fd_sc_hd__dfrtp_2 _28944_ (.CLK(clk),
    .D(_02742_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[492] ));
 sky130_fd_sc_hd__dfrtp_2 _28945_ (.CLK(clk),
    .D(_02743_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[493] ));
 sky130_fd_sc_hd__dfrtp_2 _28946_ (.CLK(clk),
    .D(_02744_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[494] ));
 sky130_fd_sc_hd__dfrtp_2 _28947_ (.CLK(clk),
    .D(_02745_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[495] ));
 sky130_fd_sc_hd__dfrtp_2 _28948_ (.CLK(clk),
    .D(_02746_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[496] ));
 sky130_fd_sc_hd__dfrtp_2 _28949_ (.CLK(clk),
    .D(_02747_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[497] ));
 sky130_fd_sc_hd__dfrtp_2 _28950_ (.CLK(clk),
    .D(_02748_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[498] ));
 sky130_fd_sc_hd__dfrtp_2 _28951_ (.CLK(clk),
    .D(_02749_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[499] ));
 sky130_fd_sc_hd__dfrtp_2 _28952_ (.CLK(clk),
    .D(_02750_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[500] ));
 sky130_fd_sc_hd__dfrtp_2 _28953_ (.CLK(clk),
    .D(_02751_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[501] ));
 sky130_fd_sc_hd__dfrtp_2 _28954_ (.CLK(clk),
    .D(_02752_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[502] ));
 sky130_fd_sc_hd__dfrtp_2 _28955_ (.CLK(clk),
    .D(_02753_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[503] ));
 sky130_fd_sc_hd__dfrtp_2 _28956_ (.CLK(clk),
    .D(_02754_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[504] ));
 sky130_fd_sc_hd__dfrtp_2 _28957_ (.CLK(clk),
    .D(_02755_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[505] ));
 sky130_fd_sc_hd__dfrtp_2 _28958_ (.CLK(clk),
    .D(_02756_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[506] ));
 sky130_fd_sc_hd__dfrtp_2 _28959_ (.CLK(clk),
    .D(_02757_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[507] ));
 sky130_fd_sc_hd__dfrtp_2 _28960_ (.CLK(clk),
    .D(_02758_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[508] ));
 sky130_fd_sc_hd__dfrtp_2 _28961_ (.CLK(clk),
    .D(_02759_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[509] ));
 sky130_fd_sc_hd__dfrtp_2 _28962_ (.CLK(clk),
    .D(_02760_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[510] ));
 sky130_fd_sc_hd__dfrtp_2 _28963_ (.CLK(clk),
    .D(_02761_),
    .RESET_B(rst_n),
    .Q(\ser_C.shift_reg[511] ));
 sky130_fd_sc_hd__dfxtp_2 _28964_ (.CLK(clk),
    .D(_02762_),
    .Q(\systolic_inst.B_shift[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28965_ (.CLK(clk),
    .D(_02763_),
    .Q(\systolic_inst.B_shift[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28966_ (.CLK(clk),
    .D(_02764_),
    .Q(\systolic_inst.B_shift[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28967_ (.CLK(clk),
    .D(_02765_),
    .Q(\systolic_inst.B_shift[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28968_ (.CLK(clk),
    .D(_02766_),
    .Q(\systolic_inst.B_shift[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28969_ (.CLK(clk),
    .D(_02767_),
    .Q(\systolic_inst.B_shift[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28970_ (.CLK(clk),
    .D(_02768_),
    .Q(\systolic_inst.B_shift[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28971_ (.CLK(clk),
    .D(_02769_),
    .Q(\systolic_inst.B_shift[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28972_ (.CLK(clk),
    .D(_02770_),
    .Q(\systolic_inst.A_shift[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28973_ (.CLK(clk),
    .D(_02771_),
    .Q(\systolic_inst.A_shift[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28974_ (.CLK(clk),
    .D(_02772_),
    .Q(\systolic_inst.A_shift[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28975_ (.CLK(clk),
    .D(_02773_),
    .Q(\systolic_inst.A_shift[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28976_ (.CLK(clk),
    .D(_02774_),
    .Q(\systolic_inst.A_shift[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28977_ (.CLK(clk),
    .D(_02775_),
    .Q(\systolic_inst.A_shift[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28978_ (.CLK(clk),
    .D(_02776_),
    .Q(\systolic_inst.A_shift[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28979_ (.CLK(clk),
    .D(_02777_),
    .Q(\systolic_inst.A_shift[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28980_ (.CLK(clk),
    .D(_02778_),
    .Q(\systolic_inst.A_shift[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28981_ (.CLK(clk),
    .D(_02779_),
    .Q(\systolic_inst.A_shift[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28982_ (.CLK(clk),
    .D(_02780_),
    .Q(\systolic_inst.A_shift[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28983_ (.CLK(clk),
    .D(_02781_),
    .Q(\systolic_inst.A_shift[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28984_ (.CLK(clk),
    .D(_02782_),
    .Q(\systolic_inst.A_shift[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28985_ (.CLK(clk),
    .D(_02783_),
    .Q(\systolic_inst.A_shift[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28986_ (.CLK(clk),
    .D(_02784_),
    .Q(\systolic_inst.A_shift[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28987_ (.CLK(clk),
    .D(_02785_),
    .Q(\systolic_inst.A_shift[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28988_ (.CLK(clk),
    .D(_02786_),
    .Q(\systolic_inst.A_shift[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28989_ (.CLK(clk),
    .D(_02787_),
    .Q(\systolic_inst.A_shift[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28990_ (.CLK(clk),
    .D(_02788_),
    .Q(\systolic_inst.A_shift[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28991_ (.CLK(clk),
    .D(_02789_),
    .Q(\systolic_inst.A_shift[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28992_ (.CLK(clk),
    .D(_02790_),
    .Q(\systolic_inst.A_shift[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28993_ (.CLK(clk),
    .D(_02791_),
    .Q(\systolic_inst.A_shift[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28994_ (.CLK(clk),
    .D(_02792_),
    .Q(\systolic_inst.A_shift[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28995_ (.CLK(clk),
    .D(_02793_),
    .Q(\systolic_inst.A_shift[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28996_ (.CLK(clk),
    .D(_02794_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _28997_ (.CLK(clk),
    .D(_02795_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_2 _28998_ (.CLK(clk),
    .D(_02796_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _28999_ (.CLK(clk),
    .D(_02797_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_2 _29000_ (.CLK(clk),
    .D(_02798_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _29001_ (.CLK(clk),
    .D(_02799_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_2 _29002_ (.CLK(clk),
    .D(_02800_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_2 _29003_ (.CLK(clk),
    .D(_02801_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_2 _29004_ (.CLK(clk),
    .D(_02802_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _29005_ (.CLK(clk),
    .D(_02803_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_2 _29006_ (.CLK(clk),
    .D(_02804_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_2 _29007_ (.CLK(clk),
    .D(_02805_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_2 _29008_ (.CLK(clk),
    .D(_02806_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_2 _29009_ (.CLK(clk),
    .D(_02807_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_2 _29010_ (.CLK(clk),
    .D(_02808_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_2 _29011_ (.CLK(clk),
    .D(_02809_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_2 _29012_ (.CLK(clk),
    .D(_02810_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[16] ));
 sky130_fd_sc_hd__dfrtp_2 _29013_ (.CLK(clk),
    .D(_02811_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[17] ));
 sky130_fd_sc_hd__dfrtp_2 _29014_ (.CLK(clk),
    .D(_02812_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[18] ));
 sky130_fd_sc_hd__dfrtp_2 _29015_ (.CLK(clk),
    .D(_02813_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[19] ));
 sky130_fd_sc_hd__dfrtp_2 _29016_ (.CLK(clk),
    .D(_02814_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[20] ));
 sky130_fd_sc_hd__dfrtp_2 _29017_ (.CLK(clk),
    .D(_02815_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[21] ));
 sky130_fd_sc_hd__dfrtp_2 _29018_ (.CLK(clk),
    .D(_02816_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[22] ));
 sky130_fd_sc_hd__dfrtp_2 _29019_ (.CLK(clk),
    .D(_02817_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[23] ));
 sky130_fd_sc_hd__dfrtp_2 _29020_ (.CLK(clk),
    .D(_02818_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[24] ));
 sky130_fd_sc_hd__dfrtp_2 _29021_ (.CLK(clk),
    .D(_02819_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[25] ));
 sky130_fd_sc_hd__dfrtp_2 _29022_ (.CLK(clk),
    .D(_02820_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[26] ));
 sky130_fd_sc_hd__dfrtp_2 _29023_ (.CLK(clk),
    .D(_02821_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[27] ));
 sky130_fd_sc_hd__dfrtp_2 _29024_ (.CLK(clk),
    .D(_02822_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[28] ));
 sky130_fd_sc_hd__dfrtp_2 _29025_ (.CLK(clk),
    .D(_02823_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[29] ));
 sky130_fd_sc_hd__dfrtp_2 _29026_ (.CLK(clk),
    .D(_02824_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[30] ));
 sky130_fd_sc_hd__dfrtp_2 _29027_ (.CLK(clk),
    .D(_02825_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.cycle_cnt[31] ));
 sky130_fd_sc_hd__dfrtp_2 _29028_ (.CLK(clk),
    .D(_02826_),
    .RESET_B(rst_n),
    .Q(\C_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _29029_ (.CLK(clk),
    .D(_02827_),
    .RESET_B(rst_n),
    .Q(\C_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _29030_ (.CLK(clk),
    .D(_02828_),
    .RESET_B(rst_n),
    .Q(\C_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _29031_ (.CLK(clk),
    .D(_02829_),
    .RESET_B(rst_n),
    .Q(\C_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _29032_ (.CLK(clk),
    .D(_02830_),
    .RESET_B(rst_n),
    .Q(\C_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _29033_ (.CLK(clk),
    .D(_02831_),
    .RESET_B(rst_n),
    .Q(\C_out[5] ));
 sky130_fd_sc_hd__dfrtp_2 _29034_ (.CLK(clk),
    .D(_02832_),
    .RESET_B(rst_n),
    .Q(\C_out[6] ));
 sky130_fd_sc_hd__dfrtp_2 _29035_ (.CLK(clk),
    .D(_02833_),
    .RESET_B(rst_n),
    .Q(\C_out[7] ));
 sky130_fd_sc_hd__dfrtp_2 _29036_ (.CLK(clk),
    .D(_02834_),
    .RESET_B(rst_n),
    .Q(\C_out[8] ));
 sky130_fd_sc_hd__dfrtp_2 _29037_ (.CLK(clk),
    .D(_02835_),
    .RESET_B(rst_n),
    .Q(\C_out[9] ));
 sky130_fd_sc_hd__dfrtp_2 _29038_ (.CLK(clk),
    .D(_02836_),
    .RESET_B(rst_n),
    .Q(\C_out[10] ));
 sky130_fd_sc_hd__dfrtp_2 _29039_ (.CLK(clk),
    .D(_02837_),
    .RESET_B(rst_n),
    .Q(\C_out[11] ));
 sky130_fd_sc_hd__dfrtp_2 _29040_ (.CLK(clk),
    .D(_02838_),
    .RESET_B(rst_n),
    .Q(\C_out[12] ));
 sky130_fd_sc_hd__dfrtp_2 _29041_ (.CLK(clk),
    .D(_02839_),
    .RESET_B(rst_n),
    .Q(\C_out[13] ));
 sky130_fd_sc_hd__dfrtp_2 _29042_ (.CLK(clk),
    .D(_02840_),
    .RESET_B(rst_n),
    .Q(\C_out[14] ));
 sky130_fd_sc_hd__dfrtp_2 _29043_ (.CLK(clk),
    .D(_02841_),
    .RESET_B(rst_n),
    .Q(\C_out[15] ));
 sky130_fd_sc_hd__dfrtp_2 _29044_ (.CLK(clk),
    .D(_02842_),
    .RESET_B(rst_n),
    .Q(\C_out[16] ));
 sky130_fd_sc_hd__dfrtp_2 _29045_ (.CLK(clk),
    .D(_02843_),
    .RESET_B(rst_n),
    .Q(\C_out[17] ));
 sky130_fd_sc_hd__dfrtp_2 _29046_ (.CLK(clk),
    .D(_02844_),
    .RESET_B(rst_n),
    .Q(\C_out[18] ));
 sky130_fd_sc_hd__dfrtp_2 _29047_ (.CLK(clk),
    .D(_02845_),
    .RESET_B(rst_n),
    .Q(\C_out[19] ));
 sky130_fd_sc_hd__dfrtp_2 _29048_ (.CLK(clk),
    .D(_02846_),
    .RESET_B(rst_n),
    .Q(\C_out[20] ));
 sky130_fd_sc_hd__dfrtp_2 _29049_ (.CLK(clk),
    .D(_02847_),
    .RESET_B(rst_n),
    .Q(\C_out[21] ));
 sky130_fd_sc_hd__dfrtp_2 _29050_ (.CLK(clk),
    .D(_02848_),
    .RESET_B(rst_n),
    .Q(\C_out[22] ));
 sky130_fd_sc_hd__dfrtp_2 _29051_ (.CLK(clk),
    .D(_02849_),
    .RESET_B(rst_n),
    .Q(\C_out[23] ));
 sky130_fd_sc_hd__dfrtp_2 _29052_ (.CLK(clk),
    .D(_02850_),
    .RESET_B(rst_n),
    .Q(\C_out[24] ));
 sky130_fd_sc_hd__dfrtp_2 _29053_ (.CLK(clk),
    .D(_02851_),
    .RESET_B(rst_n),
    .Q(\C_out[25] ));
 sky130_fd_sc_hd__dfrtp_2 _29054_ (.CLK(clk),
    .D(_02852_),
    .RESET_B(rst_n),
    .Q(\C_out[26] ));
 sky130_fd_sc_hd__dfrtp_2 _29055_ (.CLK(clk),
    .D(_02853_),
    .RESET_B(rst_n),
    .Q(\C_out[27] ));
 sky130_fd_sc_hd__dfrtp_2 _29056_ (.CLK(clk),
    .D(_02854_),
    .RESET_B(rst_n),
    .Q(\C_out[28] ));
 sky130_fd_sc_hd__dfrtp_2 _29057_ (.CLK(clk),
    .D(_02855_),
    .RESET_B(rst_n),
    .Q(\C_out[29] ));
 sky130_fd_sc_hd__dfrtp_2 _29058_ (.CLK(clk),
    .D(_02856_),
    .RESET_B(rst_n),
    .Q(\C_out[30] ));
 sky130_fd_sc_hd__dfrtp_2 _29059_ (.CLK(clk),
    .D(_02857_),
    .RESET_B(rst_n),
    .Q(\C_out[31] ));
 sky130_fd_sc_hd__dfrtp_2 _29060_ (.CLK(clk),
    .D(_02858_),
    .RESET_B(rst_n),
    .Q(\C_out[32] ));
 sky130_fd_sc_hd__dfrtp_2 _29061_ (.CLK(clk),
    .D(_02859_),
    .RESET_B(rst_n),
    .Q(\C_out[33] ));
 sky130_fd_sc_hd__dfrtp_2 _29062_ (.CLK(clk),
    .D(_02860_),
    .RESET_B(rst_n),
    .Q(\C_out[34] ));
 sky130_fd_sc_hd__dfrtp_2 _29063_ (.CLK(clk),
    .D(_02861_),
    .RESET_B(rst_n),
    .Q(\C_out[35] ));
 sky130_fd_sc_hd__dfrtp_2 _29064_ (.CLK(clk),
    .D(_02862_),
    .RESET_B(rst_n),
    .Q(\C_out[36] ));
 sky130_fd_sc_hd__dfrtp_2 _29065_ (.CLK(clk),
    .D(_02863_),
    .RESET_B(rst_n),
    .Q(\C_out[37] ));
 sky130_fd_sc_hd__dfrtp_2 _29066_ (.CLK(clk),
    .D(_02864_),
    .RESET_B(rst_n),
    .Q(\C_out[38] ));
 sky130_fd_sc_hd__dfrtp_2 _29067_ (.CLK(clk),
    .D(_02865_),
    .RESET_B(rst_n),
    .Q(\C_out[39] ));
 sky130_fd_sc_hd__dfrtp_2 _29068_ (.CLK(clk),
    .D(_02866_),
    .RESET_B(rst_n),
    .Q(\C_out[40] ));
 sky130_fd_sc_hd__dfrtp_2 _29069_ (.CLK(clk),
    .D(_02867_),
    .RESET_B(rst_n),
    .Q(\C_out[41] ));
 sky130_fd_sc_hd__dfrtp_2 _29070_ (.CLK(clk),
    .D(_02868_),
    .RESET_B(rst_n),
    .Q(\C_out[42] ));
 sky130_fd_sc_hd__dfrtp_2 _29071_ (.CLK(clk),
    .D(_02869_),
    .RESET_B(rst_n),
    .Q(\C_out[43] ));
 sky130_fd_sc_hd__dfrtp_2 _29072_ (.CLK(clk),
    .D(_02870_),
    .RESET_B(rst_n),
    .Q(\C_out[44] ));
 sky130_fd_sc_hd__dfrtp_2 _29073_ (.CLK(clk),
    .D(_02871_),
    .RESET_B(rst_n),
    .Q(\C_out[45] ));
 sky130_fd_sc_hd__dfrtp_2 _29074_ (.CLK(clk),
    .D(_02872_),
    .RESET_B(rst_n),
    .Q(\C_out[46] ));
 sky130_fd_sc_hd__dfrtp_2 _29075_ (.CLK(clk),
    .D(_02873_),
    .RESET_B(rst_n),
    .Q(\C_out[47] ));
 sky130_fd_sc_hd__dfrtp_2 _29076_ (.CLK(clk),
    .D(_02874_),
    .RESET_B(rst_n),
    .Q(\C_out[48] ));
 sky130_fd_sc_hd__dfrtp_2 _29077_ (.CLK(clk),
    .D(_02875_),
    .RESET_B(rst_n),
    .Q(\C_out[49] ));
 sky130_fd_sc_hd__dfrtp_2 _29078_ (.CLK(clk),
    .D(_02876_),
    .RESET_B(rst_n),
    .Q(\C_out[50] ));
 sky130_fd_sc_hd__dfrtp_2 _29079_ (.CLK(clk),
    .D(_02877_),
    .RESET_B(rst_n),
    .Q(\C_out[51] ));
 sky130_fd_sc_hd__dfrtp_2 _29080_ (.CLK(clk),
    .D(_02878_),
    .RESET_B(rst_n),
    .Q(\C_out[52] ));
 sky130_fd_sc_hd__dfrtp_2 _29081_ (.CLK(clk),
    .D(_02879_),
    .RESET_B(rst_n),
    .Q(\C_out[53] ));
 sky130_fd_sc_hd__dfrtp_2 _29082_ (.CLK(clk),
    .D(_02880_),
    .RESET_B(rst_n),
    .Q(\C_out[54] ));
 sky130_fd_sc_hd__dfrtp_2 _29083_ (.CLK(clk),
    .D(_02881_),
    .RESET_B(rst_n),
    .Q(\C_out[55] ));
 sky130_fd_sc_hd__dfrtp_2 _29084_ (.CLK(clk),
    .D(_02882_),
    .RESET_B(rst_n),
    .Q(\C_out[56] ));
 sky130_fd_sc_hd__dfrtp_2 _29085_ (.CLK(clk),
    .D(_02883_),
    .RESET_B(rst_n),
    .Q(\C_out[57] ));
 sky130_fd_sc_hd__dfrtp_2 _29086_ (.CLK(clk),
    .D(_02884_),
    .RESET_B(rst_n),
    .Q(\C_out[58] ));
 sky130_fd_sc_hd__dfrtp_2 _29087_ (.CLK(clk),
    .D(_02885_),
    .RESET_B(rst_n),
    .Q(\C_out[59] ));
 sky130_fd_sc_hd__dfrtp_2 _29088_ (.CLK(clk),
    .D(_02886_),
    .RESET_B(rst_n),
    .Q(\C_out[60] ));
 sky130_fd_sc_hd__dfrtp_2 _29089_ (.CLK(clk),
    .D(_02887_),
    .RESET_B(rst_n),
    .Q(\C_out[61] ));
 sky130_fd_sc_hd__dfrtp_2 _29090_ (.CLK(clk),
    .D(_02888_),
    .RESET_B(rst_n),
    .Q(\C_out[62] ));
 sky130_fd_sc_hd__dfrtp_2 _29091_ (.CLK(clk),
    .D(_02889_),
    .RESET_B(rst_n),
    .Q(\C_out[63] ));
 sky130_fd_sc_hd__dfrtp_2 _29092_ (.CLK(clk),
    .D(_02890_),
    .RESET_B(rst_n),
    .Q(\C_out[64] ));
 sky130_fd_sc_hd__dfrtp_2 _29093_ (.CLK(clk),
    .D(_02891_),
    .RESET_B(rst_n),
    .Q(\C_out[65] ));
 sky130_fd_sc_hd__dfrtp_2 _29094_ (.CLK(clk),
    .D(_02892_),
    .RESET_B(rst_n),
    .Q(\C_out[66] ));
 sky130_fd_sc_hd__dfrtp_2 _29095_ (.CLK(clk),
    .D(_02893_),
    .RESET_B(rst_n),
    .Q(\C_out[67] ));
 sky130_fd_sc_hd__dfrtp_2 _29096_ (.CLK(clk),
    .D(_02894_),
    .RESET_B(rst_n),
    .Q(\C_out[68] ));
 sky130_fd_sc_hd__dfrtp_2 _29097_ (.CLK(clk),
    .D(_02895_),
    .RESET_B(rst_n),
    .Q(\C_out[69] ));
 sky130_fd_sc_hd__dfrtp_2 _29098_ (.CLK(clk),
    .D(_02896_),
    .RESET_B(rst_n),
    .Q(\C_out[70] ));
 sky130_fd_sc_hd__dfrtp_2 _29099_ (.CLK(clk),
    .D(_02897_),
    .RESET_B(rst_n),
    .Q(\C_out[71] ));
 sky130_fd_sc_hd__dfrtp_2 _29100_ (.CLK(clk),
    .D(_02898_),
    .RESET_B(rst_n),
    .Q(\C_out[72] ));
 sky130_fd_sc_hd__dfrtp_2 _29101_ (.CLK(clk),
    .D(_02899_),
    .RESET_B(rst_n),
    .Q(\C_out[73] ));
 sky130_fd_sc_hd__dfrtp_2 _29102_ (.CLK(clk),
    .D(_02900_),
    .RESET_B(rst_n),
    .Q(\C_out[74] ));
 sky130_fd_sc_hd__dfrtp_2 _29103_ (.CLK(clk),
    .D(_02901_),
    .RESET_B(rst_n),
    .Q(\C_out[75] ));
 sky130_fd_sc_hd__dfrtp_2 _29104_ (.CLK(clk),
    .D(_02902_),
    .RESET_B(rst_n),
    .Q(\C_out[76] ));
 sky130_fd_sc_hd__dfrtp_2 _29105_ (.CLK(clk),
    .D(_02903_),
    .RESET_B(rst_n),
    .Q(\C_out[77] ));
 sky130_fd_sc_hd__dfrtp_2 _29106_ (.CLK(clk),
    .D(_02904_),
    .RESET_B(rst_n),
    .Q(\C_out[78] ));
 sky130_fd_sc_hd__dfrtp_2 _29107_ (.CLK(clk),
    .D(_02905_),
    .RESET_B(rst_n),
    .Q(\C_out[79] ));
 sky130_fd_sc_hd__dfrtp_2 _29108_ (.CLK(clk),
    .D(_02906_),
    .RESET_B(rst_n),
    .Q(\C_out[80] ));
 sky130_fd_sc_hd__dfrtp_2 _29109_ (.CLK(clk),
    .D(_02907_),
    .RESET_B(rst_n),
    .Q(\C_out[81] ));
 sky130_fd_sc_hd__dfrtp_2 _29110_ (.CLK(clk),
    .D(_02908_),
    .RESET_B(rst_n),
    .Q(\C_out[82] ));
 sky130_fd_sc_hd__dfrtp_2 _29111_ (.CLK(clk),
    .D(_02909_),
    .RESET_B(rst_n),
    .Q(\C_out[83] ));
 sky130_fd_sc_hd__dfrtp_2 _29112_ (.CLK(clk),
    .D(_02910_),
    .RESET_B(rst_n),
    .Q(\C_out[84] ));
 sky130_fd_sc_hd__dfrtp_2 _29113_ (.CLK(clk),
    .D(_02911_),
    .RESET_B(rst_n),
    .Q(\C_out[85] ));
 sky130_fd_sc_hd__dfrtp_2 _29114_ (.CLK(clk),
    .D(_02912_),
    .RESET_B(rst_n),
    .Q(\C_out[86] ));
 sky130_fd_sc_hd__dfrtp_2 _29115_ (.CLK(clk),
    .D(_02913_),
    .RESET_B(rst_n),
    .Q(\C_out[87] ));
 sky130_fd_sc_hd__dfrtp_2 _29116_ (.CLK(clk),
    .D(_02914_),
    .RESET_B(rst_n),
    .Q(\C_out[88] ));
 sky130_fd_sc_hd__dfrtp_2 _29117_ (.CLK(clk),
    .D(_02915_),
    .RESET_B(rst_n),
    .Q(\C_out[89] ));
 sky130_fd_sc_hd__dfrtp_2 _29118_ (.CLK(clk),
    .D(_02916_),
    .RESET_B(rst_n),
    .Q(\C_out[90] ));
 sky130_fd_sc_hd__dfrtp_2 _29119_ (.CLK(clk),
    .D(_02917_),
    .RESET_B(rst_n),
    .Q(\C_out[91] ));
 sky130_fd_sc_hd__dfrtp_2 _29120_ (.CLK(clk),
    .D(_02918_),
    .RESET_B(rst_n),
    .Q(\C_out[92] ));
 sky130_fd_sc_hd__dfrtp_2 _29121_ (.CLK(clk),
    .D(_02919_),
    .RESET_B(rst_n),
    .Q(\C_out[93] ));
 sky130_fd_sc_hd__dfrtp_2 _29122_ (.CLK(clk),
    .D(_02920_),
    .RESET_B(rst_n),
    .Q(\C_out[94] ));
 sky130_fd_sc_hd__dfrtp_2 _29123_ (.CLK(clk),
    .D(_02921_),
    .RESET_B(rst_n),
    .Q(\C_out[95] ));
 sky130_fd_sc_hd__dfrtp_2 _29124_ (.CLK(clk),
    .D(_02922_),
    .RESET_B(rst_n),
    .Q(\C_out[96] ));
 sky130_fd_sc_hd__dfrtp_2 _29125_ (.CLK(clk),
    .D(_02923_),
    .RESET_B(rst_n),
    .Q(\C_out[97] ));
 sky130_fd_sc_hd__dfrtp_2 _29126_ (.CLK(clk),
    .D(_02924_),
    .RESET_B(rst_n),
    .Q(\C_out[98] ));
 sky130_fd_sc_hd__dfrtp_2 _29127_ (.CLK(clk),
    .D(_02925_),
    .RESET_B(rst_n),
    .Q(\C_out[99] ));
 sky130_fd_sc_hd__dfrtp_2 _29128_ (.CLK(clk),
    .D(_02926_),
    .RESET_B(rst_n),
    .Q(\C_out[100] ));
 sky130_fd_sc_hd__dfrtp_2 _29129_ (.CLK(clk),
    .D(_02927_),
    .RESET_B(rst_n),
    .Q(\C_out[101] ));
 sky130_fd_sc_hd__dfrtp_2 _29130_ (.CLK(clk),
    .D(_02928_),
    .RESET_B(rst_n),
    .Q(\C_out[102] ));
 sky130_fd_sc_hd__dfrtp_2 _29131_ (.CLK(clk),
    .D(_02929_),
    .RESET_B(rst_n),
    .Q(\C_out[103] ));
 sky130_fd_sc_hd__dfrtp_2 _29132_ (.CLK(clk),
    .D(_02930_),
    .RESET_B(rst_n),
    .Q(\C_out[104] ));
 sky130_fd_sc_hd__dfrtp_2 _29133_ (.CLK(clk),
    .D(_02931_),
    .RESET_B(rst_n),
    .Q(\C_out[105] ));
 sky130_fd_sc_hd__dfrtp_2 _29134_ (.CLK(clk),
    .D(_02932_),
    .RESET_B(rst_n),
    .Q(\C_out[106] ));
 sky130_fd_sc_hd__dfrtp_2 _29135_ (.CLK(clk),
    .D(_02933_),
    .RESET_B(rst_n),
    .Q(\C_out[107] ));
 sky130_fd_sc_hd__dfrtp_2 _29136_ (.CLK(clk),
    .D(_02934_),
    .RESET_B(rst_n),
    .Q(\C_out[108] ));
 sky130_fd_sc_hd__dfrtp_2 _29137_ (.CLK(clk),
    .D(_02935_),
    .RESET_B(rst_n),
    .Q(\C_out[109] ));
 sky130_fd_sc_hd__dfrtp_2 _29138_ (.CLK(clk),
    .D(_02936_),
    .RESET_B(rst_n),
    .Q(\C_out[110] ));
 sky130_fd_sc_hd__dfrtp_2 _29139_ (.CLK(clk),
    .D(_02937_),
    .RESET_B(rst_n),
    .Q(\C_out[111] ));
 sky130_fd_sc_hd__dfrtp_2 _29140_ (.CLK(clk),
    .D(_02938_),
    .RESET_B(rst_n),
    .Q(\C_out[112] ));
 sky130_fd_sc_hd__dfrtp_2 _29141_ (.CLK(clk),
    .D(_02939_),
    .RESET_B(rst_n),
    .Q(\C_out[113] ));
 sky130_fd_sc_hd__dfrtp_2 _29142_ (.CLK(clk),
    .D(_02940_),
    .RESET_B(rst_n),
    .Q(\C_out[114] ));
 sky130_fd_sc_hd__dfrtp_2 _29143_ (.CLK(clk),
    .D(_02941_),
    .RESET_B(rst_n),
    .Q(\C_out[115] ));
 sky130_fd_sc_hd__dfrtp_2 _29144_ (.CLK(clk),
    .D(_02942_),
    .RESET_B(rst_n),
    .Q(\C_out[116] ));
 sky130_fd_sc_hd__dfrtp_2 _29145_ (.CLK(clk),
    .D(_02943_),
    .RESET_B(rst_n),
    .Q(\C_out[117] ));
 sky130_fd_sc_hd__dfrtp_2 _29146_ (.CLK(clk),
    .D(_02944_),
    .RESET_B(rst_n),
    .Q(\C_out[118] ));
 sky130_fd_sc_hd__dfrtp_2 _29147_ (.CLK(clk),
    .D(_02945_),
    .RESET_B(rst_n),
    .Q(\C_out[119] ));
 sky130_fd_sc_hd__dfrtp_2 _29148_ (.CLK(clk),
    .D(_02946_),
    .RESET_B(rst_n),
    .Q(\C_out[120] ));
 sky130_fd_sc_hd__dfrtp_2 _29149_ (.CLK(clk),
    .D(_02947_),
    .RESET_B(rst_n),
    .Q(\C_out[121] ));
 sky130_fd_sc_hd__dfrtp_2 _29150_ (.CLK(clk),
    .D(_02948_),
    .RESET_B(rst_n),
    .Q(\C_out[122] ));
 sky130_fd_sc_hd__dfrtp_2 _29151_ (.CLK(clk),
    .D(_02949_),
    .RESET_B(rst_n),
    .Q(\C_out[123] ));
 sky130_fd_sc_hd__dfrtp_2 _29152_ (.CLK(clk),
    .D(_02950_),
    .RESET_B(rst_n),
    .Q(\C_out[124] ));
 sky130_fd_sc_hd__dfrtp_2 _29153_ (.CLK(clk),
    .D(_02951_),
    .RESET_B(rst_n),
    .Q(\C_out[125] ));
 sky130_fd_sc_hd__dfrtp_2 _29154_ (.CLK(clk),
    .D(_02952_),
    .RESET_B(rst_n),
    .Q(\C_out[126] ));
 sky130_fd_sc_hd__dfrtp_2 _29155_ (.CLK(clk),
    .D(_02953_),
    .RESET_B(rst_n),
    .Q(\C_out[127] ));
 sky130_fd_sc_hd__dfrtp_2 _29156_ (.CLK(clk),
    .D(_02954_),
    .RESET_B(rst_n),
    .Q(\C_out[128] ));
 sky130_fd_sc_hd__dfrtp_2 _29157_ (.CLK(clk),
    .D(_02955_),
    .RESET_B(rst_n),
    .Q(\C_out[129] ));
 sky130_fd_sc_hd__dfrtp_2 _29158_ (.CLK(clk),
    .D(_02956_),
    .RESET_B(rst_n),
    .Q(\C_out[130] ));
 sky130_fd_sc_hd__dfrtp_2 _29159_ (.CLK(clk),
    .D(_02957_),
    .RESET_B(rst_n),
    .Q(\C_out[131] ));
 sky130_fd_sc_hd__dfrtp_2 _29160_ (.CLK(clk),
    .D(_02958_),
    .RESET_B(rst_n),
    .Q(\C_out[132] ));
 sky130_fd_sc_hd__dfrtp_2 _29161_ (.CLK(clk),
    .D(_02959_),
    .RESET_B(rst_n),
    .Q(\C_out[133] ));
 sky130_fd_sc_hd__dfrtp_2 _29162_ (.CLK(clk),
    .D(_02960_),
    .RESET_B(rst_n),
    .Q(\C_out[134] ));
 sky130_fd_sc_hd__dfrtp_2 _29163_ (.CLK(clk),
    .D(_02961_),
    .RESET_B(rst_n),
    .Q(\C_out[135] ));
 sky130_fd_sc_hd__dfrtp_2 _29164_ (.CLK(clk),
    .D(_02962_),
    .RESET_B(rst_n),
    .Q(\C_out[136] ));
 sky130_fd_sc_hd__dfrtp_2 _29165_ (.CLK(clk),
    .D(_02963_),
    .RESET_B(rst_n),
    .Q(\C_out[137] ));
 sky130_fd_sc_hd__dfrtp_2 _29166_ (.CLK(clk),
    .D(_02964_),
    .RESET_B(rst_n),
    .Q(\C_out[138] ));
 sky130_fd_sc_hd__dfrtp_2 _29167_ (.CLK(clk),
    .D(_02965_),
    .RESET_B(rst_n),
    .Q(\C_out[139] ));
 sky130_fd_sc_hd__dfrtp_2 _29168_ (.CLK(clk),
    .D(_02966_),
    .RESET_B(rst_n),
    .Q(\C_out[140] ));
 sky130_fd_sc_hd__dfrtp_2 _29169_ (.CLK(clk),
    .D(_02967_),
    .RESET_B(rst_n),
    .Q(\C_out[141] ));
 sky130_fd_sc_hd__dfrtp_2 _29170_ (.CLK(clk),
    .D(_02968_),
    .RESET_B(rst_n),
    .Q(\C_out[142] ));
 sky130_fd_sc_hd__dfrtp_2 _29171_ (.CLK(clk),
    .D(_02969_),
    .RESET_B(rst_n),
    .Q(\C_out[143] ));
 sky130_fd_sc_hd__dfrtp_2 _29172_ (.CLK(clk),
    .D(_02970_),
    .RESET_B(rst_n),
    .Q(\C_out[144] ));
 sky130_fd_sc_hd__dfrtp_2 _29173_ (.CLK(clk),
    .D(_02971_),
    .RESET_B(rst_n),
    .Q(\C_out[145] ));
 sky130_fd_sc_hd__dfrtp_2 _29174_ (.CLK(clk),
    .D(_02972_),
    .RESET_B(rst_n),
    .Q(\C_out[146] ));
 sky130_fd_sc_hd__dfrtp_2 _29175_ (.CLK(clk),
    .D(_02973_),
    .RESET_B(rst_n),
    .Q(\C_out[147] ));
 sky130_fd_sc_hd__dfrtp_2 _29176_ (.CLK(clk),
    .D(_02974_),
    .RESET_B(rst_n),
    .Q(\C_out[148] ));
 sky130_fd_sc_hd__dfrtp_2 _29177_ (.CLK(clk),
    .D(_02975_),
    .RESET_B(rst_n),
    .Q(\C_out[149] ));
 sky130_fd_sc_hd__dfrtp_2 _29178_ (.CLK(clk),
    .D(_02976_),
    .RESET_B(rst_n),
    .Q(\C_out[150] ));
 sky130_fd_sc_hd__dfrtp_2 _29179_ (.CLK(clk),
    .D(_02977_),
    .RESET_B(rst_n),
    .Q(\C_out[151] ));
 sky130_fd_sc_hd__dfrtp_2 _29180_ (.CLK(clk),
    .D(_02978_),
    .RESET_B(rst_n),
    .Q(\C_out[152] ));
 sky130_fd_sc_hd__dfrtp_2 _29181_ (.CLK(clk),
    .D(_02979_),
    .RESET_B(rst_n),
    .Q(\C_out[153] ));
 sky130_fd_sc_hd__dfrtp_2 _29182_ (.CLK(clk),
    .D(_02980_),
    .RESET_B(rst_n),
    .Q(\C_out[154] ));
 sky130_fd_sc_hd__dfrtp_2 _29183_ (.CLK(clk),
    .D(_02981_),
    .RESET_B(rst_n),
    .Q(\C_out[155] ));
 sky130_fd_sc_hd__dfrtp_2 _29184_ (.CLK(clk),
    .D(_02982_),
    .RESET_B(rst_n),
    .Q(\C_out[156] ));
 sky130_fd_sc_hd__dfrtp_2 _29185_ (.CLK(clk),
    .D(_02983_),
    .RESET_B(rst_n),
    .Q(\C_out[157] ));
 sky130_fd_sc_hd__dfrtp_2 _29186_ (.CLK(clk),
    .D(_02984_),
    .RESET_B(rst_n),
    .Q(\C_out[158] ));
 sky130_fd_sc_hd__dfrtp_2 _29187_ (.CLK(clk),
    .D(_02985_),
    .RESET_B(rst_n),
    .Q(\C_out[159] ));
 sky130_fd_sc_hd__dfrtp_2 _29188_ (.CLK(clk),
    .D(_02986_),
    .RESET_B(rst_n),
    .Q(\C_out[160] ));
 sky130_fd_sc_hd__dfrtp_2 _29189_ (.CLK(clk),
    .D(_02987_),
    .RESET_B(rst_n),
    .Q(\C_out[161] ));
 sky130_fd_sc_hd__dfrtp_2 _29190_ (.CLK(clk),
    .D(_02988_),
    .RESET_B(rst_n),
    .Q(\C_out[162] ));
 sky130_fd_sc_hd__dfrtp_2 _29191_ (.CLK(clk),
    .D(_02989_),
    .RESET_B(rst_n),
    .Q(\C_out[163] ));
 sky130_fd_sc_hd__dfrtp_2 _29192_ (.CLK(clk),
    .D(_02990_),
    .RESET_B(rst_n),
    .Q(\C_out[164] ));
 sky130_fd_sc_hd__dfrtp_2 _29193_ (.CLK(clk),
    .D(_02991_),
    .RESET_B(rst_n),
    .Q(\C_out[165] ));
 sky130_fd_sc_hd__dfrtp_2 _29194_ (.CLK(clk),
    .D(_02992_),
    .RESET_B(rst_n),
    .Q(\C_out[166] ));
 sky130_fd_sc_hd__dfrtp_2 _29195_ (.CLK(clk),
    .D(_02993_),
    .RESET_B(rst_n),
    .Q(\C_out[167] ));
 sky130_fd_sc_hd__dfrtp_2 _29196_ (.CLK(clk),
    .D(_02994_),
    .RESET_B(rst_n),
    .Q(\C_out[168] ));
 sky130_fd_sc_hd__dfrtp_2 _29197_ (.CLK(clk),
    .D(_02995_),
    .RESET_B(rst_n),
    .Q(\C_out[169] ));
 sky130_fd_sc_hd__dfrtp_2 _29198_ (.CLK(clk),
    .D(_02996_),
    .RESET_B(rst_n),
    .Q(\C_out[170] ));
 sky130_fd_sc_hd__dfrtp_2 _29199_ (.CLK(clk),
    .D(_02997_),
    .RESET_B(rst_n),
    .Q(\C_out[171] ));
 sky130_fd_sc_hd__dfrtp_2 _29200_ (.CLK(clk),
    .D(_02998_),
    .RESET_B(rst_n),
    .Q(\C_out[172] ));
 sky130_fd_sc_hd__dfrtp_2 _29201_ (.CLK(clk),
    .D(_02999_),
    .RESET_B(rst_n),
    .Q(\C_out[173] ));
 sky130_fd_sc_hd__dfrtp_2 _29202_ (.CLK(clk),
    .D(_03000_),
    .RESET_B(rst_n),
    .Q(\C_out[174] ));
 sky130_fd_sc_hd__dfrtp_2 _29203_ (.CLK(clk),
    .D(_03001_),
    .RESET_B(rst_n),
    .Q(\C_out[175] ));
 sky130_fd_sc_hd__dfrtp_2 _29204_ (.CLK(clk),
    .D(_03002_),
    .RESET_B(rst_n),
    .Q(\C_out[176] ));
 sky130_fd_sc_hd__dfrtp_2 _29205_ (.CLK(clk),
    .D(_03003_),
    .RESET_B(rst_n),
    .Q(\C_out[177] ));
 sky130_fd_sc_hd__dfrtp_2 _29206_ (.CLK(clk),
    .D(_03004_),
    .RESET_B(rst_n),
    .Q(\C_out[178] ));
 sky130_fd_sc_hd__dfrtp_2 _29207_ (.CLK(clk),
    .D(_03005_),
    .RESET_B(rst_n),
    .Q(\C_out[179] ));
 sky130_fd_sc_hd__dfrtp_2 _29208_ (.CLK(clk),
    .D(_03006_),
    .RESET_B(rst_n),
    .Q(\C_out[180] ));
 sky130_fd_sc_hd__dfrtp_2 _29209_ (.CLK(clk),
    .D(_03007_),
    .RESET_B(rst_n),
    .Q(\C_out[181] ));
 sky130_fd_sc_hd__dfrtp_2 _29210_ (.CLK(clk),
    .D(_03008_),
    .RESET_B(rst_n),
    .Q(\C_out[182] ));
 sky130_fd_sc_hd__dfrtp_2 _29211_ (.CLK(clk),
    .D(_03009_),
    .RESET_B(rst_n),
    .Q(\C_out[183] ));
 sky130_fd_sc_hd__dfrtp_2 _29212_ (.CLK(clk),
    .D(_03010_),
    .RESET_B(rst_n),
    .Q(\C_out[184] ));
 sky130_fd_sc_hd__dfrtp_2 _29213_ (.CLK(clk),
    .D(_03011_),
    .RESET_B(rst_n),
    .Q(\C_out[185] ));
 sky130_fd_sc_hd__dfrtp_2 _29214_ (.CLK(clk),
    .D(_03012_),
    .RESET_B(rst_n),
    .Q(\C_out[186] ));
 sky130_fd_sc_hd__dfrtp_2 _29215_ (.CLK(clk),
    .D(_03013_),
    .RESET_B(rst_n),
    .Q(\C_out[187] ));
 sky130_fd_sc_hd__dfrtp_2 _29216_ (.CLK(clk),
    .D(_03014_),
    .RESET_B(rst_n),
    .Q(\C_out[188] ));
 sky130_fd_sc_hd__dfrtp_2 _29217_ (.CLK(clk),
    .D(_03015_),
    .RESET_B(rst_n),
    .Q(\C_out[189] ));
 sky130_fd_sc_hd__dfrtp_2 _29218_ (.CLK(clk),
    .D(_03016_),
    .RESET_B(rst_n),
    .Q(\C_out[190] ));
 sky130_fd_sc_hd__dfrtp_2 _29219_ (.CLK(clk),
    .D(_03017_),
    .RESET_B(rst_n),
    .Q(\C_out[191] ));
 sky130_fd_sc_hd__dfrtp_2 _29220_ (.CLK(clk),
    .D(_03018_),
    .RESET_B(rst_n),
    .Q(\C_out[192] ));
 sky130_fd_sc_hd__dfrtp_2 _29221_ (.CLK(clk),
    .D(_03019_),
    .RESET_B(rst_n),
    .Q(\C_out[193] ));
 sky130_fd_sc_hd__dfrtp_2 _29222_ (.CLK(clk),
    .D(_03020_),
    .RESET_B(rst_n),
    .Q(\C_out[194] ));
 sky130_fd_sc_hd__dfrtp_2 _29223_ (.CLK(clk),
    .D(_03021_),
    .RESET_B(rst_n),
    .Q(\C_out[195] ));
 sky130_fd_sc_hd__dfrtp_2 _29224_ (.CLK(clk),
    .D(_03022_),
    .RESET_B(rst_n),
    .Q(\C_out[196] ));
 sky130_fd_sc_hd__dfrtp_2 _29225_ (.CLK(clk),
    .D(_03023_),
    .RESET_B(rst_n),
    .Q(\C_out[197] ));
 sky130_fd_sc_hd__dfrtp_2 _29226_ (.CLK(clk),
    .D(_03024_),
    .RESET_B(rst_n),
    .Q(\C_out[198] ));
 sky130_fd_sc_hd__dfrtp_2 _29227_ (.CLK(clk),
    .D(_03025_),
    .RESET_B(rst_n),
    .Q(\C_out[199] ));
 sky130_fd_sc_hd__dfrtp_2 _29228_ (.CLK(clk),
    .D(_03026_),
    .RESET_B(rst_n),
    .Q(\C_out[200] ));
 sky130_fd_sc_hd__dfrtp_2 _29229_ (.CLK(clk),
    .D(_03027_),
    .RESET_B(rst_n),
    .Q(\C_out[201] ));
 sky130_fd_sc_hd__dfrtp_2 _29230_ (.CLK(clk),
    .D(_03028_),
    .RESET_B(rst_n),
    .Q(\C_out[202] ));
 sky130_fd_sc_hd__dfrtp_2 _29231_ (.CLK(clk),
    .D(_03029_),
    .RESET_B(rst_n),
    .Q(\C_out[203] ));
 sky130_fd_sc_hd__dfrtp_2 _29232_ (.CLK(clk),
    .D(_03030_),
    .RESET_B(rst_n),
    .Q(\C_out[204] ));
 sky130_fd_sc_hd__dfrtp_2 _29233_ (.CLK(clk),
    .D(_03031_),
    .RESET_B(rst_n),
    .Q(\C_out[205] ));
 sky130_fd_sc_hd__dfrtp_2 _29234_ (.CLK(clk),
    .D(_03032_),
    .RESET_B(rst_n),
    .Q(\C_out[206] ));
 sky130_fd_sc_hd__dfrtp_2 _29235_ (.CLK(clk),
    .D(_03033_),
    .RESET_B(rst_n),
    .Q(\C_out[207] ));
 sky130_fd_sc_hd__dfrtp_2 _29236_ (.CLK(clk),
    .D(_03034_),
    .RESET_B(rst_n),
    .Q(\C_out[208] ));
 sky130_fd_sc_hd__dfrtp_2 _29237_ (.CLK(clk),
    .D(_03035_),
    .RESET_B(rst_n),
    .Q(\C_out[209] ));
 sky130_fd_sc_hd__dfrtp_2 _29238_ (.CLK(clk),
    .D(_03036_),
    .RESET_B(rst_n),
    .Q(\C_out[210] ));
 sky130_fd_sc_hd__dfrtp_2 _29239_ (.CLK(clk),
    .D(_03037_),
    .RESET_B(rst_n),
    .Q(\C_out[211] ));
 sky130_fd_sc_hd__dfrtp_2 _29240_ (.CLK(clk),
    .D(_03038_),
    .RESET_B(rst_n),
    .Q(\C_out[212] ));
 sky130_fd_sc_hd__dfrtp_2 _29241_ (.CLK(clk),
    .D(_03039_),
    .RESET_B(rst_n),
    .Q(\C_out[213] ));
 sky130_fd_sc_hd__dfrtp_2 _29242_ (.CLK(clk),
    .D(_03040_),
    .RESET_B(rst_n),
    .Q(\C_out[214] ));
 sky130_fd_sc_hd__dfrtp_2 _29243_ (.CLK(clk),
    .D(_03041_),
    .RESET_B(rst_n),
    .Q(\C_out[215] ));
 sky130_fd_sc_hd__dfrtp_2 _29244_ (.CLK(clk),
    .D(_03042_),
    .RESET_B(rst_n),
    .Q(\C_out[216] ));
 sky130_fd_sc_hd__dfrtp_2 _29245_ (.CLK(clk),
    .D(_03043_),
    .RESET_B(rst_n),
    .Q(\C_out[217] ));
 sky130_fd_sc_hd__dfrtp_2 _29246_ (.CLK(clk),
    .D(_03044_),
    .RESET_B(rst_n),
    .Q(\C_out[218] ));
 sky130_fd_sc_hd__dfrtp_2 _29247_ (.CLK(clk),
    .D(_03045_),
    .RESET_B(rst_n),
    .Q(\C_out[219] ));
 sky130_fd_sc_hd__dfrtp_2 _29248_ (.CLK(clk),
    .D(_03046_),
    .RESET_B(rst_n),
    .Q(\C_out[220] ));
 sky130_fd_sc_hd__dfrtp_2 _29249_ (.CLK(clk),
    .D(_03047_),
    .RESET_B(rst_n),
    .Q(\C_out[221] ));
 sky130_fd_sc_hd__dfrtp_2 _29250_ (.CLK(clk),
    .D(_03048_),
    .RESET_B(rst_n),
    .Q(\C_out[222] ));
 sky130_fd_sc_hd__dfrtp_2 _29251_ (.CLK(clk),
    .D(_03049_),
    .RESET_B(rst_n),
    .Q(\C_out[223] ));
 sky130_fd_sc_hd__dfrtp_2 _29252_ (.CLK(clk),
    .D(_03050_),
    .RESET_B(rst_n),
    .Q(\C_out[224] ));
 sky130_fd_sc_hd__dfrtp_2 _29253_ (.CLK(clk),
    .D(_03051_),
    .RESET_B(rst_n),
    .Q(\C_out[225] ));
 sky130_fd_sc_hd__dfrtp_2 _29254_ (.CLK(clk),
    .D(_03052_),
    .RESET_B(rst_n),
    .Q(\C_out[226] ));
 sky130_fd_sc_hd__dfrtp_2 _29255_ (.CLK(clk),
    .D(_03053_),
    .RESET_B(rst_n),
    .Q(\C_out[227] ));
 sky130_fd_sc_hd__dfrtp_2 _29256_ (.CLK(clk),
    .D(_03054_),
    .RESET_B(rst_n),
    .Q(\C_out[228] ));
 sky130_fd_sc_hd__dfrtp_2 _29257_ (.CLK(clk),
    .D(_03055_),
    .RESET_B(rst_n),
    .Q(\C_out[229] ));
 sky130_fd_sc_hd__dfrtp_2 _29258_ (.CLK(clk),
    .D(_03056_),
    .RESET_B(rst_n),
    .Q(\C_out[230] ));
 sky130_fd_sc_hd__dfrtp_2 _29259_ (.CLK(clk),
    .D(_03057_),
    .RESET_B(rst_n),
    .Q(\C_out[231] ));
 sky130_fd_sc_hd__dfrtp_2 _29260_ (.CLK(clk),
    .D(_03058_),
    .RESET_B(rst_n),
    .Q(\C_out[232] ));
 sky130_fd_sc_hd__dfrtp_2 _29261_ (.CLK(clk),
    .D(_03059_),
    .RESET_B(rst_n),
    .Q(\C_out[233] ));
 sky130_fd_sc_hd__dfrtp_2 _29262_ (.CLK(clk),
    .D(_03060_),
    .RESET_B(rst_n),
    .Q(\C_out[234] ));
 sky130_fd_sc_hd__dfrtp_2 _29263_ (.CLK(clk),
    .D(_03061_),
    .RESET_B(rst_n),
    .Q(\C_out[235] ));
 sky130_fd_sc_hd__dfrtp_2 _29264_ (.CLK(clk),
    .D(_03062_),
    .RESET_B(rst_n),
    .Q(\C_out[236] ));
 sky130_fd_sc_hd__dfrtp_2 _29265_ (.CLK(clk),
    .D(_03063_),
    .RESET_B(rst_n),
    .Q(\C_out[237] ));
 sky130_fd_sc_hd__dfrtp_2 _29266_ (.CLK(clk),
    .D(_03064_),
    .RESET_B(rst_n),
    .Q(\C_out[238] ));
 sky130_fd_sc_hd__dfrtp_2 _29267_ (.CLK(clk),
    .D(_03065_),
    .RESET_B(rst_n),
    .Q(\C_out[239] ));
 sky130_fd_sc_hd__dfrtp_2 _29268_ (.CLK(clk),
    .D(_03066_),
    .RESET_B(rst_n),
    .Q(\C_out[240] ));
 sky130_fd_sc_hd__dfrtp_2 _29269_ (.CLK(clk),
    .D(_03067_),
    .RESET_B(rst_n),
    .Q(\C_out[241] ));
 sky130_fd_sc_hd__dfrtp_2 _29270_ (.CLK(clk),
    .D(_03068_),
    .RESET_B(rst_n),
    .Q(\C_out[242] ));
 sky130_fd_sc_hd__dfrtp_2 _29271_ (.CLK(clk),
    .D(_03069_),
    .RESET_B(rst_n),
    .Q(\C_out[243] ));
 sky130_fd_sc_hd__dfrtp_2 _29272_ (.CLK(clk),
    .D(_03070_),
    .RESET_B(rst_n),
    .Q(\C_out[244] ));
 sky130_fd_sc_hd__dfrtp_2 _29273_ (.CLK(clk),
    .D(_03071_),
    .RESET_B(rst_n),
    .Q(\C_out[245] ));
 sky130_fd_sc_hd__dfrtp_2 _29274_ (.CLK(clk),
    .D(_03072_),
    .RESET_B(rst_n),
    .Q(\C_out[246] ));
 sky130_fd_sc_hd__dfrtp_2 _29275_ (.CLK(clk),
    .D(_03073_),
    .RESET_B(rst_n),
    .Q(\C_out[247] ));
 sky130_fd_sc_hd__dfrtp_2 _29276_ (.CLK(clk),
    .D(_03074_),
    .RESET_B(rst_n),
    .Q(\C_out[248] ));
 sky130_fd_sc_hd__dfrtp_2 _29277_ (.CLK(clk),
    .D(_03075_),
    .RESET_B(rst_n),
    .Q(\C_out[249] ));
 sky130_fd_sc_hd__dfrtp_2 _29278_ (.CLK(clk),
    .D(_03076_),
    .RESET_B(rst_n),
    .Q(\C_out[250] ));
 sky130_fd_sc_hd__dfrtp_2 _29279_ (.CLK(clk),
    .D(_03077_),
    .RESET_B(rst_n),
    .Q(\C_out[251] ));
 sky130_fd_sc_hd__dfrtp_2 _29280_ (.CLK(clk),
    .D(_03078_),
    .RESET_B(rst_n),
    .Q(\C_out[252] ));
 sky130_fd_sc_hd__dfrtp_2 _29281_ (.CLK(clk),
    .D(_03079_),
    .RESET_B(rst_n),
    .Q(\C_out[253] ));
 sky130_fd_sc_hd__dfrtp_2 _29282_ (.CLK(clk),
    .D(_03080_),
    .RESET_B(rst_n),
    .Q(\C_out[254] ));
 sky130_fd_sc_hd__dfrtp_2 _29283_ (.CLK(clk),
    .D(_03081_),
    .RESET_B(rst_n),
    .Q(\C_out[255] ));
 sky130_fd_sc_hd__dfrtp_2 _29284_ (.CLK(clk),
    .D(_03082_),
    .RESET_B(rst_n),
    .Q(\C_out[256] ));
 sky130_fd_sc_hd__dfrtp_2 _29285_ (.CLK(clk),
    .D(_03083_),
    .RESET_B(rst_n),
    .Q(\C_out[257] ));
 sky130_fd_sc_hd__dfrtp_2 _29286_ (.CLK(clk),
    .D(_03084_),
    .RESET_B(rst_n),
    .Q(\C_out[258] ));
 sky130_fd_sc_hd__dfrtp_2 _29287_ (.CLK(clk),
    .D(_03085_),
    .RESET_B(rst_n),
    .Q(\C_out[259] ));
 sky130_fd_sc_hd__dfrtp_2 _29288_ (.CLK(clk),
    .D(_03086_),
    .RESET_B(rst_n),
    .Q(\C_out[260] ));
 sky130_fd_sc_hd__dfrtp_2 _29289_ (.CLK(clk),
    .D(_03087_),
    .RESET_B(rst_n),
    .Q(\C_out[261] ));
 sky130_fd_sc_hd__dfrtp_2 _29290_ (.CLK(clk),
    .D(_03088_),
    .RESET_B(rst_n),
    .Q(\C_out[262] ));
 sky130_fd_sc_hd__dfrtp_2 _29291_ (.CLK(clk),
    .D(_03089_),
    .RESET_B(rst_n),
    .Q(\C_out[263] ));
 sky130_fd_sc_hd__dfrtp_2 _29292_ (.CLK(clk),
    .D(_03090_),
    .RESET_B(rst_n),
    .Q(\C_out[264] ));
 sky130_fd_sc_hd__dfrtp_2 _29293_ (.CLK(clk),
    .D(_03091_),
    .RESET_B(rst_n),
    .Q(\C_out[265] ));
 sky130_fd_sc_hd__dfrtp_2 _29294_ (.CLK(clk),
    .D(_03092_),
    .RESET_B(rst_n),
    .Q(\C_out[266] ));
 sky130_fd_sc_hd__dfrtp_2 _29295_ (.CLK(clk),
    .D(_03093_),
    .RESET_B(rst_n),
    .Q(\C_out[267] ));
 sky130_fd_sc_hd__dfrtp_2 _29296_ (.CLK(clk),
    .D(_03094_),
    .RESET_B(rst_n),
    .Q(\C_out[268] ));
 sky130_fd_sc_hd__dfrtp_2 _29297_ (.CLK(clk),
    .D(_03095_),
    .RESET_B(rst_n),
    .Q(\C_out[269] ));
 sky130_fd_sc_hd__dfrtp_2 _29298_ (.CLK(clk),
    .D(_03096_),
    .RESET_B(rst_n),
    .Q(\C_out[270] ));
 sky130_fd_sc_hd__dfrtp_2 _29299_ (.CLK(clk),
    .D(_03097_),
    .RESET_B(rst_n),
    .Q(\C_out[271] ));
 sky130_fd_sc_hd__dfrtp_2 _29300_ (.CLK(clk),
    .D(_03098_),
    .RESET_B(rst_n),
    .Q(\C_out[272] ));
 sky130_fd_sc_hd__dfrtp_2 _29301_ (.CLK(clk),
    .D(_03099_),
    .RESET_B(rst_n),
    .Q(\C_out[273] ));
 sky130_fd_sc_hd__dfrtp_2 _29302_ (.CLK(clk),
    .D(_03100_),
    .RESET_B(rst_n),
    .Q(\C_out[274] ));
 sky130_fd_sc_hd__dfrtp_2 _29303_ (.CLK(clk),
    .D(_03101_),
    .RESET_B(rst_n),
    .Q(\C_out[275] ));
 sky130_fd_sc_hd__dfrtp_2 _29304_ (.CLK(clk),
    .D(_03102_),
    .RESET_B(rst_n),
    .Q(\C_out[276] ));
 sky130_fd_sc_hd__dfrtp_2 _29305_ (.CLK(clk),
    .D(_03103_),
    .RESET_B(rst_n),
    .Q(\C_out[277] ));
 sky130_fd_sc_hd__dfrtp_2 _29306_ (.CLK(clk),
    .D(_03104_),
    .RESET_B(rst_n),
    .Q(\C_out[278] ));
 sky130_fd_sc_hd__dfrtp_2 _29307_ (.CLK(clk),
    .D(_03105_),
    .RESET_B(rst_n),
    .Q(\C_out[279] ));
 sky130_fd_sc_hd__dfrtp_2 _29308_ (.CLK(clk),
    .D(_03106_),
    .RESET_B(rst_n),
    .Q(\C_out[280] ));
 sky130_fd_sc_hd__dfrtp_2 _29309_ (.CLK(clk),
    .D(_03107_),
    .RESET_B(rst_n),
    .Q(\C_out[281] ));
 sky130_fd_sc_hd__dfrtp_2 _29310_ (.CLK(clk),
    .D(_03108_),
    .RESET_B(rst_n),
    .Q(\C_out[282] ));
 sky130_fd_sc_hd__dfrtp_2 _29311_ (.CLK(clk),
    .D(_03109_),
    .RESET_B(rst_n),
    .Q(\C_out[283] ));
 sky130_fd_sc_hd__dfrtp_2 _29312_ (.CLK(clk),
    .D(_03110_),
    .RESET_B(rst_n),
    .Q(\C_out[284] ));
 sky130_fd_sc_hd__dfrtp_2 _29313_ (.CLK(clk),
    .D(_03111_),
    .RESET_B(rst_n),
    .Q(\C_out[285] ));
 sky130_fd_sc_hd__dfrtp_2 _29314_ (.CLK(clk),
    .D(_03112_),
    .RESET_B(rst_n),
    .Q(\C_out[286] ));
 sky130_fd_sc_hd__dfrtp_2 _29315_ (.CLK(clk),
    .D(_03113_),
    .RESET_B(rst_n),
    .Q(\C_out[287] ));
 sky130_fd_sc_hd__dfrtp_2 _29316_ (.CLK(clk),
    .D(_03114_),
    .RESET_B(rst_n),
    .Q(\C_out[288] ));
 sky130_fd_sc_hd__dfrtp_2 _29317_ (.CLK(clk),
    .D(_03115_),
    .RESET_B(rst_n),
    .Q(\C_out[289] ));
 sky130_fd_sc_hd__dfrtp_2 _29318_ (.CLK(clk),
    .D(_03116_),
    .RESET_B(rst_n),
    .Q(\C_out[290] ));
 sky130_fd_sc_hd__dfrtp_2 _29319_ (.CLK(clk),
    .D(_03117_),
    .RESET_B(rst_n),
    .Q(\C_out[291] ));
 sky130_fd_sc_hd__dfrtp_2 _29320_ (.CLK(clk),
    .D(_03118_),
    .RESET_B(rst_n),
    .Q(\C_out[292] ));
 sky130_fd_sc_hd__dfrtp_2 _29321_ (.CLK(clk),
    .D(_03119_),
    .RESET_B(rst_n),
    .Q(\C_out[293] ));
 sky130_fd_sc_hd__dfrtp_2 _29322_ (.CLK(clk),
    .D(_03120_),
    .RESET_B(rst_n),
    .Q(\C_out[294] ));
 sky130_fd_sc_hd__dfrtp_2 _29323_ (.CLK(clk),
    .D(_03121_),
    .RESET_B(rst_n),
    .Q(\C_out[295] ));
 sky130_fd_sc_hd__dfrtp_2 _29324_ (.CLK(clk),
    .D(_03122_),
    .RESET_B(rst_n),
    .Q(\C_out[296] ));
 sky130_fd_sc_hd__dfrtp_2 _29325_ (.CLK(clk),
    .D(_03123_),
    .RESET_B(rst_n),
    .Q(\C_out[297] ));
 sky130_fd_sc_hd__dfrtp_2 _29326_ (.CLK(clk),
    .D(_03124_),
    .RESET_B(rst_n),
    .Q(\C_out[298] ));
 sky130_fd_sc_hd__dfrtp_2 _29327_ (.CLK(clk),
    .D(_03125_),
    .RESET_B(rst_n),
    .Q(\C_out[299] ));
 sky130_fd_sc_hd__dfrtp_2 _29328_ (.CLK(clk),
    .D(_03126_),
    .RESET_B(rst_n),
    .Q(\C_out[300] ));
 sky130_fd_sc_hd__dfrtp_2 _29329_ (.CLK(clk),
    .D(_03127_),
    .RESET_B(rst_n),
    .Q(\C_out[301] ));
 sky130_fd_sc_hd__dfrtp_2 _29330_ (.CLK(clk),
    .D(_03128_),
    .RESET_B(rst_n),
    .Q(\C_out[302] ));
 sky130_fd_sc_hd__dfrtp_2 _29331_ (.CLK(clk),
    .D(_03129_),
    .RESET_B(rst_n),
    .Q(\C_out[303] ));
 sky130_fd_sc_hd__dfrtp_2 _29332_ (.CLK(clk),
    .D(_03130_),
    .RESET_B(rst_n),
    .Q(\C_out[304] ));
 sky130_fd_sc_hd__dfrtp_2 _29333_ (.CLK(clk),
    .D(_03131_),
    .RESET_B(rst_n),
    .Q(\C_out[305] ));
 sky130_fd_sc_hd__dfrtp_2 _29334_ (.CLK(clk),
    .D(_03132_),
    .RESET_B(rst_n),
    .Q(\C_out[306] ));
 sky130_fd_sc_hd__dfrtp_2 _29335_ (.CLK(clk),
    .D(_03133_),
    .RESET_B(rst_n),
    .Q(\C_out[307] ));
 sky130_fd_sc_hd__dfrtp_2 _29336_ (.CLK(clk),
    .D(_03134_),
    .RESET_B(rst_n),
    .Q(\C_out[308] ));
 sky130_fd_sc_hd__dfrtp_2 _29337_ (.CLK(clk),
    .D(_03135_),
    .RESET_B(rst_n),
    .Q(\C_out[309] ));
 sky130_fd_sc_hd__dfrtp_2 _29338_ (.CLK(clk),
    .D(_03136_),
    .RESET_B(rst_n),
    .Q(\C_out[310] ));
 sky130_fd_sc_hd__dfrtp_2 _29339_ (.CLK(clk),
    .D(_03137_),
    .RESET_B(rst_n),
    .Q(\C_out[311] ));
 sky130_fd_sc_hd__dfrtp_2 _29340_ (.CLK(clk),
    .D(_03138_),
    .RESET_B(rst_n),
    .Q(\C_out[312] ));
 sky130_fd_sc_hd__dfrtp_2 _29341_ (.CLK(clk),
    .D(_03139_),
    .RESET_B(rst_n),
    .Q(\C_out[313] ));
 sky130_fd_sc_hd__dfrtp_2 _29342_ (.CLK(clk),
    .D(_03140_),
    .RESET_B(rst_n),
    .Q(\C_out[314] ));
 sky130_fd_sc_hd__dfrtp_2 _29343_ (.CLK(clk),
    .D(_03141_),
    .RESET_B(rst_n),
    .Q(\C_out[315] ));
 sky130_fd_sc_hd__dfrtp_2 _29344_ (.CLK(clk),
    .D(_03142_),
    .RESET_B(rst_n),
    .Q(\C_out[316] ));
 sky130_fd_sc_hd__dfrtp_2 _29345_ (.CLK(clk),
    .D(_03143_),
    .RESET_B(rst_n),
    .Q(\C_out[317] ));
 sky130_fd_sc_hd__dfrtp_2 _29346_ (.CLK(clk),
    .D(_03144_),
    .RESET_B(rst_n),
    .Q(\C_out[318] ));
 sky130_fd_sc_hd__dfrtp_2 _29347_ (.CLK(clk),
    .D(_03145_),
    .RESET_B(rst_n),
    .Q(\C_out[319] ));
 sky130_fd_sc_hd__dfrtp_2 _29348_ (.CLK(clk),
    .D(_03146_),
    .RESET_B(rst_n),
    .Q(\C_out[320] ));
 sky130_fd_sc_hd__dfrtp_2 _29349_ (.CLK(clk),
    .D(_03147_),
    .RESET_B(rst_n),
    .Q(\C_out[321] ));
 sky130_fd_sc_hd__dfrtp_2 _29350_ (.CLK(clk),
    .D(_03148_),
    .RESET_B(rst_n),
    .Q(\C_out[322] ));
 sky130_fd_sc_hd__dfrtp_2 _29351_ (.CLK(clk),
    .D(_03149_),
    .RESET_B(rst_n),
    .Q(\C_out[323] ));
 sky130_fd_sc_hd__dfrtp_2 _29352_ (.CLK(clk),
    .D(_03150_),
    .RESET_B(rst_n),
    .Q(\C_out[324] ));
 sky130_fd_sc_hd__dfrtp_2 _29353_ (.CLK(clk),
    .D(_03151_),
    .RESET_B(rst_n),
    .Q(\C_out[325] ));
 sky130_fd_sc_hd__dfrtp_2 _29354_ (.CLK(clk),
    .D(_03152_),
    .RESET_B(rst_n),
    .Q(\C_out[326] ));
 sky130_fd_sc_hd__dfrtp_2 _29355_ (.CLK(clk),
    .D(_03153_),
    .RESET_B(rst_n),
    .Q(\C_out[327] ));
 sky130_fd_sc_hd__dfrtp_2 _29356_ (.CLK(clk),
    .D(_03154_),
    .RESET_B(rst_n),
    .Q(\C_out[328] ));
 sky130_fd_sc_hd__dfrtp_2 _29357_ (.CLK(clk),
    .D(_03155_),
    .RESET_B(rst_n),
    .Q(\C_out[329] ));
 sky130_fd_sc_hd__dfrtp_2 _29358_ (.CLK(clk),
    .D(_03156_),
    .RESET_B(rst_n),
    .Q(\C_out[330] ));
 sky130_fd_sc_hd__dfrtp_2 _29359_ (.CLK(clk),
    .D(_03157_),
    .RESET_B(rst_n),
    .Q(\C_out[331] ));
 sky130_fd_sc_hd__dfrtp_2 _29360_ (.CLK(clk),
    .D(_03158_),
    .RESET_B(rst_n),
    .Q(\C_out[332] ));
 sky130_fd_sc_hd__dfrtp_2 _29361_ (.CLK(clk),
    .D(_03159_),
    .RESET_B(rst_n),
    .Q(\C_out[333] ));
 sky130_fd_sc_hd__dfrtp_2 _29362_ (.CLK(clk),
    .D(_03160_),
    .RESET_B(rst_n),
    .Q(\C_out[334] ));
 sky130_fd_sc_hd__dfrtp_2 _29363_ (.CLK(clk),
    .D(_03161_),
    .RESET_B(rst_n),
    .Q(\C_out[335] ));
 sky130_fd_sc_hd__dfrtp_2 _29364_ (.CLK(clk),
    .D(_03162_),
    .RESET_B(rst_n),
    .Q(\C_out[336] ));
 sky130_fd_sc_hd__dfrtp_2 _29365_ (.CLK(clk),
    .D(_03163_),
    .RESET_B(rst_n),
    .Q(\C_out[337] ));
 sky130_fd_sc_hd__dfrtp_2 _29366_ (.CLK(clk),
    .D(_03164_),
    .RESET_B(rst_n),
    .Q(\C_out[338] ));
 sky130_fd_sc_hd__dfrtp_2 _29367_ (.CLK(clk),
    .D(_03165_),
    .RESET_B(rst_n),
    .Q(\C_out[339] ));
 sky130_fd_sc_hd__dfrtp_2 _29368_ (.CLK(clk),
    .D(_03166_),
    .RESET_B(rst_n),
    .Q(\C_out[340] ));
 sky130_fd_sc_hd__dfrtp_2 _29369_ (.CLK(clk),
    .D(_03167_),
    .RESET_B(rst_n),
    .Q(\C_out[341] ));
 sky130_fd_sc_hd__dfrtp_2 _29370_ (.CLK(clk),
    .D(_03168_),
    .RESET_B(rst_n),
    .Q(\C_out[342] ));
 sky130_fd_sc_hd__dfrtp_2 _29371_ (.CLK(clk),
    .D(_03169_),
    .RESET_B(rst_n),
    .Q(\C_out[343] ));
 sky130_fd_sc_hd__dfrtp_2 _29372_ (.CLK(clk),
    .D(_03170_),
    .RESET_B(rst_n),
    .Q(\C_out[344] ));
 sky130_fd_sc_hd__dfrtp_2 _29373_ (.CLK(clk),
    .D(_03171_),
    .RESET_B(rst_n),
    .Q(\C_out[345] ));
 sky130_fd_sc_hd__dfrtp_2 _29374_ (.CLK(clk),
    .D(_03172_),
    .RESET_B(rst_n),
    .Q(\C_out[346] ));
 sky130_fd_sc_hd__dfrtp_2 _29375_ (.CLK(clk),
    .D(_03173_),
    .RESET_B(rst_n),
    .Q(\C_out[347] ));
 sky130_fd_sc_hd__dfrtp_2 _29376_ (.CLK(clk),
    .D(_03174_),
    .RESET_B(rst_n),
    .Q(\C_out[348] ));
 sky130_fd_sc_hd__dfrtp_2 _29377_ (.CLK(clk),
    .D(_03175_),
    .RESET_B(rst_n),
    .Q(\C_out[349] ));
 sky130_fd_sc_hd__dfrtp_2 _29378_ (.CLK(clk),
    .D(_03176_),
    .RESET_B(rst_n),
    .Q(\C_out[350] ));
 sky130_fd_sc_hd__dfrtp_2 _29379_ (.CLK(clk),
    .D(_03177_),
    .RESET_B(rst_n),
    .Q(\C_out[351] ));
 sky130_fd_sc_hd__dfrtp_2 _29380_ (.CLK(clk),
    .D(_03178_),
    .RESET_B(rst_n),
    .Q(\C_out[352] ));
 sky130_fd_sc_hd__dfrtp_2 _29381_ (.CLK(clk),
    .D(_03179_),
    .RESET_B(rst_n),
    .Q(\C_out[353] ));
 sky130_fd_sc_hd__dfrtp_2 _29382_ (.CLK(clk),
    .D(_03180_),
    .RESET_B(rst_n),
    .Q(\C_out[354] ));
 sky130_fd_sc_hd__dfrtp_2 _29383_ (.CLK(clk),
    .D(_03181_),
    .RESET_B(rst_n),
    .Q(\C_out[355] ));
 sky130_fd_sc_hd__dfrtp_2 _29384_ (.CLK(clk),
    .D(_03182_),
    .RESET_B(rst_n),
    .Q(\C_out[356] ));
 sky130_fd_sc_hd__dfrtp_2 _29385_ (.CLK(clk),
    .D(_03183_),
    .RESET_B(rst_n),
    .Q(\C_out[357] ));
 sky130_fd_sc_hd__dfrtp_2 _29386_ (.CLK(clk),
    .D(_03184_),
    .RESET_B(rst_n),
    .Q(\C_out[358] ));
 sky130_fd_sc_hd__dfrtp_2 _29387_ (.CLK(clk),
    .D(_03185_),
    .RESET_B(rst_n),
    .Q(\C_out[359] ));
 sky130_fd_sc_hd__dfrtp_2 _29388_ (.CLK(clk),
    .D(_03186_),
    .RESET_B(rst_n),
    .Q(\C_out[360] ));
 sky130_fd_sc_hd__dfrtp_2 _29389_ (.CLK(clk),
    .D(_03187_),
    .RESET_B(rst_n),
    .Q(\C_out[361] ));
 sky130_fd_sc_hd__dfrtp_2 _29390_ (.CLK(clk),
    .D(_03188_),
    .RESET_B(rst_n),
    .Q(\C_out[362] ));
 sky130_fd_sc_hd__dfrtp_2 _29391_ (.CLK(clk),
    .D(_03189_),
    .RESET_B(rst_n),
    .Q(\C_out[363] ));
 sky130_fd_sc_hd__dfrtp_2 _29392_ (.CLK(clk),
    .D(_03190_),
    .RESET_B(rst_n),
    .Q(\C_out[364] ));
 sky130_fd_sc_hd__dfrtp_2 _29393_ (.CLK(clk),
    .D(_03191_),
    .RESET_B(rst_n),
    .Q(\C_out[365] ));
 sky130_fd_sc_hd__dfrtp_2 _29394_ (.CLK(clk),
    .D(_03192_),
    .RESET_B(rst_n),
    .Q(\C_out[366] ));
 sky130_fd_sc_hd__dfrtp_2 _29395_ (.CLK(clk),
    .D(_03193_),
    .RESET_B(rst_n),
    .Q(\C_out[367] ));
 sky130_fd_sc_hd__dfrtp_2 _29396_ (.CLK(clk),
    .D(_03194_),
    .RESET_B(rst_n),
    .Q(\C_out[368] ));
 sky130_fd_sc_hd__dfrtp_2 _29397_ (.CLK(clk),
    .D(_03195_),
    .RESET_B(rst_n),
    .Q(\C_out[369] ));
 sky130_fd_sc_hd__dfrtp_2 _29398_ (.CLK(clk),
    .D(_03196_),
    .RESET_B(rst_n),
    .Q(\C_out[370] ));
 sky130_fd_sc_hd__dfrtp_2 _29399_ (.CLK(clk),
    .D(_03197_),
    .RESET_B(rst_n),
    .Q(\C_out[371] ));
 sky130_fd_sc_hd__dfrtp_2 _29400_ (.CLK(clk),
    .D(_03198_),
    .RESET_B(rst_n),
    .Q(\C_out[372] ));
 sky130_fd_sc_hd__dfrtp_2 _29401_ (.CLK(clk),
    .D(_03199_),
    .RESET_B(rst_n),
    .Q(\C_out[373] ));
 sky130_fd_sc_hd__dfrtp_2 _29402_ (.CLK(clk),
    .D(_03200_),
    .RESET_B(rst_n),
    .Q(\C_out[374] ));
 sky130_fd_sc_hd__dfrtp_2 _29403_ (.CLK(clk),
    .D(_03201_),
    .RESET_B(rst_n),
    .Q(\C_out[375] ));
 sky130_fd_sc_hd__dfrtp_2 _29404_ (.CLK(clk),
    .D(_03202_),
    .RESET_B(rst_n),
    .Q(\C_out[376] ));
 sky130_fd_sc_hd__dfrtp_2 _29405_ (.CLK(clk),
    .D(_03203_),
    .RESET_B(rst_n),
    .Q(\C_out[377] ));
 sky130_fd_sc_hd__dfrtp_2 _29406_ (.CLK(clk),
    .D(_03204_),
    .RESET_B(rst_n),
    .Q(\C_out[378] ));
 sky130_fd_sc_hd__dfrtp_2 _29407_ (.CLK(clk),
    .D(_03205_),
    .RESET_B(rst_n),
    .Q(\C_out[379] ));
 sky130_fd_sc_hd__dfrtp_2 _29408_ (.CLK(clk),
    .D(_03206_),
    .RESET_B(rst_n),
    .Q(\C_out[380] ));
 sky130_fd_sc_hd__dfrtp_2 _29409_ (.CLK(clk),
    .D(_03207_),
    .RESET_B(rst_n),
    .Q(\C_out[381] ));
 sky130_fd_sc_hd__dfrtp_2 _29410_ (.CLK(clk),
    .D(_03208_),
    .RESET_B(rst_n),
    .Q(\C_out[382] ));
 sky130_fd_sc_hd__dfrtp_2 _29411_ (.CLK(clk),
    .D(_03209_),
    .RESET_B(rst_n),
    .Q(\C_out[383] ));
 sky130_fd_sc_hd__dfrtp_2 _29412_ (.CLK(clk),
    .D(_03210_),
    .RESET_B(rst_n),
    .Q(\C_out[384] ));
 sky130_fd_sc_hd__dfrtp_2 _29413_ (.CLK(clk),
    .D(_03211_),
    .RESET_B(rst_n),
    .Q(\C_out[385] ));
 sky130_fd_sc_hd__dfrtp_2 _29414_ (.CLK(clk),
    .D(_03212_),
    .RESET_B(rst_n),
    .Q(\C_out[386] ));
 sky130_fd_sc_hd__dfrtp_2 _29415_ (.CLK(clk),
    .D(_03213_),
    .RESET_B(rst_n),
    .Q(\C_out[387] ));
 sky130_fd_sc_hd__dfrtp_2 _29416_ (.CLK(clk),
    .D(_03214_),
    .RESET_B(rst_n),
    .Q(\C_out[388] ));
 sky130_fd_sc_hd__dfrtp_2 _29417_ (.CLK(clk),
    .D(_03215_),
    .RESET_B(rst_n),
    .Q(\C_out[389] ));
 sky130_fd_sc_hd__dfrtp_2 _29418_ (.CLK(clk),
    .D(_03216_),
    .RESET_B(rst_n),
    .Q(\C_out[390] ));
 sky130_fd_sc_hd__dfrtp_2 _29419_ (.CLK(clk),
    .D(_03217_),
    .RESET_B(rst_n),
    .Q(\C_out[391] ));
 sky130_fd_sc_hd__dfrtp_2 _29420_ (.CLK(clk),
    .D(_03218_),
    .RESET_B(rst_n),
    .Q(\C_out[392] ));
 sky130_fd_sc_hd__dfrtp_2 _29421_ (.CLK(clk),
    .D(_03219_),
    .RESET_B(rst_n),
    .Q(\C_out[393] ));
 sky130_fd_sc_hd__dfrtp_2 _29422_ (.CLK(clk),
    .D(_03220_),
    .RESET_B(rst_n),
    .Q(\C_out[394] ));
 sky130_fd_sc_hd__dfrtp_2 _29423_ (.CLK(clk),
    .D(_03221_),
    .RESET_B(rst_n),
    .Q(\C_out[395] ));
 sky130_fd_sc_hd__dfrtp_2 _29424_ (.CLK(clk),
    .D(_03222_),
    .RESET_B(rst_n),
    .Q(\C_out[396] ));
 sky130_fd_sc_hd__dfrtp_2 _29425_ (.CLK(clk),
    .D(_03223_),
    .RESET_B(rst_n),
    .Q(\C_out[397] ));
 sky130_fd_sc_hd__dfrtp_2 _29426_ (.CLK(clk),
    .D(_03224_),
    .RESET_B(rst_n),
    .Q(\C_out[398] ));
 sky130_fd_sc_hd__dfrtp_2 _29427_ (.CLK(clk),
    .D(_03225_),
    .RESET_B(rst_n),
    .Q(\C_out[399] ));
 sky130_fd_sc_hd__dfrtp_2 _29428_ (.CLK(clk),
    .D(_03226_),
    .RESET_B(rst_n),
    .Q(\C_out[400] ));
 sky130_fd_sc_hd__dfrtp_2 _29429_ (.CLK(clk),
    .D(_03227_),
    .RESET_B(rst_n),
    .Q(\C_out[401] ));
 sky130_fd_sc_hd__dfrtp_2 _29430_ (.CLK(clk),
    .D(_03228_),
    .RESET_B(rst_n),
    .Q(\C_out[402] ));
 sky130_fd_sc_hd__dfrtp_2 _29431_ (.CLK(clk),
    .D(_03229_),
    .RESET_B(rst_n),
    .Q(\C_out[403] ));
 sky130_fd_sc_hd__dfrtp_2 _29432_ (.CLK(clk),
    .D(_03230_),
    .RESET_B(rst_n),
    .Q(\C_out[404] ));
 sky130_fd_sc_hd__dfrtp_2 _29433_ (.CLK(clk),
    .D(_03231_),
    .RESET_B(rst_n),
    .Q(\C_out[405] ));
 sky130_fd_sc_hd__dfrtp_2 _29434_ (.CLK(clk),
    .D(_03232_),
    .RESET_B(rst_n),
    .Q(\C_out[406] ));
 sky130_fd_sc_hd__dfrtp_2 _29435_ (.CLK(clk),
    .D(_03233_),
    .RESET_B(rst_n),
    .Q(\C_out[407] ));
 sky130_fd_sc_hd__dfrtp_2 _29436_ (.CLK(clk),
    .D(_03234_),
    .RESET_B(rst_n),
    .Q(\C_out[408] ));
 sky130_fd_sc_hd__dfrtp_2 _29437_ (.CLK(clk),
    .D(_03235_),
    .RESET_B(rst_n),
    .Q(\C_out[409] ));
 sky130_fd_sc_hd__dfrtp_2 _29438_ (.CLK(clk),
    .D(_03236_),
    .RESET_B(rst_n),
    .Q(\C_out[410] ));
 sky130_fd_sc_hd__dfrtp_2 _29439_ (.CLK(clk),
    .D(_03237_),
    .RESET_B(rst_n),
    .Q(\C_out[411] ));
 sky130_fd_sc_hd__dfrtp_2 _29440_ (.CLK(clk),
    .D(_03238_),
    .RESET_B(rst_n),
    .Q(\C_out[412] ));
 sky130_fd_sc_hd__dfrtp_2 _29441_ (.CLK(clk),
    .D(_03239_),
    .RESET_B(rst_n),
    .Q(\C_out[413] ));
 sky130_fd_sc_hd__dfrtp_2 _29442_ (.CLK(clk),
    .D(_03240_),
    .RESET_B(rst_n),
    .Q(\C_out[414] ));
 sky130_fd_sc_hd__dfrtp_2 _29443_ (.CLK(clk),
    .D(_03241_),
    .RESET_B(rst_n),
    .Q(\C_out[415] ));
 sky130_fd_sc_hd__dfrtp_2 _29444_ (.CLK(clk),
    .D(_03242_),
    .RESET_B(rst_n),
    .Q(\C_out[416] ));
 sky130_fd_sc_hd__dfrtp_2 _29445_ (.CLK(clk),
    .D(_03243_),
    .RESET_B(rst_n),
    .Q(\C_out[417] ));
 sky130_fd_sc_hd__dfrtp_2 _29446_ (.CLK(clk),
    .D(_03244_),
    .RESET_B(rst_n),
    .Q(\C_out[418] ));
 sky130_fd_sc_hd__dfrtp_2 _29447_ (.CLK(clk),
    .D(_03245_),
    .RESET_B(rst_n),
    .Q(\C_out[419] ));
 sky130_fd_sc_hd__dfrtp_2 _29448_ (.CLK(clk),
    .D(_03246_),
    .RESET_B(rst_n),
    .Q(\C_out[420] ));
 sky130_fd_sc_hd__dfrtp_2 _29449_ (.CLK(clk),
    .D(_03247_),
    .RESET_B(rst_n),
    .Q(\C_out[421] ));
 sky130_fd_sc_hd__dfrtp_2 _29450_ (.CLK(clk),
    .D(_03248_),
    .RESET_B(rst_n),
    .Q(\C_out[422] ));
 sky130_fd_sc_hd__dfrtp_2 _29451_ (.CLK(clk),
    .D(_03249_),
    .RESET_B(rst_n),
    .Q(\C_out[423] ));
 sky130_fd_sc_hd__dfrtp_2 _29452_ (.CLK(clk),
    .D(_03250_),
    .RESET_B(rst_n),
    .Q(\C_out[424] ));
 sky130_fd_sc_hd__dfrtp_2 _29453_ (.CLK(clk),
    .D(_03251_),
    .RESET_B(rst_n),
    .Q(\C_out[425] ));
 sky130_fd_sc_hd__dfrtp_2 _29454_ (.CLK(clk),
    .D(_03252_),
    .RESET_B(rst_n),
    .Q(\C_out[426] ));
 sky130_fd_sc_hd__dfrtp_2 _29455_ (.CLK(clk),
    .D(_03253_),
    .RESET_B(rst_n),
    .Q(\C_out[427] ));
 sky130_fd_sc_hd__dfrtp_2 _29456_ (.CLK(clk),
    .D(_03254_),
    .RESET_B(rst_n),
    .Q(\C_out[428] ));
 sky130_fd_sc_hd__dfrtp_2 _29457_ (.CLK(clk),
    .D(_03255_),
    .RESET_B(rst_n),
    .Q(\C_out[429] ));
 sky130_fd_sc_hd__dfrtp_2 _29458_ (.CLK(clk),
    .D(_03256_),
    .RESET_B(rst_n),
    .Q(\C_out[430] ));
 sky130_fd_sc_hd__dfrtp_2 _29459_ (.CLK(clk),
    .D(_03257_),
    .RESET_B(rst_n),
    .Q(\C_out[431] ));
 sky130_fd_sc_hd__dfrtp_2 _29460_ (.CLK(clk),
    .D(_03258_),
    .RESET_B(rst_n),
    .Q(\C_out[432] ));
 sky130_fd_sc_hd__dfrtp_2 _29461_ (.CLK(clk),
    .D(_03259_),
    .RESET_B(rst_n),
    .Q(\C_out[433] ));
 sky130_fd_sc_hd__dfrtp_2 _29462_ (.CLK(clk),
    .D(_03260_),
    .RESET_B(rst_n),
    .Q(\C_out[434] ));
 sky130_fd_sc_hd__dfrtp_2 _29463_ (.CLK(clk),
    .D(_03261_),
    .RESET_B(rst_n),
    .Q(\C_out[435] ));
 sky130_fd_sc_hd__dfrtp_2 _29464_ (.CLK(clk),
    .D(_03262_),
    .RESET_B(rst_n),
    .Q(\C_out[436] ));
 sky130_fd_sc_hd__dfrtp_2 _29465_ (.CLK(clk),
    .D(_03263_),
    .RESET_B(rst_n),
    .Q(\C_out[437] ));
 sky130_fd_sc_hd__dfrtp_2 _29466_ (.CLK(clk),
    .D(_03264_),
    .RESET_B(rst_n),
    .Q(\C_out[438] ));
 sky130_fd_sc_hd__dfrtp_2 _29467_ (.CLK(clk),
    .D(_03265_),
    .RESET_B(rst_n),
    .Q(\C_out[439] ));
 sky130_fd_sc_hd__dfrtp_2 _29468_ (.CLK(clk),
    .D(_03266_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[440] ));
 sky130_fd_sc_hd__dfrtp_2 _29469_ (.CLK(clk),
    .D(_03267_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[441] ));
 sky130_fd_sc_hd__dfrtp_2 _29470_ (.CLK(clk),
    .D(_03268_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[442] ));
 sky130_fd_sc_hd__dfrtp_2 _29471_ (.CLK(clk),
    .D(_03269_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[443] ));
 sky130_fd_sc_hd__dfrtp_2 _29472_ (.CLK(clk),
    .D(_03270_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[444] ));
 sky130_fd_sc_hd__dfrtp_2 _29473_ (.CLK(clk),
    .D(_03271_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[445] ));
 sky130_fd_sc_hd__dfrtp_2 _29474_ (.CLK(clk),
    .D(_03272_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[446] ));
 sky130_fd_sc_hd__dfrtp_2 _29475_ (.CLK(clk),
    .D(_03273_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[447] ));
 sky130_fd_sc_hd__dfrtp_2 _29476_ (.CLK(clk),
    .D(_03274_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[448] ));
 sky130_fd_sc_hd__dfrtp_2 _29477_ (.CLK(clk),
    .D(_03275_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[449] ));
 sky130_fd_sc_hd__dfrtp_2 _29478_ (.CLK(clk),
    .D(_03276_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[450] ));
 sky130_fd_sc_hd__dfrtp_2 _29479_ (.CLK(clk),
    .D(_03277_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[451] ));
 sky130_fd_sc_hd__dfrtp_2 _29480_ (.CLK(clk),
    .D(_03278_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[452] ));
 sky130_fd_sc_hd__dfrtp_2 _29481_ (.CLK(clk),
    .D(_03279_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[453] ));
 sky130_fd_sc_hd__dfrtp_2 _29482_ (.CLK(clk),
    .D(_03280_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[454] ));
 sky130_fd_sc_hd__dfrtp_2 _29483_ (.CLK(clk),
    .D(_03281_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[455] ));
 sky130_fd_sc_hd__dfrtp_2 _29484_ (.CLK(clk),
    .D(_03282_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[456] ));
 sky130_fd_sc_hd__dfrtp_2 _29485_ (.CLK(clk),
    .D(_03283_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[457] ));
 sky130_fd_sc_hd__dfrtp_2 _29486_ (.CLK(clk),
    .D(_03284_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[458] ));
 sky130_fd_sc_hd__dfrtp_2 _29487_ (.CLK(clk),
    .D(_03285_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[459] ));
 sky130_fd_sc_hd__dfrtp_2 _29488_ (.CLK(clk),
    .D(_03286_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[460] ));
 sky130_fd_sc_hd__dfrtp_2 _29489_ (.CLK(clk),
    .D(_03287_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[461] ));
 sky130_fd_sc_hd__dfrtp_2 _29490_ (.CLK(clk),
    .D(_03288_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[462] ));
 sky130_fd_sc_hd__dfrtp_2 _29491_ (.CLK(clk),
    .D(_03289_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[463] ));
 sky130_fd_sc_hd__dfrtp_2 _29492_ (.CLK(clk),
    .D(_03290_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[464] ));
 sky130_fd_sc_hd__dfrtp_2 _29493_ (.CLK(clk),
    .D(_03291_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[465] ));
 sky130_fd_sc_hd__dfrtp_2 _29494_ (.CLK(clk),
    .D(_03292_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[466] ));
 sky130_fd_sc_hd__dfrtp_2 _29495_ (.CLK(clk),
    .D(_03293_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[467] ));
 sky130_fd_sc_hd__dfrtp_2 _29496_ (.CLK(clk),
    .D(_03294_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[468] ));
 sky130_fd_sc_hd__dfrtp_2 _29497_ (.CLK(clk),
    .D(_03295_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[469] ));
 sky130_fd_sc_hd__dfrtp_2 _29498_ (.CLK(clk),
    .D(_03296_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[470] ));
 sky130_fd_sc_hd__dfrtp_2 _29499_ (.CLK(clk),
    .D(_03297_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[471] ));
 sky130_fd_sc_hd__dfrtp_2 _29500_ (.CLK(clk),
    .D(_03298_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[472] ));
 sky130_fd_sc_hd__dfrtp_2 _29501_ (.CLK(clk),
    .D(_03299_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[473] ));
 sky130_fd_sc_hd__dfrtp_2 _29502_ (.CLK(clk),
    .D(_03300_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[474] ));
 sky130_fd_sc_hd__dfrtp_2 _29503_ (.CLK(clk),
    .D(_03301_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[475] ));
 sky130_fd_sc_hd__dfrtp_2 _29504_ (.CLK(clk),
    .D(_03302_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[476] ));
 sky130_fd_sc_hd__dfrtp_2 _29505_ (.CLK(clk),
    .D(_03303_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[477] ));
 sky130_fd_sc_hd__dfrtp_2 _29506_ (.CLK(clk),
    .D(_03304_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[478] ));
 sky130_fd_sc_hd__dfrtp_2 _29507_ (.CLK(clk),
    .D(_03305_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[479] ));
 sky130_fd_sc_hd__dfrtp_2 _29508_ (.CLK(clk),
    .D(_03306_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[480] ));
 sky130_fd_sc_hd__dfrtp_2 _29509_ (.CLK(clk),
    .D(_03307_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[481] ));
 sky130_fd_sc_hd__dfrtp_2 _29510_ (.CLK(clk),
    .D(_03308_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[482] ));
 sky130_fd_sc_hd__dfrtp_2 _29511_ (.CLK(clk),
    .D(_03309_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[483] ));
 sky130_fd_sc_hd__dfrtp_2 _29512_ (.CLK(clk),
    .D(_03310_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[484] ));
 sky130_fd_sc_hd__dfrtp_2 _29513_ (.CLK(clk),
    .D(_03311_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[485] ));
 sky130_fd_sc_hd__dfrtp_2 _29514_ (.CLK(clk),
    .D(_03312_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[486] ));
 sky130_fd_sc_hd__dfrtp_2 _29515_ (.CLK(clk),
    .D(_03313_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[487] ));
 sky130_fd_sc_hd__dfrtp_2 _29516_ (.CLK(clk),
    .D(_03314_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[488] ));
 sky130_fd_sc_hd__dfrtp_2 _29517_ (.CLK(clk),
    .D(_03315_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[489] ));
 sky130_fd_sc_hd__dfrtp_2 _29518_ (.CLK(clk),
    .D(_03316_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[490] ));
 sky130_fd_sc_hd__dfrtp_2 _29519_ (.CLK(clk),
    .D(_03317_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[491] ));
 sky130_fd_sc_hd__dfrtp_2 _29520_ (.CLK(clk),
    .D(_03318_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[492] ));
 sky130_fd_sc_hd__dfrtp_2 _29521_ (.CLK(clk),
    .D(_03319_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[493] ));
 sky130_fd_sc_hd__dfrtp_2 _29522_ (.CLK(clk),
    .D(_03320_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[494] ));
 sky130_fd_sc_hd__dfrtp_2 _29523_ (.CLK(clk),
    .D(_03321_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[495] ));
 sky130_fd_sc_hd__dfrtp_2 _29524_ (.CLK(clk),
    .D(_03322_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[496] ));
 sky130_fd_sc_hd__dfrtp_2 _29525_ (.CLK(clk),
    .D(_03323_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[497] ));
 sky130_fd_sc_hd__dfrtp_2 _29526_ (.CLK(clk),
    .D(_03324_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[498] ));
 sky130_fd_sc_hd__dfrtp_2 _29527_ (.CLK(clk),
    .D(_03325_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[499] ));
 sky130_fd_sc_hd__dfrtp_2 _29528_ (.CLK(clk),
    .D(_03326_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[500] ));
 sky130_fd_sc_hd__dfrtp_2 _29529_ (.CLK(clk),
    .D(_03327_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[501] ));
 sky130_fd_sc_hd__dfrtp_2 _29530_ (.CLK(clk),
    .D(_03328_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[502] ));
 sky130_fd_sc_hd__dfrtp_2 _29531_ (.CLK(clk),
    .D(_03329_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[503] ));
 sky130_fd_sc_hd__dfrtp_2 _29532_ (.CLK(clk),
    .D(_03330_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[504] ));
 sky130_fd_sc_hd__dfrtp_2 _29533_ (.CLK(clk),
    .D(_03331_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[505] ));
 sky130_fd_sc_hd__dfrtp_2 _29534_ (.CLK(clk),
    .D(_03332_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[506] ));
 sky130_fd_sc_hd__dfrtp_2 _29535_ (.CLK(clk),
    .D(_03333_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[507] ));
 sky130_fd_sc_hd__dfrtp_2 _29536_ (.CLK(clk),
    .D(_03334_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[508] ));
 sky130_fd_sc_hd__dfrtp_2 _29537_ (.CLK(clk),
    .D(_03335_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[509] ));
 sky130_fd_sc_hd__dfrtp_2 _29538_ (.CLK(clk),
    .D(_03336_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[510] ));
 sky130_fd_sc_hd__dfrtp_2 _29539_ (.CLK(clk),
    .D(_03337_),
    .RESET_B(rst_n),
    .Q(\ser_C.parallel_data[511] ));
 sky130_fd_sc_hd__dfrtp_2 _29540_ (.CLK(clk),
    .D(_00008_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.load_acc ));
 sky130_fd_sc_hd__dfrtp_2 _29541_ (.CLK(clk),
    .D(_00009_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.ce_local ));
 sky130_fd_sc_hd__dfrtp_2 _29542_ (.CLK(clk),
    .D(_00000_),
    .RESET_B(rst_n),
    .Q(done));
 sky130_fd_sc_hd__dfrtp_2 _29543_ (.CLK(clk),
    .D(_03338_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[15][0] ));
 sky130_fd_sc_hd__dfrtp_2 _29544_ (.CLK(clk),
    .D(_03339_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[15][1] ));
 sky130_fd_sc_hd__dfrtp_2 _29545_ (.CLK(clk),
    .D(_03340_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[15][2] ));
 sky130_fd_sc_hd__dfrtp_2 _29546_ (.CLK(clk),
    .D(_03341_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[15][3] ));
 sky130_fd_sc_hd__dfrtp_2 _29547_ (.CLK(clk),
    .D(_03342_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[15][4] ));
 sky130_fd_sc_hd__dfrtp_2 _29548_ (.CLK(clk),
    .D(_03343_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[15][5] ));
 sky130_fd_sc_hd__dfrtp_2 _29549_ (.CLK(clk),
    .D(_03344_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[15][6] ));
 sky130_fd_sc_hd__dfrtp_2 _29550_ (.CLK(clk),
    .D(_03345_),
    .RESET_B(rst_n),
    .Q(\systolic_inst.B_outs[15][7] ));
 sky130_fd_sc_hd__dfrtp_2 _29551_ (.CLK(clk),
    .D(_03346_),
    .RESET_B(rst_n),
    .Q(C_out_serial_data));
 sky130_fd_sc_hd__dfrtp_2 _29552_ (.CLK(B_in_serial_clk),
    .D(_03347_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[0] ));
 sky130_fd_sc_hd__dfrtp_2 _29553_ (.CLK(B_in_serial_clk),
    .D(_03348_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[1] ));
 sky130_fd_sc_hd__dfrtp_2 _29554_ (.CLK(B_in_serial_clk),
    .D(_03349_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[2] ));
 sky130_fd_sc_hd__dfrtp_2 _29555_ (.CLK(B_in_serial_clk),
    .D(_03350_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[3] ));
 sky130_fd_sc_hd__dfrtp_2 _29556_ (.CLK(B_in_serial_clk),
    .D(_03351_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[4] ));
 sky130_fd_sc_hd__dfrtp_2 _29557_ (.CLK(B_in_serial_clk),
    .D(_03352_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[5] ));
 sky130_fd_sc_hd__dfrtp_2 _29558_ (.CLK(B_in_serial_clk),
    .D(_03353_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[6] ));
 sky130_fd_sc_hd__dfrtp_2 _29559_ (.CLK(B_in_serial_clk),
    .D(_03354_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[7] ));
 sky130_fd_sc_hd__dfrtp_2 _29560_ (.CLK(B_in_serial_clk),
    .D(_03355_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[8] ));
 sky130_fd_sc_hd__dfrtp_2 _29561_ (.CLK(B_in_serial_clk),
    .D(_03356_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[9] ));
 sky130_fd_sc_hd__dfrtp_2 _29562_ (.CLK(B_in_serial_clk),
    .D(_03357_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[10] ));
 sky130_fd_sc_hd__dfrtp_2 _29563_ (.CLK(B_in_serial_clk),
    .D(_03358_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[11] ));
 sky130_fd_sc_hd__dfrtp_2 _29564_ (.CLK(B_in_serial_clk),
    .D(_03359_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[12] ));
 sky130_fd_sc_hd__dfrtp_2 _29565_ (.CLK(B_in_serial_clk),
    .D(_03360_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[13] ));
 sky130_fd_sc_hd__dfrtp_2 _29566_ (.CLK(B_in_serial_clk),
    .D(_03361_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[14] ));
 sky130_fd_sc_hd__dfrtp_2 _29567_ (.CLK(B_in_serial_clk),
    .D(_03362_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[15] ));
 sky130_fd_sc_hd__dfrtp_2 _29568_ (.CLK(B_in_serial_clk),
    .D(_03363_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[16] ));
 sky130_fd_sc_hd__dfrtp_2 _29569_ (.CLK(B_in_serial_clk),
    .D(_03364_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[17] ));
 sky130_fd_sc_hd__dfrtp_2 _29570_ (.CLK(B_in_serial_clk),
    .D(_03365_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[18] ));
 sky130_fd_sc_hd__dfrtp_2 _29571_ (.CLK(B_in_serial_clk),
    .D(_03366_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[19] ));
 sky130_fd_sc_hd__dfrtp_2 _29572_ (.CLK(B_in_serial_clk),
    .D(_03367_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[20] ));
 sky130_fd_sc_hd__dfrtp_2 _29573_ (.CLK(B_in_serial_clk),
    .D(_03368_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[21] ));
 sky130_fd_sc_hd__dfrtp_2 _29574_ (.CLK(B_in_serial_clk),
    .D(_03369_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[22] ));
 sky130_fd_sc_hd__dfrtp_2 _29575_ (.CLK(B_in_serial_clk),
    .D(_03370_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[23] ));
 sky130_fd_sc_hd__dfrtp_2 _29576_ (.CLK(B_in_serial_clk),
    .D(_03371_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[24] ));
 sky130_fd_sc_hd__dfrtp_2 _29577_ (.CLK(B_in_serial_clk),
    .D(_03372_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[25] ));
 sky130_fd_sc_hd__dfrtp_2 _29578_ (.CLK(B_in_serial_clk),
    .D(_03373_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[26] ));
 sky130_fd_sc_hd__dfrtp_2 _29579_ (.CLK(B_in_serial_clk),
    .D(_03374_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[27] ));
 sky130_fd_sc_hd__dfrtp_2 _29580_ (.CLK(B_in_serial_clk),
    .D(_03375_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[28] ));
 sky130_fd_sc_hd__dfrtp_2 _29581_ (.CLK(B_in_serial_clk),
    .D(_03376_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[29] ));
 sky130_fd_sc_hd__dfrtp_2 _29582_ (.CLK(B_in_serial_clk),
    .D(_03377_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[30] ));
 sky130_fd_sc_hd__dfrtp_2 _29583_ (.CLK(B_in_serial_clk),
    .D(_03378_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[31] ));
 sky130_fd_sc_hd__dfrtp_2 _29584_ (.CLK(B_in_serial_clk),
    .D(_03379_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[32] ));
 sky130_fd_sc_hd__dfrtp_2 _29585_ (.CLK(B_in_serial_clk),
    .D(_03380_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[33] ));
 sky130_fd_sc_hd__dfrtp_2 _29586_ (.CLK(B_in_serial_clk),
    .D(_03381_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[34] ));
 sky130_fd_sc_hd__dfrtp_2 _29587_ (.CLK(B_in_serial_clk),
    .D(_03382_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[35] ));
 sky130_fd_sc_hd__dfrtp_2 _29588_ (.CLK(B_in_serial_clk),
    .D(_03383_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[36] ));
 sky130_fd_sc_hd__dfrtp_2 _29589_ (.CLK(B_in_serial_clk),
    .D(_03384_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[37] ));
 sky130_fd_sc_hd__dfrtp_2 _29590_ (.CLK(B_in_serial_clk),
    .D(_03385_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[38] ));
 sky130_fd_sc_hd__dfrtp_2 _29591_ (.CLK(B_in_serial_clk),
    .D(_03386_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[39] ));
 sky130_fd_sc_hd__dfrtp_2 _29592_ (.CLK(B_in_serial_clk),
    .D(_03387_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[40] ));
 sky130_fd_sc_hd__dfrtp_2 _29593_ (.CLK(B_in_serial_clk),
    .D(_03388_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[41] ));
 sky130_fd_sc_hd__dfrtp_2 _29594_ (.CLK(B_in_serial_clk),
    .D(_03389_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[42] ));
 sky130_fd_sc_hd__dfrtp_2 _29595_ (.CLK(B_in_serial_clk),
    .D(_03390_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[43] ));
 sky130_fd_sc_hd__dfrtp_2 _29596_ (.CLK(B_in_serial_clk),
    .D(_03391_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[44] ));
 sky130_fd_sc_hd__dfrtp_2 _29597_ (.CLK(B_in_serial_clk),
    .D(_03392_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[45] ));
 sky130_fd_sc_hd__dfrtp_2 _29598_ (.CLK(B_in_serial_clk),
    .D(_03393_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[46] ));
 sky130_fd_sc_hd__dfrtp_2 _29599_ (.CLK(B_in_serial_clk),
    .D(_03394_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[47] ));
 sky130_fd_sc_hd__dfrtp_2 _29600_ (.CLK(B_in_serial_clk),
    .D(_03395_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[48] ));
 sky130_fd_sc_hd__dfrtp_2 _29601_ (.CLK(B_in_serial_clk),
    .D(_03396_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[49] ));
 sky130_fd_sc_hd__dfrtp_2 _29602_ (.CLK(B_in_serial_clk),
    .D(_03397_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[50] ));
 sky130_fd_sc_hd__dfrtp_2 _29603_ (.CLK(B_in_serial_clk),
    .D(_03398_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[51] ));
 sky130_fd_sc_hd__dfrtp_2 _29604_ (.CLK(B_in_serial_clk),
    .D(_03399_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[52] ));
 sky130_fd_sc_hd__dfrtp_2 _29605_ (.CLK(B_in_serial_clk),
    .D(_03400_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[53] ));
 sky130_fd_sc_hd__dfrtp_2 _29606_ (.CLK(B_in_serial_clk),
    .D(_03401_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[54] ));
 sky130_fd_sc_hd__dfrtp_2 _29607_ (.CLK(B_in_serial_clk),
    .D(_03402_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[55] ));
 sky130_fd_sc_hd__dfrtp_2 _29608_ (.CLK(B_in_serial_clk),
    .D(_03403_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[56] ));
 sky130_fd_sc_hd__dfrtp_2 _29609_ (.CLK(B_in_serial_clk),
    .D(_03404_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[57] ));
 sky130_fd_sc_hd__dfrtp_2 _29610_ (.CLK(B_in_serial_clk),
    .D(_03405_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[58] ));
 sky130_fd_sc_hd__dfrtp_2 _29611_ (.CLK(B_in_serial_clk),
    .D(_03406_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[59] ));
 sky130_fd_sc_hd__dfrtp_2 _29612_ (.CLK(B_in_serial_clk),
    .D(_03407_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[60] ));
 sky130_fd_sc_hd__dfrtp_2 _29613_ (.CLK(B_in_serial_clk),
    .D(_03408_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[61] ));
 sky130_fd_sc_hd__dfrtp_2 _29614_ (.CLK(B_in_serial_clk),
    .D(_03409_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[62] ));
 sky130_fd_sc_hd__dfrtp_2 _29615_ (.CLK(B_in_serial_clk),
    .D(_03410_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[63] ));
 sky130_fd_sc_hd__dfrtp_2 _29616_ (.CLK(B_in_serial_clk),
    .D(_03411_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[64] ));
 sky130_fd_sc_hd__dfrtp_2 _29617_ (.CLK(B_in_serial_clk),
    .D(_03412_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[65] ));
 sky130_fd_sc_hd__dfrtp_2 _29618_ (.CLK(B_in_serial_clk),
    .D(_03413_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[66] ));
 sky130_fd_sc_hd__dfrtp_2 _29619_ (.CLK(B_in_serial_clk),
    .D(_03414_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[67] ));
 sky130_fd_sc_hd__dfrtp_2 _29620_ (.CLK(B_in_serial_clk),
    .D(_03415_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[68] ));
 sky130_fd_sc_hd__dfrtp_2 _29621_ (.CLK(B_in_serial_clk),
    .D(_03416_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[69] ));
 sky130_fd_sc_hd__dfrtp_2 _29622_ (.CLK(B_in_serial_clk),
    .D(_03417_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[70] ));
 sky130_fd_sc_hd__dfrtp_2 _29623_ (.CLK(B_in_serial_clk),
    .D(_03418_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[71] ));
 sky130_fd_sc_hd__dfrtp_2 _29624_ (.CLK(B_in_serial_clk),
    .D(_03419_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[72] ));
 sky130_fd_sc_hd__dfrtp_2 _29625_ (.CLK(B_in_serial_clk),
    .D(_03420_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[73] ));
 sky130_fd_sc_hd__dfrtp_2 _29626_ (.CLK(B_in_serial_clk),
    .D(_03421_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[74] ));
 sky130_fd_sc_hd__dfrtp_2 _29627_ (.CLK(B_in_serial_clk),
    .D(_03422_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[75] ));
 sky130_fd_sc_hd__dfrtp_2 _29628_ (.CLK(B_in_serial_clk),
    .D(_03423_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[76] ));
 sky130_fd_sc_hd__dfrtp_2 _29629_ (.CLK(B_in_serial_clk),
    .D(_03424_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[77] ));
 sky130_fd_sc_hd__dfrtp_2 _29630_ (.CLK(B_in_serial_clk),
    .D(_03425_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[78] ));
 sky130_fd_sc_hd__dfrtp_2 _29631_ (.CLK(B_in_serial_clk),
    .D(_03426_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[79] ));
 sky130_fd_sc_hd__dfrtp_2 _29632_ (.CLK(B_in_serial_clk),
    .D(_03427_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[80] ));
 sky130_fd_sc_hd__dfrtp_2 _29633_ (.CLK(B_in_serial_clk),
    .D(_03428_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[81] ));
 sky130_fd_sc_hd__dfrtp_2 _29634_ (.CLK(B_in_serial_clk),
    .D(_03429_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[82] ));
 sky130_fd_sc_hd__dfrtp_2 _29635_ (.CLK(B_in_serial_clk),
    .D(_03430_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[83] ));
 sky130_fd_sc_hd__dfrtp_2 _29636_ (.CLK(B_in_serial_clk),
    .D(_03431_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[84] ));
 sky130_fd_sc_hd__dfrtp_2 _29637_ (.CLK(B_in_serial_clk),
    .D(_03432_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[85] ));
 sky130_fd_sc_hd__dfrtp_2 _29638_ (.CLK(B_in_serial_clk),
    .D(_03433_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[86] ));
 sky130_fd_sc_hd__dfrtp_2 _29639_ (.CLK(B_in_serial_clk),
    .D(_03434_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[87] ));
 sky130_fd_sc_hd__dfrtp_2 _29640_ (.CLK(B_in_serial_clk),
    .D(_03435_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[88] ));
 sky130_fd_sc_hd__dfrtp_2 _29641_ (.CLK(B_in_serial_clk),
    .D(_03436_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[89] ));
 sky130_fd_sc_hd__dfrtp_2 _29642_ (.CLK(B_in_serial_clk),
    .D(_03437_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[90] ));
 sky130_fd_sc_hd__dfrtp_2 _29643_ (.CLK(B_in_serial_clk),
    .D(_03438_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[91] ));
 sky130_fd_sc_hd__dfrtp_2 _29644_ (.CLK(B_in_serial_clk),
    .D(_03439_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[92] ));
 sky130_fd_sc_hd__dfrtp_2 _29645_ (.CLK(B_in_serial_clk),
    .D(_03440_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[93] ));
 sky130_fd_sc_hd__dfrtp_2 _29646_ (.CLK(B_in_serial_clk),
    .D(_03441_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[94] ));
 sky130_fd_sc_hd__dfrtp_2 _29647_ (.CLK(B_in_serial_clk),
    .D(_03442_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[95] ));
 sky130_fd_sc_hd__dfrtp_2 _29648_ (.CLK(B_in_serial_clk),
    .D(_03443_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[96] ));
 sky130_fd_sc_hd__dfrtp_2 _29649_ (.CLK(B_in_serial_clk),
    .D(_03444_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[97] ));
 sky130_fd_sc_hd__dfrtp_2 _29650_ (.CLK(B_in_serial_clk),
    .D(_03445_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[98] ));
 sky130_fd_sc_hd__dfrtp_2 _29651_ (.CLK(B_in_serial_clk),
    .D(_03446_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[99] ));
 sky130_fd_sc_hd__dfrtp_2 _29652_ (.CLK(B_in_serial_clk),
    .D(_03447_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[100] ));
 sky130_fd_sc_hd__dfrtp_2 _29653_ (.CLK(B_in_serial_clk),
    .D(_03448_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[101] ));
 sky130_fd_sc_hd__dfrtp_2 _29654_ (.CLK(B_in_serial_clk),
    .D(_03449_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[102] ));
 sky130_fd_sc_hd__dfrtp_2 _29655_ (.CLK(B_in_serial_clk),
    .D(_03450_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[103] ));
 sky130_fd_sc_hd__dfrtp_2 _29656_ (.CLK(B_in_serial_clk),
    .D(_03451_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[104] ));
 sky130_fd_sc_hd__dfrtp_2 _29657_ (.CLK(B_in_serial_clk),
    .D(_03452_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[105] ));
 sky130_fd_sc_hd__dfrtp_2 _29658_ (.CLK(B_in_serial_clk),
    .D(_03453_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[106] ));
 sky130_fd_sc_hd__dfrtp_2 _29659_ (.CLK(B_in_serial_clk),
    .D(_03454_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[107] ));
 sky130_fd_sc_hd__dfrtp_2 _29660_ (.CLK(B_in_serial_clk),
    .D(_03455_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[108] ));
 sky130_fd_sc_hd__dfrtp_2 _29661_ (.CLK(B_in_serial_clk),
    .D(_03456_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[109] ));
 sky130_fd_sc_hd__dfrtp_2 _29662_ (.CLK(B_in_serial_clk),
    .D(_03457_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[110] ));
 sky130_fd_sc_hd__dfrtp_2 _29663_ (.CLK(B_in_serial_clk),
    .D(_03458_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[111] ));
 sky130_fd_sc_hd__dfrtp_2 _29664_ (.CLK(B_in_serial_clk),
    .D(_03459_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[112] ));
 sky130_fd_sc_hd__dfrtp_2 _29665_ (.CLK(B_in_serial_clk),
    .D(_03460_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[113] ));
 sky130_fd_sc_hd__dfrtp_2 _29666_ (.CLK(B_in_serial_clk),
    .D(_03461_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[114] ));
 sky130_fd_sc_hd__dfrtp_2 _29667_ (.CLK(B_in_serial_clk),
    .D(_03462_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[115] ));
 sky130_fd_sc_hd__dfrtp_2 _29668_ (.CLK(B_in_serial_clk),
    .D(_03463_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[116] ));
 sky130_fd_sc_hd__dfrtp_2 _29669_ (.CLK(B_in_serial_clk),
    .D(_03464_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[117] ));
 sky130_fd_sc_hd__dfrtp_2 _29670_ (.CLK(B_in_serial_clk),
    .D(_03465_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[118] ));
 sky130_fd_sc_hd__dfrtp_2 _29671_ (.CLK(B_in_serial_clk),
    .D(_03466_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[119] ));
 sky130_fd_sc_hd__dfrtp_2 _29672_ (.CLK(B_in_serial_clk),
    .D(_03467_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[120] ));
 sky130_fd_sc_hd__dfrtp_2 _29673_ (.CLK(B_in_serial_clk),
    .D(_03468_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[121] ));
 sky130_fd_sc_hd__dfrtp_2 _29674_ (.CLK(B_in_serial_clk),
    .D(_03469_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[122] ));
 sky130_fd_sc_hd__dfrtp_2 _29675_ (.CLK(B_in_serial_clk),
    .D(_03470_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[123] ));
 sky130_fd_sc_hd__dfrtp_2 _29676_ (.CLK(B_in_serial_clk),
    .D(_03471_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[124] ));
 sky130_fd_sc_hd__dfrtp_2 _29677_ (.CLK(B_in_serial_clk),
    .D(_03472_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[125] ));
 sky130_fd_sc_hd__dfrtp_2 _29678_ (.CLK(B_in_serial_clk),
    .D(_03473_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[126] ));
 sky130_fd_sc_hd__dfrtp_2 _29679_ (.CLK(B_in_serial_clk),
    .D(_03474_),
    .RESET_B(rst_n),
    .Q(\deser_B.serial_word[127] ));
 sky130_fd_sc_hd__dfrtp_2 _29680_ (.CLK(clk),
    .D(_03475_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[0] ));
 sky130_fd_sc_hd__dfrtp_2 _29681_ (.CLK(clk),
    .D(_03476_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[1] ));
 sky130_fd_sc_hd__dfrtp_2 _29682_ (.CLK(clk),
    .D(_03477_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[2] ));
 sky130_fd_sc_hd__dfrtp_2 _29683_ (.CLK(clk),
    .D(_03478_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[3] ));
 sky130_fd_sc_hd__dfrtp_2 _29684_ (.CLK(clk),
    .D(_03479_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[4] ));
 sky130_fd_sc_hd__dfrtp_2 _29685_ (.CLK(clk),
    .D(_03480_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[5] ));
 sky130_fd_sc_hd__dfrtp_2 _29686_ (.CLK(clk),
    .D(_03481_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[6] ));
 sky130_fd_sc_hd__dfrtp_2 _29687_ (.CLK(clk),
    .D(_03482_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[7] ));
 sky130_fd_sc_hd__dfrtp_2 _29688_ (.CLK(clk),
    .D(_03483_),
    .RESET_B(rst_n),
    .Q(\ser_C.bit_idx[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29689_ (.CLK(clk),
    .D(_03484_),
    .Q(\systolic_inst.A_shift[30][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29690_ (.CLK(clk),
    .D(_03485_),
    .Q(\systolic_inst.A_shift[30][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29691_ (.CLK(clk),
    .D(_03486_),
    .Q(\systolic_inst.A_shift[30][2] ));
 sky130_fd_sc_hd__dfxtp_2 _29692_ (.CLK(clk),
    .D(_03487_),
    .Q(\systolic_inst.A_shift[30][3] ));
 sky130_fd_sc_hd__dfxtp_2 _29693_ (.CLK(clk),
    .D(_03488_),
    .Q(\systolic_inst.A_shift[30][4] ));
 sky130_fd_sc_hd__dfxtp_2 _29694_ (.CLK(clk),
    .D(_03489_),
    .Q(\systolic_inst.A_shift[30][5] ));
 sky130_fd_sc_hd__dfxtp_2 _29695_ (.CLK(clk),
    .D(_03490_),
    .Q(\systolic_inst.A_shift[30][6] ));
 sky130_fd_sc_hd__dfxtp_2 _29696_ (.CLK(clk),
    .D(_03491_),
    .Q(\systolic_inst.A_shift[30][7] ));
 sky130_fd_sc_hd__dfrtp_2 _29697_ (.CLK(clk),
    .D(_00007_),
    .RESET_B(rst_n),
    .Q(C_out_frame_sync));
 sky130_fd_sc_hd__buf_2 _29698_ (.A(clk),
    .X(C_out_serial_clk));
endmodule
